VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_mattvenn_inverter
  CLASS BLOCK ;
  FOREIGN tt_um_mattvenn_inverter ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 154.870 224.760 155.170 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 158.550 224.760 158.850 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 151.190 224.760 151.490 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.300000 ;
    PORT
      LAYER met4 ;
        RECT 156.560 0.000 157.160 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.180000 ;
    PORT
      LAYER met4 ;
        RECT 134.480 0.000 135.080 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 112.400 0.000 113.000 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 90.320 0.000 90.920 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 68.240 0.000 68.840 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 46.160 0.000 46.760 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 24.080 0.000 24.680 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 2.000 0.000 2.600 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 147.510 224.760 147.810 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 140.150 224.760 140.450 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 136.470 224.760 136.770 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 129.110 224.760 129.410 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 125.430 224.760 125.730 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.070 224.760 118.370 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 114.390 224.760 114.690 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.030 224.760 107.330 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 103.350 224.760 103.650 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 95.990 224.760 96.290 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 92.310 224.760 92.610 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 9.526400 ;
    PORT
      LAYER met4 ;
        RECT 29.750 224.760 30.050 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 9.526400 ;
    PORT
      LAYER met4 ;
        RECT 26.070 224.760 26.370 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 9.526400 ;
    PORT
      LAYER met4 ;
        RECT 22.390 224.760 22.690 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 9.526400 ;
    PORT
      LAYER met4 ;
        RECT 18.710 224.760 19.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 9.526400 ;
    PORT
      LAYER met4 ;
        RECT 15.030 224.760 15.330 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 9.526400 ;
    PORT
      LAYER met4 ;
        RECT 11.350 224.760 11.650 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 9.526400 ;
    PORT
      LAYER met4 ;
        RECT 7.670 224.760 7.970 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 9.526400 ;
    PORT
      LAYER met4 ;
        RECT 3.990 224.760 4.290 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 9.526400 ;
    PORT
      LAYER met4 ;
        RECT 59.190 224.760 59.490 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 9.526400 ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 9.526400 ;
    PORT
      LAYER met4 ;
        RECT 51.830 224.760 52.130 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 9.526400 ;
    PORT
      LAYER met4 ;
        RECT 48.150 224.760 48.450 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 9.526400 ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 9.526400 ;
    PORT
      LAYER met4 ;
        RECT 40.790 224.760 41.090 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 9.526400 ;
    PORT
      LAYER met4 ;
        RECT 37.110 224.760 37.410 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 9.526400 ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 9.526400 ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 9.526400 ;
    PORT
      LAYER met4 ;
        RECT 84.950 224.760 85.250 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 9.526400 ;
    PORT
      LAYER met4 ;
        RECT 81.270 224.760 81.570 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 9.526400 ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 9.526400 ;
    PORT
      LAYER met4 ;
        RECT 73.910 224.760 74.210 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 9.526400 ;
    PORT
      LAYER met4 ;
        RECT 70.230 224.760 70.530 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 9.526400 ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 9.526400 ;
    PORT
      LAYER met4 ;
        RECT 62.870 224.760 63.170 225.760 ;
    END
  END uo_out[7]
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 2.500 220.760 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 49.000 5.000 50.500 220.760 ;
    END
  END VGND
  OBS
      LAYER nwell ;
        RECT 102.410 26.970 104.520 30.160 ;
        RECT 106.680 26.920 117.950 30.110 ;
      LAYER pwell ;
        RECT 102.390 22.970 104.500 26.070 ;
        RECT 106.650 22.930 117.920 26.030 ;
      LAYER li1 ;
        RECT 103.150 29.980 103.750 30.020 ;
        RECT 102.590 29.810 104.340 29.980 ;
        RECT 109.070 29.930 114.840 29.970 ;
        RECT 102.590 27.320 102.760 29.810 ;
        RECT 103.150 29.800 103.750 29.810 ;
        RECT 103.300 29.300 103.630 29.470 ;
        RECT 103.160 28.045 103.330 29.085 ;
        RECT 103.600 28.045 103.770 29.085 ;
        RECT 103.300 27.660 103.630 27.830 ;
        RECT 104.170 27.320 104.340 29.810 ;
        RECT 102.590 27.150 104.340 27.320 ;
        RECT 106.860 29.760 117.770 29.930 ;
        RECT 106.860 27.270 107.030 29.760 ;
        RECT 109.070 29.730 114.840 29.760 ;
        RECT 108.070 29.250 108.400 29.420 ;
        RECT 109.030 29.250 109.360 29.420 ;
        RECT 109.990 29.250 110.320 29.420 ;
        RECT 110.950 29.250 111.280 29.420 ;
        RECT 111.910 29.250 112.240 29.420 ;
        RECT 112.870 29.250 113.200 29.420 ;
        RECT 113.830 29.250 114.160 29.420 ;
        RECT 114.790 29.250 115.120 29.420 ;
        RECT 115.750 29.250 116.080 29.420 ;
        RECT 116.710 29.250 117.040 29.420 ;
        RECT 107.430 27.995 107.600 29.035 ;
        RECT 107.910 27.995 108.080 29.035 ;
        RECT 108.390 27.995 108.560 29.035 ;
        RECT 108.870 27.995 109.040 29.035 ;
        RECT 109.350 27.995 109.520 29.035 ;
        RECT 109.830 27.995 110.000 29.035 ;
        RECT 110.310 27.995 110.480 29.035 ;
        RECT 110.790 27.995 110.960 29.035 ;
        RECT 111.270 27.995 111.440 29.035 ;
        RECT 111.750 27.995 111.920 29.035 ;
        RECT 112.230 27.995 112.400 29.035 ;
        RECT 112.710 27.995 112.880 29.035 ;
        RECT 113.190 27.995 113.360 29.035 ;
        RECT 113.670 27.995 113.840 29.035 ;
        RECT 114.150 27.995 114.320 29.035 ;
        RECT 114.630 27.995 114.800 29.035 ;
        RECT 115.110 27.995 115.280 29.035 ;
        RECT 115.590 27.995 115.760 29.035 ;
        RECT 116.070 27.995 116.240 29.035 ;
        RECT 116.550 27.995 116.720 29.035 ;
        RECT 117.030 27.995 117.200 29.035 ;
        RECT 107.590 27.610 107.920 27.780 ;
        RECT 108.550 27.610 108.880 27.780 ;
        RECT 109.510 27.610 109.840 27.780 ;
        RECT 110.470 27.610 110.800 27.780 ;
        RECT 111.430 27.610 111.760 27.780 ;
        RECT 112.390 27.610 112.720 27.780 ;
        RECT 113.350 27.610 113.680 27.780 ;
        RECT 114.310 27.610 114.640 27.780 ;
        RECT 115.270 27.610 115.600 27.780 ;
        RECT 116.230 27.610 116.560 27.780 ;
        RECT 117.600 27.270 117.770 29.760 ;
        RECT 106.860 27.100 117.770 27.270 ;
        RECT 102.570 25.720 104.320 25.890 ;
        RECT 102.570 23.320 102.740 25.720 ;
        RECT 103.280 25.210 103.610 25.380 ;
        RECT 103.140 24.000 103.310 25.040 ;
        RECT 103.580 24.000 103.750 25.040 ;
        RECT 103.280 23.660 103.610 23.830 ;
        RECT 103.180 23.320 103.730 23.340 ;
        RECT 104.150 23.320 104.320 25.720 ;
        RECT 102.570 23.150 104.320 23.320 ;
        RECT 106.830 25.680 117.740 25.850 ;
        RECT 106.830 23.280 107.000 25.680 ;
        RECT 108.040 25.170 108.370 25.340 ;
        RECT 109.000 25.170 109.330 25.340 ;
        RECT 109.960 25.170 110.290 25.340 ;
        RECT 110.920 25.170 111.250 25.340 ;
        RECT 111.880 25.170 112.210 25.340 ;
        RECT 112.840 25.170 113.170 25.340 ;
        RECT 113.800 25.170 114.130 25.340 ;
        RECT 114.760 25.170 115.090 25.340 ;
        RECT 115.720 25.170 116.050 25.340 ;
        RECT 116.680 25.170 117.010 25.340 ;
        RECT 107.400 23.960 107.570 25.000 ;
        RECT 107.880 23.960 108.050 25.000 ;
        RECT 108.360 23.960 108.530 25.000 ;
        RECT 108.840 23.960 109.010 25.000 ;
        RECT 109.320 23.960 109.490 25.000 ;
        RECT 109.800 23.960 109.970 25.000 ;
        RECT 110.280 23.960 110.450 25.000 ;
        RECT 110.760 23.960 110.930 25.000 ;
        RECT 111.240 23.960 111.410 25.000 ;
        RECT 111.720 23.960 111.890 25.000 ;
        RECT 112.200 23.960 112.370 25.000 ;
        RECT 112.680 23.960 112.850 25.000 ;
        RECT 113.160 23.960 113.330 25.000 ;
        RECT 113.640 23.960 113.810 25.000 ;
        RECT 114.120 23.960 114.290 25.000 ;
        RECT 114.600 23.960 114.770 25.000 ;
        RECT 115.080 23.960 115.250 25.000 ;
        RECT 115.560 23.960 115.730 25.000 ;
        RECT 116.040 23.960 116.210 25.000 ;
        RECT 116.520 23.960 116.690 25.000 ;
        RECT 117.000 23.960 117.170 25.000 ;
        RECT 107.560 23.620 107.890 23.790 ;
        RECT 108.520 23.620 108.850 23.790 ;
        RECT 109.480 23.620 109.810 23.790 ;
        RECT 110.440 23.620 110.770 23.790 ;
        RECT 111.400 23.620 111.730 23.790 ;
        RECT 112.360 23.620 112.690 23.790 ;
        RECT 113.320 23.620 113.650 23.790 ;
        RECT 114.280 23.620 114.610 23.790 ;
        RECT 115.240 23.620 115.570 23.790 ;
        RECT 116.200 23.620 116.530 23.790 ;
        RECT 109.200 23.280 114.880 23.310 ;
        RECT 117.570 23.280 117.740 25.680 ;
        RECT 103.180 23.130 103.730 23.150 ;
        RECT 106.830 23.110 117.740 23.280 ;
        RECT 109.200 23.050 114.880 23.110 ;
      LAYER mcon ;
        RECT 103.380 29.300 103.550 29.470 ;
        RECT 103.160 28.125 103.330 29.005 ;
        RECT 103.600 28.125 103.770 29.005 ;
        RECT 103.380 27.660 103.550 27.830 ;
        RECT 108.150 29.250 108.320 29.420 ;
        RECT 109.110 29.250 109.280 29.420 ;
        RECT 110.070 29.250 110.240 29.420 ;
        RECT 111.030 29.250 111.200 29.420 ;
        RECT 111.990 29.250 112.160 29.420 ;
        RECT 112.950 29.250 113.120 29.420 ;
        RECT 113.910 29.250 114.080 29.420 ;
        RECT 114.870 29.250 115.040 29.420 ;
        RECT 115.830 29.250 116.000 29.420 ;
        RECT 116.790 29.250 116.960 29.420 ;
        RECT 107.430 28.075 107.600 28.955 ;
        RECT 107.910 28.075 108.080 28.955 ;
        RECT 108.390 28.075 108.560 28.955 ;
        RECT 108.870 28.075 109.040 28.955 ;
        RECT 109.350 28.075 109.520 28.955 ;
        RECT 109.830 28.075 110.000 28.955 ;
        RECT 110.310 28.075 110.480 28.955 ;
        RECT 110.790 28.075 110.960 28.955 ;
        RECT 111.270 28.075 111.440 28.955 ;
        RECT 111.750 28.075 111.920 28.955 ;
        RECT 112.230 28.075 112.400 28.955 ;
        RECT 112.710 28.075 112.880 28.955 ;
        RECT 113.190 28.075 113.360 28.955 ;
        RECT 113.670 28.075 113.840 28.955 ;
        RECT 114.150 28.075 114.320 28.955 ;
        RECT 114.630 28.075 114.800 28.955 ;
        RECT 115.110 28.075 115.280 28.955 ;
        RECT 115.590 28.075 115.760 28.955 ;
        RECT 116.070 28.075 116.240 28.955 ;
        RECT 116.550 28.075 116.720 28.955 ;
        RECT 117.030 28.075 117.200 28.955 ;
        RECT 107.670 27.610 107.840 27.780 ;
        RECT 108.630 27.610 108.800 27.780 ;
        RECT 109.590 27.610 109.760 27.780 ;
        RECT 110.550 27.610 110.720 27.780 ;
        RECT 111.510 27.610 111.680 27.780 ;
        RECT 112.470 27.610 112.640 27.780 ;
        RECT 113.430 27.610 113.600 27.780 ;
        RECT 114.390 27.610 114.560 27.780 ;
        RECT 115.350 27.610 115.520 27.780 ;
        RECT 116.310 27.610 116.480 27.780 ;
        RECT 103.360 25.210 103.530 25.380 ;
        RECT 103.140 24.080 103.310 24.960 ;
        RECT 103.580 24.080 103.750 24.960 ;
        RECT 103.360 23.660 103.530 23.830 ;
        RECT 108.120 25.170 108.290 25.340 ;
        RECT 109.080 25.170 109.250 25.340 ;
        RECT 110.040 25.170 110.210 25.340 ;
        RECT 111.000 25.170 111.170 25.340 ;
        RECT 111.960 25.170 112.130 25.340 ;
        RECT 112.920 25.170 113.090 25.340 ;
        RECT 113.880 25.170 114.050 25.340 ;
        RECT 114.840 25.170 115.010 25.340 ;
        RECT 115.800 25.170 115.970 25.340 ;
        RECT 116.760 25.170 116.930 25.340 ;
        RECT 107.400 24.040 107.570 24.920 ;
        RECT 107.880 24.040 108.050 24.920 ;
        RECT 108.360 24.040 108.530 24.920 ;
        RECT 108.840 24.040 109.010 24.920 ;
        RECT 109.320 24.040 109.490 24.920 ;
        RECT 109.800 24.040 109.970 24.920 ;
        RECT 110.280 24.040 110.450 24.920 ;
        RECT 110.760 24.040 110.930 24.920 ;
        RECT 111.240 24.040 111.410 24.920 ;
        RECT 111.720 24.040 111.890 24.920 ;
        RECT 112.200 24.040 112.370 24.920 ;
        RECT 112.680 24.040 112.850 24.920 ;
        RECT 113.160 24.040 113.330 24.920 ;
        RECT 113.640 24.040 113.810 24.920 ;
        RECT 114.120 24.040 114.290 24.920 ;
        RECT 114.600 24.040 114.770 24.920 ;
        RECT 115.080 24.040 115.250 24.920 ;
        RECT 115.560 24.040 115.730 24.920 ;
        RECT 116.040 24.040 116.210 24.920 ;
        RECT 116.520 24.040 116.690 24.920 ;
        RECT 117.000 24.040 117.170 24.920 ;
        RECT 107.640 23.620 107.810 23.790 ;
        RECT 108.600 23.620 108.770 23.790 ;
        RECT 109.560 23.620 109.730 23.790 ;
        RECT 110.520 23.620 110.690 23.790 ;
        RECT 111.480 23.620 111.650 23.790 ;
        RECT 112.440 23.620 112.610 23.790 ;
        RECT 113.400 23.620 113.570 23.790 ;
        RECT 114.360 23.620 114.530 23.790 ;
        RECT 115.320 23.620 115.490 23.790 ;
        RECT 116.280 23.620 116.450 23.790 ;
      LAYER met1 ;
        RECT 92.840 32.180 94.340 32.210 ;
        RECT 97.350 32.180 120.420 32.320 ;
        RECT 92.840 30.820 120.420 32.180 ;
        RECT 92.840 30.700 99.350 30.820 ;
        RECT 92.840 30.680 99.340 30.700 ;
        RECT 92.840 30.650 94.340 30.680 ;
        RECT 101.700 28.970 102.190 30.820 ;
        RECT 103.030 29.710 103.860 30.820 ;
        RECT 106.030 30.560 106.390 30.820 ;
        RECT 106.000 30.200 106.420 30.560 ;
        RECT 108.990 30.250 114.990 30.820 ;
        RECT 108.980 29.700 114.990 30.250 ;
        RECT 104.585 29.530 105.830 29.535 ;
        RECT 103.270 29.285 105.830 29.530 ;
        RECT 103.270 29.280 104.840 29.285 ;
        RECT 103.320 29.270 103.610 29.280 ;
        RECT 103.130 28.970 103.360 29.065 ;
        RECT 101.700 28.260 103.360 28.970 ;
        RECT 102.130 28.200 103.360 28.260 ;
        RECT 103.130 28.065 103.360 28.200 ;
        RECT 103.570 28.830 103.800 29.065 ;
        RECT 103.570 28.430 105.290 28.830 ;
        RECT 103.570 28.065 103.800 28.430 ;
        RECT 105.585 27.885 105.830 29.285 ;
        RECT 103.285 27.635 105.830 27.885 ;
        RECT 106.300 29.255 117.275 29.505 ;
        RECT 106.300 27.825 106.550 29.255 ;
        RECT 108.090 29.220 108.380 29.255 ;
        RECT 109.050 29.220 109.340 29.255 ;
        RECT 110.010 29.220 110.300 29.255 ;
        RECT 110.970 29.220 111.260 29.255 ;
        RECT 111.930 29.220 112.220 29.255 ;
        RECT 112.890 29.220 113.180 29.255 ;
        RECT 113.850 29.220 114.140 29.255 ;
        RECT 114.810 29.220 115.100 29.255 ;
        RECT 115.770 29.220 116.060 29.255 ;
        RECT 116.730 29.220 117.020 29.255 ;
        RECT 107.400 28.980 107.630 29.015 ;
        RECT 107.340 28.690 107.720 28.980 ;
        RECT 107.400 28.015 107.630 28.690 ;
        RECT 107.880 28.350 108.110 29.015 ;
        RECT 108.360 29.000 108.590 29.015 ;
        RECT 108.300 28.710 108.680 29.000 ;
        RECT 107.820 28.080 108.180 28.350 ;
        RECT 107.880 28.015 108.110 28.080 ;
        RECT 108.360 28.015 108.590 28.710 ;
        RECT 108.840 28.370 109.070 29.015 ;
        RECT 109.320 29.010 109.550 29.015 ;
        RECT 109.230 28.700 109.600 29.010 ;
        RECT 108.780 28.100 109.140 28.370 ;
        RECT 108.840 28.015 109.070 28.100 ;
        RECT 109.320 28.015 109.550 28.700 ;
        RECT 109.800 28.350 110.030 29.015 ;
        RECT 110.280 28.990 110.510 29.015 ;
        RECT 110.240 28.680 110.610 28.990 ;
        RECT 109.730 28.080 110.090 28.350 ;
        RECT 109.800 28.015 110.030 28.080 ;
        RECT 110.280 28.015 110.510 28.680 ;
        RECT 110.760 28.330 110.990 29.015 ;
        RECT 111.240 28.990 111.470 29.015 ;
        RECT 111.180 28.680 111.550 28.990 ;
        RECT 110.670 28.060 111.030 28.330 ;
        RECT 110.760 28.015 110.990 28.060 ;
        RECT 111.240 28.015 111.470 28.680 ;
        RECT 111.720 28.360 111.950 29.015 ;
        RECT 112.200 29.010 112.430 29.015 ;
        RECT 112.160 28.700 112.530 29.010 ;
        RECT 111.650 28.090 112.010 28.360 ;
        RECT 111.720 28.015 111.950 28.090 ;
        RECT 112.200 28.015 112.430 28.700 ;
        RECT 112.680 28.340 112.910 29.015 ;
        RECT 113.080 28.710 113.450 29.020 ;
        RECT 112.620 28.070 112.980 28.340 ;
        RECT 112.680 28.015 112.910 28.070 ;
        RECT 113.160 28.015 113.390 28.710 ;
        RECT 113.640 28.320 113.870 29.015 ;
        RECT 114.120 28.970 114.350 29.015 ;
        RECT 114.060 28.660 114.430 28.970 ;
        RECT 113.580 28.050 113.940 28.320 ;
        RECT 113.640 28.015 113.870 28.050 ;
        RECT 114.120 28.015 114.350 28.660 ;
        RECT 114.600 28.340 114.830 29.015 ;
        RECT 115.080 28.990 115.310 29.015 ;
        RECT 115.020 28.680 115.390 28.990 ;
        RECT 114.560 28.070 114.920 28.340 ;
        RECT 114.600 28.015 114.830 28.070 ;
        RECT 115.080 28.015 115.310 28.680 ;
        RECT 115.560 28.340 115.790 29.015 ;
        RECT 115.980 28.710 116.350 29.020 ;
        RECT 115.520 28.070 115.880 28.340 ;
        RECT 115.560 28.015 115.790 28.070 ;
        RECT 116.040 28.015 116.270 28.710 ;
        RECT 116.520 28.340 116.750 29.015 ;
        RECT 116.940 28.710 117.310 29.020 ;
        RECT 116.440 28.070 116.800 28.340 ;
        RECT 116.520 28.015 116.750 28.070 ;
        RECT 117.000 28.015 117.230 28.710 ;
        RECT 106.245 27.745 106.550 27.825 ;
        RECT 107.610 27.745 107.900 27.810 ;
        RECT 108.570 27.745 108.860 27.810 ;
        RECT 109.530 27.745 109.820 27.810 ;
        RECT 110.490 27.745 110.780 27.810 ;
        RECT 111.450 27.745 111.740 27.810 ;
        RECT 112.410 27.745 112.700 27.810 ;
        RECT 113.370 27.745 113.660 27.810 ;
        RECT 114.330 27.745 114.620 27.810 ;
        RECT 115.290 27.745 115.580 27.810 ;
        RECT 116.250 27.745 116.540 27.810 ;
        RECT 103.320 27.630 103.610 27.635 ;
        RECT 98.550 26.685 100.040 27.030 ;
        RECT 105.265 26.685 105.515 27.635 ;
        RECT 106.245 27.495 116.845 27.745 ;
        RECT 106.245 26.760 106.495 27.495 ;
        RECT 119.240 27.110 120.240 27.180 ;
        RECT 119.240 26.890 121.200 27.110 ;
        RECT 98.550 26.435 105.515 26.685 ;
        RECT 98.550 25.690 100.040 26.435 ;
        RECT 98.860 25.330 99.520 25.690 ;
        RECT 103.290 25.400 103.960 25.430 ;
        RECT 105.265 25.400 105.515 26.435 ;
        RECT 106.240 26.300 106.640 26.760 ;
        RECT 118.400 26.510 121.200 26.890 ;
        RECT 118.400 26.360 120.240 26.510 ;
        RECT 106.245 25.400 106.495 26.300 ;
        RECT 119.240 26.180 120.240 26.360 ;
        RECT 120.600 26.270 121.200 26.510 ;
        RECT 134.480 26.270 135.080 26.300 ;
        RECT 120.600 25.670 135.080 26.270 ;
        RECT 134.480 25.640 135.080 25.670 ;
        RECT 103.290 25.210 105.890 25.400 ;
        RECT 103.300 25.180 103.590 25.210 ;
        RECT 103.740 25.170 105.890 25.210 ;
        RECT 104.760 25.150 105.890 25.170 ;
        RECT 106.245 25.160 117.315 25.400 ;
        RECT 106.245 25.150 115.070 25.160 ;
        RECT 115.360 25.150 117.315 25.160 ;
        RECT 103.110 24.970 103.340 25.020 ;
        RECT 102.040 24.870 103.340 24.970 ;
        RECT 101.700 24.200 103.340 24.870 ;
        RECT 101.700 22.340 102.160 24.200 ;
        RECT 103.110 24.020 103.340 24.200 ;
        RECT 103.550 24.720 103.780 25.020 ;
        RECT 103.550 24.320 105.290 24.720 ;
        RECT 103.550 24.020 103.780 24.320 ;
        RECT 103.300 23.835 103.590 23.860 ;
        RECT 105.635 23.835 105.885 25.150 ;
        RECT 106.245 23.835 106.495 25.150 ;
        RECT 108.060 25.140 108.350 25.150 ;
        RECT 109.020 25.140 109.310 25.150 ;
        RECT 109.980 25.140 110.270 25.150 ;
        RECT 110.940 25.140 111.230 25.150 ;
        RECT 111.900 25.140 112.190 25.150 ;
        RECT 112.860 25.140 113.150 25.150 ;
        RECT 113.820 25.140 114.110 25.150 ;
        RECT 114.780 25.140 115.070 25.150 ;
        RECT 115.740 25.140 116.030 25.150 ;
        RECT 116.700 25.140 116.990 25.150 ;
        RECT 107.370 24.950 107.600 24.980 ;
        RECT 107.310 24.660 107.690 24.950 ;
        RECT 107.370 23.980 107.600 24.660 ;
        RECT 107.850 24.320 108.080 24.980 ;
        RECT 108.330 24.970 108.560 24.980 ;
        RECT 108.270 24.680 108.650 24.970 ;
        RECT 107.790 24.050 108.150 24.320 ;
        RECT 107.850 23.980 108.080 24.050 ;
        RECT 108.330 23.980 108.560 24.680 ;
        RECT 108.810 24.340 109.040 24.980 ;
        RECT 109.200 24.670 109.570 24.980 ;
        RECT 108.750 24.070 109.110 24.340 ;
        RECT 108.810 23.980 109.040 24.070 ;
        RECT 109.290 23.980 109.520 24.670 ;
        RECT 109.770 24.320 110.000 24.980 ;
        RECT 110.250 24.960 110.480 24.980 ;
        RECT 110.210 24.650 110.580 24.960 ;
        RECT 109.700 24.050 110.060 24.320 ;
        RECT 109.770 23.980 110.000 24.050 ;
        RECT 110.250 23.980 110.480 24.650 ;
        RECT 110.730 24.300 110.960 24.980 ;
        RECT 111.210 24.960 111.440 24.980 ;
        RECT 111.150 24.650 111.520 24.960 ;
        RECT 110.640 24.030 111.000 24.300 ;
        RECT 110.730 23.980 110.960 24.030 ;
        RECT 111.210 23.980 111.440 24.650 ;
        RECT 111.690 24.330 111.920 24.980 ;
        RECT 112.130 24.670 112.500 24.980 ;
        RECT 111.620 24.060 111.980 24.330 ;
        RECT 111.690 23.980 111.920 24.060 ;
        RECT 112.170 23.980 112.400 24.670 ;
        RECT 112.650 24.310 112.880 24.980 ;
        RECT 113.050 24.680 113.420 24.990 ;
        RECT 112.590 24.040 112.950 24.310 ;
        RECT 112.650 23.980 112.880 24.040 ;
        RECT 113.130 23.980 113.360 24.680 ;
        RECT 113.610 24.290 113.840 24.980 ;
        RECT 114.090 24.940 114.320 24.980 ;
        RECT 114.030 24.630 114.400 24.940 ;
        RECT 113.550 24.020 113.910 24.290 ;
        RECT 113.610 23.980 113.840 24.020 ;
        RECT 114.090 23.980 114.320 24.630 ;
        RECT 114.570 24.310 114.800 24.980 ;
        RECT 115.050 24.960 115.280 24.980 ;
        RECT 114.990 24.650 115.360 24.960 ;
        RECT 114.530 24.040 114.890 24.310 ;
        RECT 114.570 23.980 114.800 24.040 ;
        RECT 115.050 23.980 115.280 24.650 ;
        RECT 115.530 24.310 115.760 24.980 ;
        RECT 115.950 24.680 116.320 24.990 ;
        RECT 115.490 24.040 115.850 24.310 ;
        RECT 115.530 23.980 115.760 24.040 ;
        RECT 116.010 23.980 116.240 24.680 ;
        RECT 116.490 24.310 116.720 24.980 ;
        RECT 116.910 24.680 117.280 24.990 ;
        RECT 116.410 24.040 116.770 24.310 ;
        RECT 116.490 23.980 116.720 24.040 ;
        RECT 116.970 23.980 117.200 24.680 ;
        RECT 103.265 23.585 105.890 23.835 ;
        RECT 106.245 23.595 116.915 23.835 ;
        RECT 106.400 23.585 116.915 23.595 ;
        RECT 103.070 23.310 103.830 23.380 ;
        RECT 103.060 22.340 103.830 23.310 ;
        RECT 105.980 22.780 106.400 23.140 ;
        RECT 106.010 22.340 106.370 22.780 ;
        RECT 108.990 22.340 114.990 23.340 ;
        RECT 97.700 22.290 120.770 22.340 ;
        RECT 96.100 21.180 120.770 22.290 ;
        RECT 94.680 20.840 120.770 21.180 ;
        RECT 94.680 20.790 99.360 20.840 ;
        RECT 94.680 19.650 97.600 20.790 ;
        RECT 94.680 19.620 96.180 19.650 ;
      LAYER via ;
        RECT 106.030 30.200 106.390 30.560 ;
        RECT 104.860 28.430 105.260 28.830 ;
        RECT 107.390 28.690 107.670 28.980 ;
        RECT 108.350 28.710 108.630 29.000 ;
        RECT 107.870 28.080 108.130 28.350 ;
        RECT 109.280 28.700 109.550 29.010 ;
        RECT 108.830 28.100 109.090 28.370 ;
        RECT 110.290 28.680 110.560 28.990 ;
        RECT 109.780 28.080 110.040 28.350 ;
        RECT 111.230 28.680 111.500 28.990 ;
        RECT 110.720 28.060 110.980 28.330 ;
        RECT 112.210 28.700 112.480 29.010 ;
        RECT 111.700 28.090 111.960 28.360 ;
        RECT 113.130 28.710 113.400 29.020 ;
        RECT 112.670 28.070 112.930 28.340 ;
        RECT 114.110 28.660 114.380 28.970 ;
        RECT 113.630 28.050 113.890 28.320 ;
        RECT 115.070 28.680 115.340 28.990 ;
        RECT 114.610 28.070 114.870 28.340 ;
        RECT 116.030 28.710 116.300 29.020 ;
        RECT 115.570 28.070 115.830 28.340 ;
        RECT 116.990 28.710 117.260 29.020 ;
        RECT 116.490 28.070 116.750 28.340 ;
        RECT 98.890 25.330 99.490 25.930 ;
        RECT 106.240 26.330 106.640 26.730 ;
        RECT 118.610 26.480 118.870 26.740 ;
        RECT 134.480 25.670 135.080 26.270 ;
        RECT 104.860 24.320 105.260 24.720 ;
        RECT 107.360 24.660 107.640 24.950 ;
        RECT 108.320 24.680 108.600 24.970 ;
        RECT 107.840 24.050 108.100 24.320 ;
        RECT 109.250 24.670 109.520 24.980 ;
        RECT 108.800 24.070 109.060 24.340 ;
        RECT 110.260 24.650 110.530 24.960 ;
        RECT 109.750 24.050 110.010 24.320 ;
        RECT 111.200 24.650 111.470 24.960 ;
        RECT 110.690 24.030 110.950 24.300 ;
        RECT 112.180 24.670 112.450 24.980 ;
        RECT 111.670 24.060 111.930 24.330 ;
        RECT 113.100 24.680 113.370 24.990 ;
        RECT 112.640 24.040 112.900 24.310 ;
        RECT 114.080 24.630 114.350 24.940 ;
        RECT 113.600 24.020 113.860 24.290 ;
        RECT 115.040 24.650 115.310 24.960 ;
        RECT 114.580 24.040 114.840 24.310 ;
        RECT 116.000 24.680 116.270 24.990 ;
        RECT 115.540 24.040 115.800 24.310 ;
        RECT 116.960 24.680 117.230 24.990 ;
        RECT 116.460 24.040 116.720 24.310 ;
        RECT 106.010 22.780 106.370 23.140 ;
      LAYER met2 ;
        RECT 89.595 32.180 91.045 32.200 ;
        RECT 89.570 30.680 94.370 32.180 ;
        RECT 89.595 30.660 91.045 30.680 ;
        RECT 104.860 26.730 105.260 28.860 ;
        RECT 106.030 28.400 106.390 30.590 ;
        RECT 107.390 28.980 107.670 29.030 ;
        RECT 108.350 28.980 108.630 29.050 ;
        RECT 109.280 28.980 109.550 29.060 ;
        RECT 110.290 28.980 110.560 29.040 ;
        RECT 111.230 28.980 111.500 29.040 ;
        RECT 112.210 28.980 112.480 29.060 ;
        RECT 113.130 28.980 113.400 29.070 ;
        RECT 114.110 28.980 114.380 29.020 ;
        RECT 115.070 28.980 115.340 29.040 ;
        RECT 116.030 28.980 116.300 29.070 ;
        RECT 116.990 28.980 117.260 29.070 ;
        RECT 107.340 28.720 118.870 28.980 ;
        RECT 107.390 28.640 107.670 28.720 ;
        RECT 108.350 28.660 108.630 28.720 ;
        RECT 109.280 28.650 109.550 28.720 ;
        RECT 110.290 28.630 110.560 28.720 ;
        RECT 111.230 28.630 111.500 28.720 ;
        RECT 112.210 28.650 112.480 28.720 ;
        RECT 113.130 28.660 113.400 28.720 ;
        RECT 114.110 28.610 114.380 28.720 ;
        RECT 115.070 28.630 115.340 28.720 ;
        RECT 116.030 28.660 116.300 28.720 ;
        RECT 116.990 28.660 117.260 28.720 ;
        RECT 108.830 28.400 109.090 28.420 ;
        RECT 111.700 28.400 111.960 28.410 ;
        RECT 106.030 28.040 118.010 28.400 ;
        RECT 107.870 28.030 108.130 28.040 ;
        RECT 109.780 28.030 110.040 28.040 ;
        RECT 110.720 28.010 110.980 28.040 ;
        RECT 112.670 28.020 112.930 28.040 ;
        RECT 113.630 28.000 113.890 28.040 ;
        RECT 114.610 28.020 114.870 28.040 ;
        RECT 115.570 28.020 115.830 28.040 ;
        RECT 116.490 28.020 116.750 28.040 ;
        RECT 118.610 27.080 118.870 28.720 ;
        RECT 104.860 26.330 106.670 26.730 ;
        RECT 98.890 25.175 99.490 25.960 ;
        RECT 98.870 24.625 99.510 25.175 ;
        RECT 98.890 24.600 99.490 24.625 ;
        RECT 104.860 24.290 105.260 26.330 ;
        RECT 118.500 26.115 118.970 27.080 ;
        RECT 118.500 25.980 119.125 26.115 ;
        RECT 118.610 25.530 119.125 25.980 ;
        RECT 134.450 25.670 135.110 26.270 ;
        RECT 107.360 24.950 107.640 25.000 ;
        RECT 108.320 24.950 108.600 25.020 ;
        RECT 109.250 24.950 109.520 25.030 ;
        RECT 110.260 24.950 110.530 25.010 ;
        RECT 111.200 24.950 111.470 25.010 ;
        RECT 112.180 24.950 112.450 25.030 ;
        RECT 113.100 24.950 113.370 25.040 ;
        RECT 114.080 24.950 114.350 24.990 ;
        RECT 115.040 24.950 115.310 25.010 ;
        RECT 116.000 24.950 116.270 25.040 ;
        RECT 116.960 24.950 117.230 25.040 ;
        RECT 118.560 24.950 119.125 25.530 ;
        RECT 107.310 24.690 119.125 24.950 ;
        RECT 107.360 24.610 107.640 24.690 ;
        RECT 108.320 24.630 108.600 24.690 ;
        RECT 109.250 24.620 109.520 24.690 ;
        RECT 110.260 24.600 110.530 24.690 ;
        RECT 111.200 24.600 111.470 24.690 ;
        RECT 112.180 24.620 112.450 24.690 ;
        RECT 113.100 24.630 113.370 24.690 ;
        RECT 114.080 24.580 114.350 24.690 ;
        RECT 115.040 24.600 115.310 24.690 ;
        RECT 116.000 24.630 116.270 24.690 ;
        RECT 116.960 24.630 117.230 24.690 ;
        RECT 118.560 24.495 119.125 24.690 ;
        RECT 118.560 24.470 118.820 24.495 ;
        RECT 108.800 24.370 109.060 24.390 ;
        RECT 111.670 24.370 111.930 24.380 ;
        RECT 106.010 24.010 117.980 24.370 ;
        RECT 106.010 22.750 106.370 24.010 ;
        RECT 107.840 24.000 108.100 24.010 ;
        RECT 109.750 24.000 110.010 24.010 ;
        RECT 110.690 23.980 110.950 24.010 ;
        RECT 112.640 23.990 112.900 24.010 ;
        RECT 113.600 23.970 113.860 24.010 ;
        RECT 114.580 23.990 114.840 24.010 ;
        RECT 115.540 23.990 115.800 24.010 ;
        RECT 116.460 23.990 116.720 24.010 ;
        RECT 134.480 21.245 135.080 25.670 ;
        RECT 93.375 21.150 94.825 21.170 ;
        RECT 93.350 19.650 96.210 21.150 ;
        RECT 134.460 20.695 135.100 21.245 ;
        RECT 134.480 20.670 135.080 20.695 ;
        RECT 93.375 19.630 94.825 19.650 ;
      LAYER via2 ;
        RECT 89.595 30.705 91.045 32.155 ;
        RECT 98.915 24.625 99.465 25.175 ;
        RECT 93.375 19.675 94.825 21.125 ;
        RECT 134.505 20.695 135.055 21.245 ;
      LAYER met3 ;
        RECT 32.815 32.180 34.305 32.205 ;
        RECT 32.810 30.680 91.070 32.180 ;
        RECT 32.815 30.655 34.305 30.680 ;
        RECT 98.890 23.965 99.490 25.200 ;
        RECT 98.865 23.375 99.515 23.965 ;
        RECT 98.890 23.370 99.490 23.375 ;
        RECT 91.965 21.150 93.455 21.175 ;
        RECT 91.960 19.650 94.850 21.150 ;
        RECT 91.965 19.625 93.455 19.650 ;
        RECT 134.480 8.525 135.080 21.270 ;
        RECT 134.455 7.935 135.105 8.525 ;
        RECT 134.480 7.930 135.080 7.935 ;
      LAYER via3 ;
        RECT 32.815 30.685 34.305 32.175 ;
        RECT 98.895 23.375 99.485 23.965 ;
        RECT 91.965 19.655 93.455 21.145 ;
        RECT 134.485 7.935 135.075 8.525 ;
      LAYER met4 ;
        RECT 3.990 223.300 4.290 224.760 ;
        RECT 7.670 223.300 7.970 224.760 ;
        RECT 11.350 223.300 11.650 224.760 ;
        RECT 15.030 223.300 15.330 224.760 ;
        RECT 18.710 223.300 19.010 224.760 ;
        RECT 22.390 223.300 22.690 224.760 ;
        RECT 26.070 223.300 26.370 224.760 ;
        RECT 29.750 223.300 30.050 224.760 ;
        RECT 33.430 223.300 33.730 224.760 ;
        RECT 37.110 223.300 37.410 224.760 ;
        RECT 40.790 223.300 41.090 224.760 ;
        RECT 44.470 223.300 44.770 224.760 ;
        RECT 48.150 223.300 48.450 224.760 ;
        RECT 51.830 223.300 52.130 224.760 ;
        RECT 55.510 223.300 55.810 224.760 ;
        RECT 59.190 223.300 59.490 224.760 ;
        RECT 62.870 223.300 63.170 224.760 ;
        RECT 66.550 223.300 66.850 224.760 ;
        RECT 70.230 223.300 70.530 224.760 ;
        RECT 73.910 223.300 74.210 224.760 ;
        RECT 77.590 223.300 77.890 224.760 ;
        RECT 81.270 223.300 81.570 224.760 ;
        RECT 84.950 223.300 85.250 224.760 ;
        RECT 88.630 223.300 88.930 224.760 ;
        RECT 3.710 221.420 88.930 223.300 ;
        RECT 49.000 220.760 50.500 221.420 ;
        RECT 88.630 221.350 88.930 221.420 ;
        RECT 2.500 30.680 34.310 32.180 ;
        RECT 50.500 19.650 93.460 21.150 ;
        RECT 98.890 16.030 99.490 23.970 ;
        RECT 98.890 15.430 157.160 16.030 ;
        RECT 134.480 1.000 135.080 8.530 ;
        RECT 156.560 1.000 157.160 15.430 ;
  END
END tt_um_mattvenn_inverter
END LIBRARY

