VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_psychogenic_wowa
  CLASS BLOCK ;
  FOREIGN tt_um_psychogenic_wowa ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met4 ;
        RECT 154.870 224.760 155.170 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 158.550 224.760 158.850 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 151.190 224.760 151.490 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 3.190000 ;
    PORT
      LAYER met4 ;
        RECT 156.560 0.000 157.160 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.060000 ;
    PORT
      LAYER met4 ;
        RECT 134.480 0.000 135.080 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.250000 ;
    PORT
      LAYER met4 ;
        RECT 112.400 0.000 113.000 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.250000 ;
    ANTENNADIFFAREA 1.160000 ;
    PORT
      LAYER met4 ;
        RECT 90.320 0.000 90.920 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.160000 ;
    PORT
      LAYER met4 ;
        RECT 68.240 0.000 68.840 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.160000 ;
    PORT
      LAYER met4 ;
        RECT 46.160 0.000 46.760 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 24.080 0.000 24.680 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 2.000 0.000 2.600 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met4 ;
        RECT 147.510 224.760 147.810 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 140.150 224.760 140.450 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 136.470 224.760 136.770 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 129.110 224.760 129.410 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 125.430 224.760 125.730 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.070 224.760 118.370 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 114.390 224.760 114.690 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.030 224.760 107.330 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 103.350 224.760 103.650 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 95.990 224.760 96.290 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 92.310 224.760 92.610 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 266.685486 ;
    ANTENNADIFFAREA 347.309570 ;
    PORT
      LAYER met4 ;
        RECT 29.750 224.760 30.050 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 266.685486 ;
    ANTENNADIFFAREA 347.309570 ;
    PORT
      LAYER met4 ;
        RECT 26.070 224.760 26.370 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 266.685486 ;
    ANTENNADIFFAREA 347.309570 ;
    PORT
      LAYER met4 ;
        RECT 22.390 224.760 22.690 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 266.685486 ;
    ANTENNADIFFAREA 347.309570 ;
    PORT
      LAYER met4 ;
        RECT 18.710 224.760 19.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 266.685486 ;
    ANTENNADIFFAREA 347.309570 ;
    PORT
      LAYER met4 ;
        RECT 15.030 224.760 15.330 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 266.685486 ;
    ANTENNADIFFAREA 347.309570 ;
    PORT
      LAYER met4 ;
        RECT 11.350 224.760 11.650 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 266.685486 ;
    ANTENNADIFFAREA 347.309570 ;
    PORT
      LAYER met4 ;
        RECT 7.670 224.760 7.970 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 266.685486 ;
    ANTENNADIFFAREA 347.309570 ;
    PORT
      LAYER met4 ;
        RECT 3.990 224.760 4.290 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met4 ;
        RECT 59.190 224.760 59.490 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 415.520691 ;
    ANTENNADIFFAREA 450.978302 ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 415.520691 ;
    ANTENNADIFFAREA 450.978302 ;
    PORT
      LAYER met4 ;
        RECT 51.830 224.760 52.130 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 415.520691 ;
    ANTENNADIFFAREA 450.978302 ;
    PORT
      LAYER met4 ;
        RECT 48.150 224.760 48.450 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 266.685486 ;
    ANTENNADIFFAREA 347.309570 ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 266.685486 ;
    ANTENNADIFFAREA 347.309570 ;
    PORT
      LAYER met4 ;
        RECT 40.790 224.760 41.090 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 266.685486 ;
    ANTENNADIFFAREA 347.309570 ;
    PORT
      LAYER met4 ;
        RECT 37.110 224.760 37.410 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 266.685486 ;
    ANTENNADIFFAREA 347.309570 ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met4 ;
        RECT 84.950 224.760 85.250 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met4 ;
        RECT 81.270 224.760 81.570 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met4 ;
        RECT 73.910 224.760 74.210 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met4 ;
        RECT 70.230 224.760 70.530 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met4 ;
        RECT 62.870 224.760 63.170 225.760 ;
    END
  END uo_out[7]
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 155.000 7.000 156.500 222.760 ;
    END
  END VPWR
  PIN VGND 
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.700 2.500 221.450 ;
    END
  END VGND 
  OBS
      LAYER li1 ;
        RECT 22.730 14.900 131.700 198.745 ;
      LAYER met1 ;
        RECT 20.500 3.220 157.915 198.900 ;
      LAYER met2 ;
        RECT 5.955 1.960 157.900 223.600 ;
      LAYER met3 ;
        RECT 1.770 0.600 157.900 224.450 ;
      LAYER met4 ;
        RECT 1.000 224.360 3.590 225.750 ;
        RECT 4.690 224.360 7.270 225.750 ;
        RECT 8.370 224.360 10.950 225.750 ;
        RECT 12.050 224.360 14.630 225.750 ;
        RECT 15.730 224.360 18.310 225.750 ;
        RECT 19.410 224.360 21.990 225.750 ;
        RECT 23.090 224.360 25.670 225.750 ;
        RECT 26.770 224.360 29.350 225.750 ;
        RECT 30.450 224.360 33.030 225.750 ;
        RECT 34.130 224.360 36.710 225.750 ;
        RECT 37.810 224.360 40.390 225.750 ;
        RECT 41.490 224.360 44.070 225.750 ;
        RECT 45.170 224.360 47.750 225.750 ;
        RECT 48.850 224.360 51.430 225.750 ;
        RECT 52.530 224.360 55.110 225.750 ;
        RECT 56.210 224.360 58.790 225.750 ;
        RECT 59.890 224.360 62.470 225.750 ;
        RECT 63.570 224.360 66.150 225.750 ;
        RECT 67.250 224.360 69.830 225.750 ;
        RECT 70.930 224.360 73.510 225.750 ;
        RECT 74.610 224.360 77.190 225.750 ;
        RECT 78.290 224.360 80.870 225.750 ;
        RECT 81.970 224.360 84.550 225.750 ;
        RECT 85.650 224.360 88.230 225.750 ;
        RECT 89.330 224.360 91.910 225.750 ;
        RECT 93.010 224.360 95.590 225.750 ;
        RECT 96.690 224.360 99.270 225.750 ;
        RECT 100.370 224.360 102.950 225.750 ;
        RECT 104.050 224.360 106.630 225.750 ;
        RECT 107.730 224.360 110.310 225.750 ;
        RECT 111.410 224.360 113.990 225.750 ;
        RECT 115.090 224.360 117.670 225.750 ;
        RECT 118.770 224.360 121.350 225.750 ;
        RECT 122.450 224.360 125.030 225.750 ;
        RECT 126.130 224.360 128.710 225.750 ;
        RECT 129.810 224.360 132.390 225.750 ;
        RECT 133.490 224.360 136.070 225.750 ;
        RECT 137.170 224.360 139.750 225.750 ;
        RECT 140.850 224.360 143.430 225.750 ;
        RECT 144.530 224.360 147.110 225.750 ;
        RECT 148.210 224.360 150.790 225.750 ;
        RECT 151.890 224.360 154.470 225.750 ;
        RECT 155.570 224.360 158.150 225.750 ;
        RECT 1.000 223.160 158.950 224.360 ;
        RECT 1.000 221.850 154.600 223.160 ;
        RECT 1.000 221.450 2.500 221.850 ;
        RECT 2.900 6.600 154.600 221.850 ;
        RECT 156.900 6.600 158.950 223.160 ;
        RECT 2.900 5.300 158.950 6.600 ;
        RECT 1.000 1.400 158.950 5.300 ;
        RECT 1.000 0.000 1.600 1.400 ;
        RECT 3.000 0.000 23.680 1.400 ;
        RECT 25.080 0.000 45.760 1.400 ;
        RECT 47.160 0.000 67.840 1.400 ;
        RECT 69.240 0.000 89.920 1.400 ;
        RECT 91.320 0.000 112.000 1.400 ;
        RECT 113.400 0.000 134.080 1.400 ;
        RECT 135.480 0.000 156.160 1.400 ;
        RECT 157.560 0.000 158.950 1.400 ;
  END
END tt_um_psychogenic_wowa
END LIBRARY

