VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_nurirfansyah_alits01
  CLASS BLOCK ;
  FOREIGN tt_um_nurirfansyah_alits01 ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 154.870 224.760 155.170 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 158.550 224.760 158.850 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 151.190 224.760 151.490 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.250000 ;
    PORT
      LAYER met4 ;
        RECT 156.560 0.000 157.160 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.500000 ;
    PORT
      LAYER met4 ;
        RECT 134.480 0.000 135.080 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 5.000000 ;
    PORT
      LAYER met4 ;
        RECT 112.400 0.000 113.000 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 90.320 0.000 90.920 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 68.240 0.000 68.840 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 46.160 0.000 46.760 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 24.080 0.000 24.680 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 2.000 0.000 2.600 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 147.510 224.760 147.810 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 140.150 224.760 140.450 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 136.470 224.760 136.770 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 129.110 224.760 129.410 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 125.430 224.760 125.730 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.070 224.760 118.370 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 114.390 224.760 114.690 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.030 224.760 107.330 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 103.350 224.760 103.650 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 95.990 224.760 96.290 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 92.310 224.760 92.610 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 29.750 224.760 30.050 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 26.070 224.760 26.370 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 22.390 224.760 22.690 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 18.710 224.760 19.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 15.030 224.760 15.330 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 11.350 224.760 11.650 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 7.670 224.760 7.970 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 3.990 224.760 4.290 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 59.190 224.760 59.490 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 51.830 224.760 52.130 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 48.150 224.760 48.450 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 40.790 224.760 41.090 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 37.110 224.760 37.410 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 84.950 224.760 85.250 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 81.270 224.760 81.570 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 73.910 224.760 74.210 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 70.230 224.760 70.530 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 62.870 224.760 63.170 225.760 ;
    END
  END uo_out[7]
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 2.500 220.760 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 49.000 5.000 50.500 220.760 ;
    END
  END VGND
  OBS
      LAYER nwell ;
        RECT 119.240 31.340 148.490 33.990 ;
      LAYER li1 ;
        RECT 119.240 34.140 148.490 34.490 ;
        RECT 119.740 31.540 119.940 34.140 ;
        RECT 119.440 30.940 119.990 31.340 ;
        RECT 120.190 30.740 120.390 33.540 ;
        RECT 119.540 30.390 120.390 30.740 ;
        RECT 119.440 29.790 119.990 30.190 ;
        RECT 119.740 28.190 119.940 29.590 ;
        RECT 120.190 28.590 120.390 30.390 ;
        RECT 121.090 30.740 121.290 33.540 ;
        RECT 122.390 31.540 122.590 34.140 ;
        RECT 122.840 31.540 123.040 34.140 ;
        RECT 123.140 30.740 123.540 31.290 ;
        RECT 121.090 30.390 121.890 30.740 ;
        RECT 121.090 28.590 121.290 30.390 ;
        RECT 122.390 30.340 123.540 30.740 ;
        RECT 123.140 29.840 123.540 30.340 ;
        RECT 123.740 30.740 123.940 33.540 ;
        RECT 124.640 31.540 124.840 34.140 ;
        RECT 125.590 31.540 125.790 34.140 ;
        RECT 125.290 30.940 125.840 31.340 ;
        RECT 126.040 30.740 126.240 33.540 ;
        RECT 123.740 30.340 124.740 30.740 ;
        RECT 125.390 30.390 126.240 30.740 ;
        RECT 122.390 28.190 122.590 29.590 ;
        RECT 122.840 28.190 123.040 29.590 ;
        RECT 123.740 28.590 123.940 30.340 ;
        RECT 125.290 29.790 125.840 30.190 ;
        RECT 124.640 28.190 124.840 29.590 ;
        RECT 125.590 28.190 125.790 29.590 ;
        RECT 126.040 28.590 126.240 30.390 ;
        RECT 126.940 30.740 127.140 33.540 ;
        RECT 128.240 31.540 128.440 34.140 ;
        RECT 128.690 31.540 128.890 34.140 ;
        RECT 128.990 30.740 129.390 31.290 ;
        RECT 126.940 30.390 127.740 30.740 ;
        RECT 126.940 28.590 127.140 30.390 ;
        RECT 128.240 30.340 129.390 30.740 ;
        RECT 128.990 29.840 129.390 30.340 ;
        RECT 129.590 30.740 129.790 33.540 ;
        RECT 130.490 31.540 130.690 34.140 ;
        RECT 131.440 31.540 131.640 34.140 ;
        RECT 131.140 30.940 131.690 31.340 ;
        RECT 131.890 30.740 132.090 33.540 ;
        RECT 129.590 30.340 130.590 30.740 ;
        RECT 131.240 30.390 132.090 30.740 ;
        RECT 128.240 28.190 128.440 29.590 ;
        RECT 128.690 28.190 128.890 29.590 ;
        RECT 129.590 28.590 129.790 30.340 ;
        RECT 131.140 29.790 131.690 30.190 ;
        RECT 130.490 28.190 130.690 29.590 ;
        RECT 131.440 28.190 131.640 29.590 ;
        RECT 131.890 28.590 132.090 30.390 ;
        RECT 132.790 30.740 132.990 33.540 ;
        RECT 134.090 31.540 134.290 34.140 ;
        RECT 134.540 31.540 134.740 34.140 ;
        RECT 134.840 30.740 135.240 31.290 ;
        RECT 132.790 30.390 133.590 30.740 ;
        RECT 132.790 28.590 132.990 30.390 ;
        RECT 134.090 30.340 135.240 30.740 ;
        RECT 134.840 29.840 135.240 30.340 ;
        RECT 135.440 30.740 135.640 33.540 ;
        RECT 136.340 31.540 136.540 34.140 ;
        RECT 137.290 31.540 137.490 34.140 ;
        RECT 136.990 30.940 137.540 31.340 ;
        RECT 137.740 30.740 137.940 33.540 ;
        RECT 135.440 30.340 136.440 30.740 ;
        RECT 137.090 30.390 137.940 30.740 ;
        RECT 134.090 28.190 134.290 29.590 ;
        RECT 134.540 28.190 134.740 29.590 ;
        RECT 135.440 28.590 135.640 30.340 ;
        RECT 136.990 29.790 137.540 30.190 ;
        RECT 136.340 28.190 136.540 29.590 ;
        RECT 137.290 28.190 137.490 29.590 ;
        RECT 137.740 28.590 137.940 30.390 ;
        RECT 138.640 30.740 138.840 33.540 ;
        RECT 139.940 31.540 140.140 34.140 ;
        RECT 140.390 31.540 140.590 34.140 ;
        RECT 140.690 30.740 141.090 31.290 ;
        RECT 138.640 30.390 139.440 30.740 ;
        RECT 138.640 28.590 138.840 30.390 ;
        RECT 139.940 30.340 141.090 30.740 ;
        RECT 140.690 29.840 141.090 30.340 ;
        RECT 141.290 30.740 141.490 33.540 ;
        RECT 142.190 31.540 142.390 34.140 ;
        RECT 143.140 31.540 143.340 34.140 ;
        RECT 142.840 30.940 143.390 31.340 ;
        RECT 143.590 30.740 143.790 33.540 ;
        RECT 141.290 30.340 142.290 30.740 ;
        RECT 142.940 30.390 143.790 30.740 ;
        RECT 139.940 28.190 140.140 29.590 ;
        RECT 140.390 28.190 140.590 29.590 ;
        RECT 141.290 28.590 141.490 30.340 ;
        RECT 142.840 29.790 143.390 30.190 ;
        RECT 142.190 28.190 142.390 29.590 ;
        RECT 143.140 28.190 143.340 29.590 ;
        RECT 143.590 28.590 143.790 30.390 ;
        RECT 144.490 30.740 144.690 33.540 ;
        RECT 145.790 31.540 145.990 34.140 ;
        RECT 146.240 31.540 146.440 34.140 ;
        RECT 146.540 30.740 146.940 31.290 ;
        RECT 144.490 30.390 145.290 30.740 ;
        RECT 144.490 28.590 144.690 30.390 ;
        RECT 145.790 30.340 146.940 30.740 ;
        RECT 146.540 29.840 146.940 30.340 ;
        RECT 147.140 30.740 147.340 33.540 ;
        RECT 148.040 31.540 148.240 34.140 ;
        RECT 147.140 30.340 148.140 30.740 ;
        RECT 145.790 28.190 145.990 29.590 ;
        RECT 146.240 28.190 146.440 29.590 ;
        RECT 147.140 28.590 147.340 30.340 ;
        RECT 148.040 28.190 148.240 29.590 ;
        RECT 119.240 27.840 148.490 28.190 ;
      LAYER met1 ;
        RECT 0.950 34.540 145.800 34.850 ;
        RECT 0.950 34.150 148.490 34.540 ;
        RECT 119.240 34.090 148.490 34.150 ;
        RECT 119.390 31.290 120.040 31.790 ;
        RECT 125.240 31.290 125.890 31.790 ;
        RECT 131.090 31.290 131.740 31.790 ;
        RECT 136.940 31.290 137.590 31.790 ;
        RECT 142.790 31.290 143.440 31.790 ;
        RECT 119.440 30.940 119.990 31.290 ;
        RECT 125.290 30.940 125.840 31.290 ;
        RECT 131.140 30.940 131.690 31.290 ;
        RECT 136.990 30.940 137.540 31.290 ;
        RECT 142.840 30.940 143.390 31.290 ;
        RECT 118.690 30.740 119.240 30.840 ;
        RECT 121.890 30.740 122.940 30.840 ;
        RECT 118.690 30.390 120.190 30.740 ;
        RECT 121.240 30.390 122.940 30.740 ;
        RECT 118.690 30.290 119.240 30.390 ;
        RECT 121.890 30.240 122.940 30.390 ;
        RECT 124.190 30.740 124.790 30.840 ;
        RECT 127.740 30.740 128.790 30.840 ;
        RECT 124.190 30.390 126.040 30.740 ;
        RECT 127.090 30.390 128.790 30.740 ;
        RECT 124.190 30.240 124.790 30.390 ;
        RECT 127.740 30.240 128.790 30.390 ;
        RECT 130.040 30.240 130.640 30.840 ;
        RECT 133.590 30.740 134.640 30.840 ;
        RECT 131.240 30.390 131.890 30.740 ;
        RECT 132.940 30.390 134.640 30.740 ;
        RECT 133.590 30.240 134.640 30.390 ;
        RECT 135.890 30.740 136.490 30.840 ;
        RECT 139.440 30.740 140.490 30.840 ;
        RECT 135.890 30.390 137.740 30.740 ;
        RECT 138.790 30.390 140.490 30.740 ;
        RECT 135.890 30.240 136.490 30.390 ;
        RECT 139.440 30.240 140.490 30.390 ;
        RECT 141.740 30.740 142.340 30.840 ;
        RECT 145.290 30.740 146.340 30.840 ;
        RECT 141.740 30.390 143.590 30.740 ;
        RECT 144.640 30.390 146.340 30.740 ;
        RECT 141.740 30.240 142.340 30.390 ;
        RECT 145.290 30.240 146.340 30.390 ;
        RECT 147.590 30.240 148.190 30.840 ;
        RECT 119.440 29.790 119.990 30.190 ;
        RECT 125.290 29.790 125.840 30.190 ;
        RECT 131.140 29.790 131.690 30.190 ;
        RECT 136.990 29.790 137.540 30.190 ;
        RECT 142.840 29.790 143.390 30.190 ;
        RECT 119.390 29.290 120.040 29.790 ;
        RECT 125.240 29.290 125.890 29.790 ;
        RECT 131.090 29.290 131.740 29.790 ;
        RECT 136.940 29.290 137.590 29.790 ;
        RECT 142.790 29.290 143.440 29.790 ;
        RECT 119.240 28.200 148.490 28.240 ;
        RECT 48.600 27.300 148.500 28.200 ;
      LAYER met2 ;
        RECT 0.950 34.850 2.550 35.550 ;
        RECT 0.950 34.150 4.850 34.850 ;
        RECT 0.950 33.500 2.550 34.150 ;
        RECT 112.050 31.790 119.400 31.800 ;
        RECT 112.050 31.690 120.040 31.790 ;
        RECT 125.240 31.690 125.890 31.790 ;
        RECT 131.090 31.690 131.740 31.790 ;
        RECT 136.940 31.690 137.590 31.790 ;
        RECT 142.790 31.690 143.440 31.790 ;
        RECT 112.050 31.340 147.840 31.690 ;
        RECT 112.050 31.300 120.040 31.340 ;
        RECT 48.600 28.200 50.750 31.300 ;
        RECT 112.050 30.850 113.300 31.300 ;
        RECT 119.390 31.290 120.040 31.300 ;
        RECT 125.240 31.290 125.890 31.340 ;
        RECT 131.090 31.290 131.740 31.340 ;
        RECT 136.940 31.290 137.590 31.340 ;
        RECT 142.790 31.290 143.440 31.340 ;
        RECT 148.200 30.840 157.200 30.850 ;
        RECT 118.690 30.740 119.240 30.840 ;
        RECT 147.590 30.740 157.200 30.840 ;
        RECT 118.690 30.390 157.200 30.740 ;
        RECT 118.690 30.290 119.240 30.390 ;
        RECT 147.590 30.250 157.200 30.390 ;
        RECT 147.590 30.240 148.340 30.250 ;
        RECT 115.600 29.640 120.050 29.800 ;
        RECT 125.240 29.640 125.890 29.790 ;
        RECT 131.090 29.640 131.740 29.790 ;
        RECT 136.940 29.640 137.590 29.790 ;
        RECT 142.790 29.640 143.440 29.790 ;
        RECT 156.250 29.700 157.200 30.250 ;
        RECT 115.600 29.300 143.440 29.640 ;
        RECT 115.600 28.900 116.850 29.300 ;
        RECT 119.390 29.290 143.440 29.300 ;
        RECT 48.600 27.300 57.600 28.200 ;
        RECT 48.600 25.300 50.750 27.300 ;
      LAYER met3 ;
        RECT 1.000 33.350 2.500 35.700 ;
        RECT 48.900 25.150 50.600 31.350 ;
        RECT 112.250 1.550 113.100 31.700 ;
        RECT 115.850 12.950 116.700 29.850 ;
        RECT 115.850 12.150 135.100 12.950 ;
        RECT 134.350 2.900 135.100 12.150 ;
        RECT 156.450 3.100 157.100 31.000 ;
        RECT 134.350 1.550 135.200 2.900 ;
        RECT 156.450 1.650 157.300 3.100 ;
      LAYER met4 ;
        RECT 112.250 1.550 113.100 2.750 ;
        RECT 134.350 1.550 135.200 2.750 ;
        RECT 156.450 1.650 157.300 2.850 ;
        RECT 112.400 1.000 113.000 1.550 ;
        RECT 134.480 1.000 135.080 1.550 ;
        RECT 156.560 1.000 157.160 1.650 ;
  END
END tt_um_nurirfansyah_alits01
END LIBRARY

