VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_calculator_muehlbb
  CLASS BLOCK ;
  FOREIGN tt_um_calculator_muehlbb ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 111.520 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 40.830 2.480 42.430 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 79.700 2.480 81.300 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 118.570 2.480 120.170 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 157.440 2.480 159.040 109.040 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.395 2.480 22.995 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 60.265 2.480 61.865 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 99.135 2.480 100.735 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 138.005 2.480 139.605 109.040 ;
    END
  END VPWR
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met4 ;
        RECT 154.870 110.520 155.170 111.520 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 158.550 110.520 158.850 111.520 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met4 ;
        RECT 151.190 110.520 151.490 111.520 ;
    END
  END rst_n
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 147.510 110.520 147.810 111.520 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 143.830 110.520 144.130 111.520 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 140.150 110.520 140.450 111.520 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 136.470 110.520 136.770 111.520 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.790 110.520 133.090 111.520 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 129.110 110.520 129.410 111.520 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 125.430 110.520 125.730 111.520 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 121.750 110.520 122.050 111.520 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met4 ;
        RECT 118.070 110.520 118.370 111.520 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met4 ;
        RECT 114.390 110.520 114.690 111.520 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met4 ;
        RECT 110.710 110.520 111.010 111.520 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met4 ;
        RECT 107.030 110.520 107.330 111.520 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 103.350 110.520 103.650 111.520 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 99.670 110.520 99.970 111.520 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 95.990 110.520 96.290 111.520 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met4 ;
        RECT 92.310 110.520 92.610 111.520 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 29.750 110.520 30.050 111.520 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 26.070 110.520 26.370 111.520 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 22.390 110.520 22.690 111.520 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 18.710 110.520 19.010 111.520 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 15.030 110.520 15.330 111.520 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 11.350 110.520 11.650 111.520 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 7.670 110.520 7.970 111.520 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.360500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met4 ;
        RECT 3.990 110.520 4.290 111.520 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 59.190 110.520 59.490 111.520 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met4 ;
        RECT 55.510 110.520 55.810 111.520 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 51.830 110.520 52.130 111.520 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 48.150 110.520 48.450 111.520 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 44.470 110.520 44.770 111.520 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 40.790 110.520 41.090 111.520 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 37.110 110.520 37.410 111.520 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 33.430 110.520 33.730 111.520 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met4 ;
        RECT 88.630 110.520 88.930 111.520 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 84.950 110.520 85.250 111.520 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 81.270 110.520 81.570 111.520 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met4 ;
        RECT 77.590 110.520 77.890 111.520 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met4 ;
        RECT 73.910 110.520 74.210 111.520 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.129500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met4 ;
        RECT 70.230 110.520 70.530 111.520 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.872000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met4 ;
        RECT 66.550 110.520 66.850 111.520 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.119500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met4 ;
        RECT 62.870 110.520 63.170 111.520 ;
    END
  END uo_out[7]
  OBS
      LAYER nwell ;
        RECT 2.570 107.385 158.430 108.990 ;
        RECT 2.570 101.945 158.430 104.775 ;
        RECT 2.570 96.505 158.430 99.335 ;
        RECT 2.570 91.065 158.430 93.895 ;
        RECT 2.570 85.625 158.430 88.455 ;
        RECT 2.570 80.185 158.430 83.015 ;
        RECT 2.570 74.745 158.430 77.575 ;
        RECT 2.570 69.305 158.430 72.135 ;
        RECT 2.570 63.865 158.430 66.695 ;
        RECT 2.570 58.425 158.430 61.255 ;
        RECT 2.570 52.985 158.430 55.815 ;
        RECT 2.570 47.545 158.430 50.375 ;
        RECT 2.570 42.105 158.430 44.935 ;
        RECT 2.570 36.665 158.430 39.495 ;
        RECT 2.570 31.225 158.430 34.055 ;
        RECT 2.570 25.785 158.430 28.615 ;
        RECT 2.570 20.345 158.430 23.175 ;
        RECT 2.570 14.905 158.430 17.735 ;
        RECT 2.570 9.465 158.430 12.295 ;
        RECT 2.570 4.025 158.430 6.855 ;
      LAYER li1 ;
        RECT 2.760 2.635 158.240 108.885 ;
      LAYER met1 ;
        RECT 2.760 2.480 159.040 109.440 ;
      LAYER met2 ;
        RECT 6.070 2.535 159.010 110.685 ;
      LAYER met3 ;
        RECT 3.950 2.555 159.030 110.665 ;
      LAYER met4 ;
        RECT 4.690 110.120 7.270 111.170 ;
        RECT 8.370 110.120 10.950 111.170 ;
        RECT 12.050 110.120 14.630 111.170 ;
        RECT 15.730 110.120 18.310 111.170 ;
        RECT 19.410 110.120 21.990 111.170 ;
        RECT 23.090 110.120 25.670 111.170 ;
        RECT 26.770 110.120 29.350 111.170 ;
        RECT 30.450 110.120 33.030 111.170 ;
        RECT 34.130 110.120 36.710 111.170 ;
        RECT 37.810 110.120 40.390 111.170 ;
        RECT 41.490 110.120 44.070 111.170 ;
        RECT 45.170 110.120 47.750 111.170 ;
        RECT 48.850 110.120 51.430 111.170 ;
        RECT 52.530 110.120 55.110 111.170 ;
        RECT 56.210 110.120 58.790 111.170 ;
        RECT 59.890 110.120 62.470 111.170 ;
        RECT 63.570 110.120 66.150 111.170 ;
        RECT 67.250 110.120 69.830 111.170 ;
        RECT 70.930 110.120 73.510 111.170 ;
        RECT 74.610 110.120 77.190 111.170 ;
        RECT 78.290 110.120 80.870 111.170 ;
        RECT 81.970 110.120 84.550 111.170 ;
        RECT 85.650 110.120 88.230 111.170 ;
        RECT 89.330 110.120 91.910 111.170 ;
        RECT 93.010 110.120 95.590 111.170 ;
        RECT 96.690 110.120 99.270 111.170 ;
        RECT 100.370 110.120 102.950 111.170 ;
        RECT 104.050 110.120 106.630 111.170 ;
        RECT 107.730 110.120 110.310 111.170 ;
        RECT 111.410 110.120 113.990 111.170 ;
        RECT 115.090 110.120 117.670 111.170 ;
        RECT 118.770 110.120 121.350 111.170 ;
        RECT 122.450 110.120 125.030 111.170 ;
        RECT 126.130 110.120 128.710 111.170 ;
        RECT 129.810 110.120 132.390 111.170 ;
        RECT 133.490 110.120 136.070 111.170 ;
        RECT 137.170 110.120 139.750 111.170 ;
        RECT 140.850 110.120 143.430 111.170 ;
        RECT 144.530 110.120 147.110 111.170 ;
        RECT 148.210 110.120 150.790 111.170 ;
        RECT 151.890 110.120 154.470 111.170 ;
        RECT 3.975 109.440 155.185 110.120 ;
        RECT 3.975 54.575 20.995 109.440 ;
        RECT 23.395 54.575 40.430 109.440 ;
        RECT 42.830 54.575 59.865 109.440 ;
        RECT 62.265 54.575 79.300 109.440 ;
        RECT 81.700 54.575 98.735 109.440 ;
        RECT 101.135 54.575 118.170 109.440 ;
        RECT 120.570 54.575 137.605 109.440 ;
        RECT 140.005 54.575 155.185 109.440 ;
  END
END tt_um_calculator_muehlbb
END LIBRARY

