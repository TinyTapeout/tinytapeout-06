VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_argunda_tiny_opamp
  CLASS BLOCK ;
  FOREIGN tt_um_argunda_tiny_opamp ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 154.870 224.760 155.170 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 158.550 224.760 158.850 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 151.190 224.760 151.490 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.350000 ;
    PORT
      LAYER met4 ;
        RECT 156.560 0.000 157.160 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.250000 ;
    PORT
      LAYER met4 ;
        RECT 134.480 0.000 135.080 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.250000 ;
    PORT
      LAYER met4 ;
        RECT 112.400 0.000 113.000 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 90.320 0.000 90.920 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 68.240 0.000 68.840 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 46.160 0.000 46.760 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 24.080 0.000 24.680 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 2.000 0.000 2.600 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 147.510 224.760 147.810 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 140.150 224.760 140.450 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 136.470 224.760 136.770 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 129.110 224.760 129.410 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 125.430 224.760 125.730 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.070 224.760 118.370 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 114.390 224.760 114.690 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.030 224.760 107.330 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 103.350 224.760 103.650 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 95.990 224.760 96.290 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 92.310 224.760 92.610 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 25.116999 ;
    PORT
      LAYER met4 ;
        RECT 29.750 224.760 30.050 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 25.116999 ;
    PORT
      LAYER met4 ;
        RECT 26.070 224.760 26.370 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 25.116999 ;
    PORT
      LAYER met4 ;
        RECT 22.390 224.760 22.690 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 25.116999 ;
    PORT
      LAYER met4 ;
        RECT 18.710 224.760 19.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 25.116999 ;
    PORT
      LAYER met4 ;
        RECT 15.030 224.760 15.330 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 25.116999 ;
    PORT
      LAYER met4 ;
        RECT 11.350 224.760 11.650 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 25.116999 ;
    PORT
      LAYER met4 ;
        RECT 7.670 224.760 7.970 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 25.116999 ;
    PORT
      LAYER met4 ;
        RECT 3.990 224.760 4.290 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 25.116999 ;
    PORT
      LAYER met4 ;
        RECT 59.190 224.760 59.490 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 25.116999 ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 25.116999 ;
    PORT
      LAYER met4 ;
        RECT 51.830 224.760 52.130 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 25.116999 ;
    PORT
      LAYER met4 ;
        RECT 48.150 224.760 48.450 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 25.116999 ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 25.116999 ;
    PORT
      LAYER met4 ;
        RECT 40.790 224.760 41.090 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 25.116999 ;
    PORT
      LAYER met4 ;
        RECT 37.110 224.760 37.410 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 25.116999 ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 25.116999 ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 25.116999 ;
    PORT
      LAYER met4 ;
        RECT 84.950 224.760 85.250 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 25.116999 ;
    PORT
      LAYER met4 ;
        RECT 81.270 224.760 81.570 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 25.116999 ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 25.116999 ;
    PORT
      LAYER met4 ;
        RECT 73.910 224.760 74.210 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 25.116999 ;
    PORT
      LAYER met4 ;
        RECT 70.230 224.760 70.530 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 25.116999 ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 25.116999 ;
    PORT
      LAYER met4 ;
        RECT 62.870 224.760 63.170 225.760 ;
    END
  END uo_out[7]
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 2.500 220.760 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 49.000 5.000 50.500 220.760 ;
    END
  END VGND
  OBS
      LAYER pwell ;
        RECT 144.740 87.580 153.360 89.590 ;
        RECT 141.570 75.160 144.670 85.990 ;
        RECT 143.140 74.190 143.370 74.220 ;
        RECT 143.180 73.860 143.370 74.190 ;
        RECT 144.710 73.860 144.940 74.220 ;
        RECT 142.490 63.030 145.590 73.860 ;
        RECT 141.560 58.940 146.160 61.400 ;
      LAYER nwell ;
        RECT 149.810 53.780 153.000 69.190 ;
      LAYER pwell ;
        RECT 141.740 42.520 146.340 44.980 ;
      LAYER nwell ;
        RECT 149.860 36.760 153.050 52.170 ;
      LAYER pwell ;
        RECT 142.510 18.030 145.610 35.730 ;
      LAYER nwell ;
        RECT 149.630 17.970 152.820 35.440 ;
      LAYER li1 ;
        RECT 144.920 89.240 153.180 89.410 ;
        RECT 144.920 89.070 145.090 89.240 ;
        RECT 144.770 88.170 145.260 89.070 ;
        RECT 153.010 88.970 153.180 89.240 ;
        RECT 145.570 88.410 147.730 88.760 ;
        RECT 150.370 88.410 152.530 88.760 ;
        RECT 152.990 88.220 153.280 88.970 ;
        RECT 144.920 87.930 145.090 88.170 ;
        RECT 153.010 87.930 153.180 88.220 ;
        RECT 144.920 87.760 153.180 87.930 ;
        RECT 141.750 85.640 144.490 85.810 ;
        RECT 141.750 75.510 141.920 85.640 ;
        RECT 142.600 85.070 143.640 85.240 ;
        RECT 142.260 83.010 142.430 85.010 ;
        RECT 143.810 83.010 143.980 85.010 ;
        RECT 142.600 82.780 143.640 82.950 ;
        RECT 142.260 80.720 142.430 82.720 ;
        RECT 143.810 80.720 143.980 82.720 ;
        RECT 142.600 80.490 143.640 80.660 ;
        RECT 142.260 78.430 142.430 80.430 ;
        RECT 143.810 78.430 143.980 80.430 ;
        RECT 142.600 78.200 143.640 78.370 ;
        RECT 142.260 76.140 142.430 78.140 ;
        RECT 143.810 76.140 143.980 78.140 ;
        RECT 142.600 75.910 143.640 76.080 ;
        RECT 144.320 75.510 144.490 85.640 ;
        RECT 141.750 75.340 144.490 75.510 ;
        RECT 142.670 73.510 145.410 73.680 ;
        RECT 142.670 63.380 142.840 73.510 ;
        RECT 143.520 72.940 144.560 73.110 ;
        RECT 143.180 70.880 143.350 72.880 ;
        RECT 144.730 70.880 144.900 72.880 ;
        RECT 143.520 70.650 144.560 70.820 ;
        RECT 143.180 68.590 143.350 70.590 ;
        RECT 144.730 68.590 144.900 70.590 ;
        RECT 143.520 68.360 144.560 68.530 ;
        RECT 143.180 66.300 143.350 68.300 ;
        RECT 144.730 66.300 144.900 68.300 ;
        RECT 143.520 66.070 144.560 66.240 ;
        RECT 143.180 64.010 143.350 66.010 ;
        RECT 144.730 64.010 144.900 66.010 ;
        RECT 143.520 63.780 144.560 63.950 ;
        RECT 145.240 63.380 145.410 73.510 ;
        RECT 142.670 63.210 145.410 63.380 ;
        RECT 149.990 68.840 152.820 69.010 ;
        RECT 141.740 61.050 145.980 61.220 ;
        RECT 141.740 59.290 141.910 61.050 ;
        RECT 142.590 60.480 145.130 60.650 ;
        RECT 142.250 59.920 142.420 60.420 ;
        RECT 145.300 59.920 145.470 60.420 ;
        RECT 142.590 59.690 145.130 59.860 ;
        RECT 145.810 59.290 145.980 61.050 ;
        RECT 141.740 59.120 145.980 59.290 ;
        RECT 149.990 54.130 150.160 68.840 ;
        RECT 150.885 68.270 151.925 68.440 ;
        RECT 150.500 66.210 150.670 68.210 ;
        RECT 152.140 66.210 152.310 68.210 ;
        RECT 150.885 65.980 151.925 66.150 ;
        RECT 150.500 63.920 150.670 65.920 ;
        RECT 152.140 63.920 152.310 65.920 ;
        RECT 150.885 63.690 151.925 63.860 ;
        RECT 150.500 61.630 150.670 63.630 ;
        RECT 152.140 61.630 152.310 63.630 ;
        RECT 150.885 61.400 151.925 61.570 ;
        RECT 150.500 59.340 150.670 61.340 ;
        RECT 152.140 59.340 152.310 61.340 ;
        RECT 150.885 59.110 151.925 59.280 ;
        RECT 150.500 57.050 150.670 59.050 ;
        RECT 152.140 57.050 152.310 59.050 ;
        RECT 150.885 56.820 151.925 56.990 ;
        RECT 150.500 54.760 150.670 56.760 ;
        RECT 152.140 54.760 152.310 56.760 ;
        RECT 150.885 54.530 151.925 54.700 ;
        RECT 152.650 54.130 152.820 68.840 ;
        RECT 149.990 53.960 152.820 54.130 ;
        RECT 150.040 51.820 152.870 51.990 ;
        RECT 141.920 44.630 146.160 44.800 ;
        RECT 141.920 44.310 142.090 44.630 ;
        RECT 141.730 43.190 142.090 44.310 ;
        RECT 142.770 44.060 145.310 44.230 ;
        RECT 142.430 43.500 142.600 44.000 ;
        RECT 145.480 43.500 145.650 44.000 ;
        RECT 142.770 43.270 145.310 43.440 ;
        RECT 141.920 42.870 142.090 43.190 ;
        RECT 145.990 42.870 146.160 44.630 ;
        RECT 141.920 42.700 146.160 42.870 ;
        RECT 150.040 37.110 150.210 51.820 ;
        RECT 150.935 51.250 151.975 51.420 ;
        RECT 150.550 49.190 150.720 51.190 ;
        RECT 152.190 49.190 152.360 51.190 ;
        RECT 150.935 48.960 151.975 49.130 ;
        RECT 150.550 46.900 150.720 48.900 ;
        RECT 152.190 46.900 152.360 48.900 ;
        RECT 150.935 46.670 151.975 46.840 ;
        RECT 150.550 44.610 150.720 46.610 ;
        RECT 152.190 44.610 152.360 46.610 ;
        RECT 150.935 44.380 151.975 44.550 ;
        RECT 150.550 42.320 150.720 44.320 ;
        RECT 152.190 42.320 152.360 44.320 ;
        RECT 150.935 42.090 151.975 42.260 ;
        RECT 150.550 40.030 150.720 42.030 ;
        RECT 152.190 40.030 152.360 42.030 ;
        RECT 150.935 39.800 151.975 39.970 ;
        RECT 150.550 37.740 150.720 39.740 ;
        RECT 152.190 37.740 152.360 39.740 ;
        RECT 150.935 37.510 151.975 37.680 ;
        RECT 152.700 37.110 152.870 51.820 ;
        RECT 150.040 36.940 152.870 37.110 ;
        RECT 142.690 35.380 145.430 35.550 ;
        RECT 142.690 18.380 142.860 35.380 ;
        RECT 143.540 34.810 144.580 34.980 ;
        RECT 143.200 32.750 143.370 34.750 ;
        RECT 144.750 32.750 144.920 34.750 ;
        RECT 143.540 32.520 144.580 32.690 ;
        RECT 143.200 30.460 143.370 32.460 ;
        RECT 144.750 30.460 144.920 32.460 ;
        RECT 143.540 30.230 144.580 30.400 ;
        RECT 143.200 28.170 143.370 30.170 ;
        RECT 144.750 28.170 144.920 30.170 ;
        RECT 143.540 27.940 144.580 28.110 ;
        RECT 143.200 25.880 143.370 27.880 ;
        RECT 144.750 25.880 144.920 27.880 ;
        RECT 143.540 25.650 144.580 25.820 ;
        RECT 143.200 23.590 143.370 25.590 ;
        RECT 144.750 23.590 144.920 25.590 ;
        RECT 143.540 23.360 144.580 23.530 ;
        RECT 143.200 21.300 143.370 23.300 ;
        RECT 144.750 21.300 144.920 23.300 ;
        RECT 143.540 21.070 144.580 21.240 ;
        RECT 143.200 19.010 143.370 21.010 ;
        RECT 144.750 19.010 144.920 21.010 ;
        RECT 143.540 18.780 144.580 18.950 ;
        RECT 145.260 18.380 145.430 35.380 ;
        RECT 142.690 18.210 145.430 18.380 ;
        RECT 149.810 35.090 152.640 35.260 ;
        RECT 149.810 18.320 149.980 35.090 ;
        RECT 150.705 34.520 151.745 34.690 ;
        RECT 150.320 33.960 150.490 34.460 ;
        RECT 151.960 33.960 152.130 34.460 ;
        RECT 150.705 33.730 151.745 33.900 ;
        RECT 150.320 33.170 150.490 33.670 ;
        RECT 151.960 33.170 152.130 33.670 ;
        RECT 150.705 32.940 151.745 33.110 ;
        RECT 150.320 32.380 150.490 32.880 ;
        RECT 151.960 32.380 152.130 32.880 ;
        RECT 150.705 32.150 151.745 32.320 ;
        RECT 150.320 31.590 150.490 32.090 ;
        RECT 151.960 31.590 152.130 32.090 ;
        RECT 150.705 31.360 151.745 31.530 ;
        RECT 150.320 30.800 150.490 31.300 ;
        RECT 151.960 30.800 152.130 31.300 ;
        RECT 150.705 30.570 151.745 30.740 ;
        RECT 150.320 30.010 150.490 30.510 ;
        RECT 151.960 30.010 152.130 30.510 ;
        RECT 150.705 29.780 151.745 29.950 ;
        RECT 150.320 29.220 150.490 29.720 ;
        RECT 151.960 29.220 152.130 29.720 ;
        RECT 150.705 28.990 151.745 29.160 ;
        RECT 150.320 28.430 150.490 28.930 ;
        RECT 151.960 28.430 152.130 28.930 ;
        RECT 150.705 28.200 151.745 28.370 ;
        RECT 150.320 27.640 150.490 28.140 ;
        RECT 151.960 27.640 152.130 28.140 ;
        RECT 150.705 27.410 151.745 27.580 ;
        RECT 150.320 26.850 150.490 27.350 ;
        RECT 151.960 26.850 152.130 27.350 ;
        RECT 150.705 26.620 151.745 26.790 ;
        RECT 150.320 26.060 150.490 26.560 ;
        RECT 151.960 26.060 152.130 26.560 ;
        RECT 150.705 25.830 151.745 26.000 ;
        RECT 150.320 25.270 150.490 25.770 ;
        RECT 151.960 25.270 152.130 25.770 ;
        RECT 150.705 25.040 151.745 25.210 ;
        RECT 150.320 24.480 150.490 24.980 ;
        RECT 151.960 24.480 152.130 24.980 ;
        RECT 150.705 24.250 151.745 24.420 ;
        RECT 150.320 23.690 150.490 24.190 ;
        RECT 151.960 23.690 152.130 24.190 ;
        RECT 150.705 23.460 151.745 23.630 ;
        RECT 150.320 22.900 150.490 23.400 ;
        RECT 151.960 22.900 152.130 23.400 ;
        RECT 150.705 22.670 151.745 22.840 ;
        RECT 150.320 22.110 150.490 22.610 ;
        RECT 151.960 22.110 152.130 22.610 ;
        RECT 150.705 21.880 151.745 22.050 ;
        RECT 150.320 21.320 150.490 21.820 ;
        RECT 151.960 21.320 152.130 21.820 ;
        RECT 150.705 21.090 151.745 21.260 ;
        RECT 150.320 20.530 150.490 21.030 ;
        RECT 151.960 20.530 152.130 21.030 ;
        RECT 150.705 20.300 151.745 20.470 ;
        RECT 150.320 19.740 150.490 20.240 ;
        RECT 151.960 19.740 152.130 20.240 ;
        RECT 150.705 19.510 151.745 19.680 ;
        RECT 150.320 18.950 150.490 19.450 ;
        RECT 151.960 18.950 152.130 19.450 ;
        RECT 150.705 18.720 151.745 18.890 ;
        RECT 152.470 18.320 152.640 35.090 ;
        RECT 149.810 18.150 152.640 18.320 ;
      LAYER mcon ;
        RECT 145.660 88.490 147.645 88.680 ;
        RECT 150.455 88.490 152.440 88.680 ;
        RECT 141.750 75.820 141.920 85.330 ;
        RECT 142.680 85.070 143.560 85.240 ;
        RECT 142.260 83.090 142.430 84.930 ;
        RECT 143.810 83.090 143.980 84.930 ;
        RECT 142.680 82.780 143.560 82.950 ;
        RECT 142.260 80.800 142.430 82.640 ;
        RECT 143.810 80.800 143.980 82.640 ;
        RECT 142.680 80.490 143.560 80.660 ;
        RECT 142.260 78.510 142.430 80.350 ;
        RECT 143.810 78.510 143.980 80.350 ;
        RECT 142.680 78.200 143.560 78.370 ;
        RECT 142.260 76.220 142.430 78.060 ;
        RECT 143.810 76.220 143.980 78.060 ;
        RECT 142.680 75.910 143.560 76.080 ;
        RECT 142.670 63.690 142.840 73.200 ;
        RECT 143.600 72.940 144.480 73.110 ;
        RECT 143.180 70.960 143.350 72.800 ;
        RECT 144.730 70.960 144.900 72.800 ;
        RECT 143.600 70.650 144.480 70.820 ;
        RECT 143.180 68.670 143.350 70.510 ;
        RECT 144.730 68.670 144.900 70.510 ;
        RECT 143.600 68.360 144.480 68.530 ;
        RECT 143.180 66.380 143.350 68.220 ;
        RECT 144.730 66.380 144.900 68.220 ;
        RECT 143.600 66.070 144.480 66.240 ;
        RECT 143.180 64.090 143.350 65.930 ;
        RECT 144.730 64.090 144.900 65.930 ;
        RECT 143.600 63.780 144.480 63.950 ;
        RECT 141.740 59.600 141.910 60.740 ;
        RECT 142.670 60.480 145.050 60.650 ;
        RECT 142.250 60.000 142.420 60.340 ;
        RECT 145.300 60.000 145.470 60.340 ;
        RECT 142.670 59.690 145.050 59.860 ;
        RECT 150.965 68.270 151.845 68.440 ;
        RECT 150.500 66.290 150.670 68.130 ;
        RECT 152.140 66.290 152.310 68.130 ;
        RECT 150.965 65.980 151.845 66.150 ;
        RECT 150.500 64.000 150.670 65.840 ;
        RECT 152.140 64.000 152.310 65.840 ;
        RECT 150.965 63.690 151.845 63.860 ;
        RECT 150.500 61.710 150.670 63.550 ;
        RECT 152.140 61.710 152.310 63.550 ;
        RECT 150.965 61.400 151.845 61.570 ;
        RECT 150.500 59.420 150.670 61.260 ;
        RECT 152.140 59.420 152.310 61.260 ;
        RECT 150.965 59.110 151.845 59.280 ;
        RECT 150.500 57.130 150.670 58.970 ;
        RECT 152.140 57.130 152.310 58.970 ;
        RECT 150.965 56.820 151.845 56.990 ;
        RECT 150.500 54.840 150.670 56.680 ;
        RECT 152.140 54.840 152.310 56.680 ;
        RECT 150.965 54.530 151.845 54.700 ;
        RECT 152.650 54.440 152.820 68.530 ;
        RECT 141.730 43.190 142.080 44.310 ;
        RECT 142.850 44.060 145.230 44.230 ;
        RECT 142.430 43.580 142.600 43.920 ;
        RECT 145.480 43.580 145.650 43.920 ;
        RECT 142.850 43.270 145.230 43.440 ;
        RECT 151.015 51.250 151.895 51.420 ;
        RECT 150.550 49.270 150.720 51.110 ;
        RECT 152.190 49.270 152.360 51.110 ;
        RECT 151.015 48.960 151.895 49.130 ;
        RECT 150.550 46.980 150.720 48.820 ;
        RECT 152.190 46.980 152.360 48.820 ;
        RECT 151.015 46.670 151.895 46.840 ;
        RECT 150.550 44.690 150.720 46.530 ;
        RECT 152.190 44.690 152.360 46.530 ;
        RECT 151.015 44.380 151.895 44.550 ;
        RECT 150.550 42.400 150.720 44.240 ;
        RECT 152.190 42.400 152.360 44.240 ;
        RECT 151.015 42.090 151.895 42.260 ;
        RECT 150.550 40.110 150.720 41.950 ;
        RECT 152.190 40.110 152.360 41.950 ;
        RECT 151.015 39.800 151.895 39.970 ;
        RECT 150.550 37.820 150.720 39.660 ;
        RECT 152.190 37.820 152.360 39.660 ;
        RECT 151.015 37.510 151.895 37.680 ;
        RECT 152.700 37.420 152.870 51.510 ;
        RECT 142.690 18.690 142.860 35.070 ;
        RECT 143.620 34.810 144.500 34.980 ;
        RECT 143.200 32.830 143.370 34.670 ;
        RECT 144.750 32.830 144.920 34.670 ;
        RECT 143.620 32.520 144.500 32.690 ;
        RECT 143.200 30.540 143.370 32.380 ;
        RECT 144.750 30.540 144.920 32.380 ;
        RECT 143.620 30.230 144.500 30.400 ;
        RECT 143.200 28.250 143.370 30.090 ;
        RECT 144.750 28.250 144.920 30.090 ;
        RECT 143.620 27.940 144.500 28.110 ;
        RECT 143.200 25.960 143.370 27.800 ;
        RECT 144.750 25.960 144.920 27.800 ;
        RECT 143.620 25.650 144.500 25.820 ;
        RECT 143.200 23.670 143.370 25.510 ;
        RECT 144.750 23.670 144.920 25.510 ;
        RECT 143.620 23.360 144.500 23.530 ;
        RECT 143.200 21.380 143.370 23.220 ;
        RECT 144.750 21.380 144.920 23.220 ;
        RECT 143.620 21.070 144.500 21.240 ;
        RECT 143.200 19.090 143.370 20.930 ;
        RECT 144.750 19.090 144.920 20.930 ;
        RECT 143.620 18.780 144.500 18.950 ;
        RECT 150.785 34.520 151.665 34.690 ;
        RECT 150.320 34.040 150.490 34.380 ;
        RECT 151.960 34.040 152.130 34.380 ;
        RECT 150.785 33.730 151.665 33.900 ;
        RECT 150.320 33.250 150.490 33.590 ;
        RECT 151.960 33.250 152.130 33.590 ;
        RECT 150.785 32.940 151.665 33.110 ;
        RECT 150.320 32.460 150.490 32.800 ;
        RECT 151.960 32.460 152.130 32.800 ;
        RECT 150.785 32.150 151.665 32.320 ;
        RECT 150.320 31.670 150.490 32.010 ;
        RECT 151.960 31.670 152.130 32.010 ;
        RECT 150.785 31.360 151.665 31.530 ;
        RECT 150.320 30.880 150.490 31.220 ;
        RECT 151.960 30.880 152.130 31.220 ;
        RECT 150.785 30.570 151.665 30.740 ;
        RECT 150.320 30.090 150.490 30.430 ;
        RECT 151.960 30.090 152.130 30.430 ;
        RECT 150.785 29.780 151.665 29.950 ;
        RECT 150.320 29.300 150.490 29.640 ;
        RECT 151.960 29.300 152.130 29.640 ;
        RECT 150.785 28.990 151.665 29.160 ;
        RECT 150.320 28.510 150.490 28.850 ;
        RECT 151.960 28.510 152.130 28.850 ;
        RECT 150.785 28.200 151.665 28.370 ;
        RECT 150.320 27.720 150.490 28.060 ;
        RECT 151.960 27.720 152.130 28.060 ;
        RECT 150.785 27.410 151.665 27.580 ;
        RECT 150.320 26.930 150.490 27.270 ;
        RECT 151.960 26.930 152.130 27.270 ;
        RECT 150.785 26.620 151.665 26.790 ;
        RECT 150.320 26.140 150.490 26.480 ;
        RECT 151.960 26.140 152.130 26.480 ;
        RECT 150.785 25.830 151.665 26.000 ;
        RECT 150.320 25.350 150.490 25.690 ;
        RECT 151.960 25.350 152.130 25.690 ;
        RECT 150.785 25.040 151.665 25.210 ;
        RECT 150.320 24.560 150.490 24.900 ;
        RECT 151.960 24.560 152.130 24.900 ;
        RECT 150.785 24.250 151.665 24.420 ;
        RECT 150.320 23.770 150.490 24.110 ;
        RECT 151.960 23.770 152.130 24.110 ;
        RECT 150.785 23.460 151.665 23.630 ;
        RECT 150.320 22.980 150.490 23.320 ;
        RECT 151.960 22.980 152.130 23.320 ;
        RECT 150.785 22.670 151.665 22.840 ;
        RECT 150.320 22.190 150.490 22.530 ;
        RECT 151.960 22.190 152.130 22.530 ;
        RECT 150.785 21.880 151.665 22.050 ;
        RECT 150.320 21.400 150.490 21.740 ;
        RECT 151.960 21.400 152.130 21.740 ;
        RECT 150.785 21.090 151.665 21.260 ;
        RECT 150.320 20.610 150.490 20.950 ;
        RECT 151.960 20.610 152.130 20.950 ;
        RECT 150.785 20.300 151.665 20.470 ;
        RECT 150.320 19.820 150.490 20.160 ;
        RECT 151.960 19.820 152.130 20.160 ;
        RECT 150.785 19.510 151.665 19.680 ;
        RECT 150.320 19.030 150.490 19.370 ;
        RECT 151.960 19.030 152.130 19.370 ;
        RECT 150.785 18.720 151.665 18.890 ;
        RECT 150.290 18.150 152.160 18.320 ;
      LAYER met1 ;
        RECT 140.180 132.070 140.540 132.370 ;
        RECT 140.210 91.000 140.510 132.070 ;
        RECT 156.780 107.820 158.340 109.320 ;
        RECT 156.810 91.030 158.310 107.820 ;
        RECT 137.690 90.020 154.010 91.000 ;
        RECT 137.700 89.670 141.190 90.020 ;
        RECT 137.700 87.550 145.340 89.670 ;
        RECT 145.640 88.710 147.740 89.700 ;
        RECT 145.600 88.460 147.740 88.710 ;
        RECT 137.700 85.810 141.190 87.550 ;
        RECT 145.640 87.030 147.740 88.460 ;
        RECT 149.650 87.460 152.800 89.620 ;
        RECT 141.970 86.400 147.740 87.030 ;
        RECT 137.700 75.070 141.950 85.810 ;
        RECT 142.260 84.990 142.450 86.400 ;
        RECT 142.590 85.990 147.740 86.400 ;
        RECT 142.230 83.030 142.460 84.990 ;
        RECT 142.600 84.980 143.640 85.990 ;
        RECT 143.780 84.930 144.010 84.990 ;
        RECT 145.640 84.930 147.740 85.990 ;
        RECT 142.260 82.700 142.450 83.030 ;
        RECT 142.640 82.980 143.620 83.370 ;
        RECT 143.780 83.090 147.740 84.930 ;
        RECT 150.640 86.910 152.800 87.460 ;
        RECT 152.950 87.380 153.980 90.020 ;
        RECT 154.770 87.810 158.310 91.030 ;
        RECT 154.770 86.910 158.270 87.810 ;
        RECT 150.640 84.750 158.270 86.910 ;
        RECT 143.780 83.030 144.010 83.090 ;
        RECT 142.620 82.750 143.620 82.980 ;
        RECT 142.230 80.740 142.460 82.700 ;
        RECT 142.640 82.420 143.620 82.750 ;
        RECT 143.780 82.640 144.010 82.700 ;
        RECT 145.640 82.640 147.740 83.090 ;
        RECT 143.780 82.220 147.740 82.640 ;
        RECT 142.630 81.310 147.740 82.220 ;
        RECT 142.260 80.410 142.450 80.740 ;
        RECT 142.640 80.690 143.610 81.310 ;
        RECT 143.780 80.790 147.740 81.310 ;
        RECT 143.780 80.740 144.010 80.790 ;
        RECT 144.810 80.760 147.740 80.790 ;
        RECT 142.620 80.460 143.620 80.690 ;
        RECT 142.230 78.450 142.460 80.410 ;
        RECT 142.640 79.880 143.610 80.460 ;
        RECT 143.780 80.350 144.010 80.410 ;
        RECT 145.640 80.350 147.740 80.760 ;
        RECT 143.780 79.880 147.740 80.350 ;
        RECT 142.620 78.970 147.740 79.880 ;
        RECT 142.640 78.920 143.610 78.970 ;
        RECT 142.260 78.120 142.450 78.450 ;
        RECT 142.640 78.400 143.620 78.740 ;
        RECT 143.780 78.510 147.740 78.970 ;
        RECT 143.780 78.450 144.010 78.510 ;
        RECT 142.620 78.170 143.620 78.400 ;
        RECT 142.230 76.160 142.460 78.120 ;
        RECT 142.640 77.790 143.620 78.170 ;
        RECT 143.780 78.060 144.010 78.120 ;
        RECT 145.640 78.060 147.740 78.510 ;
        RECT 143.780 77.220 147.740 78.060 ;
        RECT 142.640 76.220 147.740 77.220 ;
        RECT 142.640 76.210 144.180 76.220 ;
        RECT 145.640 76.210 147.740 76.220 ;
        RECT 142.640 76.160 144.010 76.210 ;
        RECT 142.260 76.050 142.450 76.160 ;
        RECT 142.640 76.110 143.780 76.160 ;
        RECT 142.620 76.040 143.780 76.110 ;
        RECT 145.640 76.080 147.750 76.210 ;
        RECT 142.620 75.880 143.620 76.040 ;
        RECT 142.640 75.870 143.570 75.880 ;
        RECT 137.700 75.050 141.940 75.070 ;
        RECT 137.700 73.890 141.190 75.050 ;
        RECT 145.640 74.430 148.995 76.080 ;
        RECT 143.140 74.190 148.995 74.430 ;
        RECT 143.180 73.960 148.995 74.190 ;
        RECT 137.700 63.080 142.870 73.890 ;
        RECT 143.180 72.860 143.370 73.960 ;
        RECT 143.580 73.140 144.500 73.490 ;
        RECT 143.540 72.910 144.540 73.140 ;
        RECT 143.150 70.900 143.380 72.860 ;
        RECT 143.580 72.460 144.500 72.910 ;
        RECT 144.710 72.860 144.940 73.960 ;
        RECT 143.180 70.570 143.370 70.900 ;
        RECT 143.560 70.850 144.550 71.440 ;
        RECT 144.700 70.900 144.940 72.860 ;
        RECT 143.540 70.620 144.550 70.850 ;
        RECT 143.150 68.610 143.380 70.570 ;
        RECT 143.560 70.050 144.550 70.620 ;
        RECT 144.710 70.570 144.940 70.900 ;
        RECT 143.180 68.280 143.370 68.610 ;
        RECT 143.600 68.560 144.520 68.930 ;
        RECT 144.700 68.610 144.940 70.570 ;
        RECT 143.540 68.330 144.540 68.560 ;
        RECT 143.150 66.320 143.380 68.280 ;
        RECT 143.600 67.900 144.520 68.330 ;
        RECT 144.710 68.280 144.940 68.610 ;
        RECT 143.180 65.990 143.370 66.320 ;
        RECT 143.540 66.270 144.530 66.860 ;
        RECT 144.700 66.320 144.940 68.280 ;
        RECT 143.540 66.040 144.540 66.270 ;
        RECT 143.150 64.030 143.380 65.990 ;
        RECT 143.540 65.470 144.530 66.040 ;
        RECT 144.710 65.990 144.940 66.320 ;
        RECT 143.570 63.980 144.490 64.360 ;
        RECT 144.700 64.050 144.940 65.990 ;
        RECT 144.700 64.030 144.930 64.050 ;
        RECT 143.540 63.750 144.540 63.980 ;
        RECT 143.570 63.330 144.490 63.750 ;
        RECT 137.700 63.050 142.860 63.080 ;
        RECT 137.700 61.290 141.190 63.050 ;
        RECT 143.590 62.740 144.480 63.330 ;
        RECT 143.590 62.030 146.450 62.740 ;
        RECT 137.700 59.050 141.980 61.290 ;
        RECT 143.590 60.680 144.480 62.030 ;
        RECT 142.610 60.450 145.110 60.680 ;
        RECT 142.250 60.400 142.420 60.430 ;
        RECT 145.300 60.400 145.470 60.420 ;
        RECT 142.220 59.940 142.450 60.400 ;
        RECT 145.270 59.940 145.500 60.400 ;
        RECT 137.700 44.930 141.190 59.050 ;
        RECT 142.250 56.970 142.420 59.940 ;
        RECT 142.610 59.660 145.110 59.890 ;
        RECT 142.670 57.780 145.060 59.660 ;
        RECT 142.140 56.780 143.140 56.970 ;
        RECT 145.300 56.780 145.470 59.940 ;
        RECT 142.140 56.610 145.470 56.780 ;
        RECT 142.140 55.970 143.140 56.610 ;
        RECT 142.360 53.950 142.960 55.970 ;
        RECT 142.330 53.350 142.990 53.950 ;
        RECT 143.765 51.125 144.475 51.155 ;
        RECT 145.740 51.125 146.450 62.030 ;
        RECT 146.885 61.350 148.995 73.960 ;
        RECT 150.500 72.000 152.400 72.010 ;
        RECT 150.460 69.420 152.400 72.000 ;
        RECT 142.380 50.300 143.040 50.900 ;
        RECT 143.765 50.415 146.450 51.125 ;
        RECT 146.650 59.245 148.995 61.350 ;
        RECT 150.470 68.570 150.730 69.420 ;
        RECT 152.130 69.270 152.400 69.420 ;
        RECT 152.130 68.570 152.310 69.270 ;
        RECT 150.470 68.380 152.310 68.570 ;
        RECT 150.470 63.860 150.730 68.380 ;
        RECT 150.905 68.240 151.905 68.380 ;
        RECT 152.130 68.190 152.310 68.380 ;
        RECT 152.620 68.530 152.880 68.630 ;
        RECT 154.780 68.530 158.270 84.750 ;
        RECT 150.930 66.180 151.920 66.420 ;
        RECT 152.110 66.230 152.340 68.190 ;
        RECT 150.905 65.950 151.920 66.180 ;
        RECT 150.930 65.750 151.920 65.950 ;
        RECT 152.130 65.900 152.310 66.230 ;
        RECT 152.110 63.940 152.340 65.900 ;
        RECT 150.905 63.860 151.905 63.890 ;
        RECT 150.470 63.690 151.970 63.860 ;
        RECT 150.470 60.060 150.730 63.690 ;
        RECT 150.905 63.660 151.905 63.690 ;
        RECT 152.130 63.610 152.310 63.940 ;
        RECT 150.900 61.600 151.890 61.830 ;
        RECT 152.110 61.650 152.340 63.610 ;
        RECT 150.900 61.370 151.905 61.600 ;
        RECT 150.900 61.160 151.890 61.370 ;
        RECT 152.130 61.320 152.310 61.650 ;
        RECT 149.900 59.280 150.730 60.060 ;
        RECT 152.110 59.360 152.340 61.320 ;
        RECT 150.905 59.280 151.905 59.310 ;
        RECT 143.765 50.385 144.475 50.415 ;
        RECT 142.410 49.260 143.010 50.300 ;
        RECT 142.160 48.285 143.160 49.260 ;
        RECT 142.160 48.260 145.665 48.285 ;
        RECT 142.430 48.095 145.665 48.260 ;
        RECT 137.700 44.340 142.090 44.930 ;
        RECT 137.700 43.160 142.120 44.340 ;
        RECT 142.430 43.980 142.620 48.095 ;
        RECT 143.765 47.535 144.460 47.585 ;
        RECT 143.765 44.260 144.610 47.535 ;
        RECT 142.790 44.030 145.290 44.260 ;
        RECT 143.765 44.000 144.610 44.030 ;
        RECT 145.475 43.980 145.665 48.095 ;
        RECT 142.400 43.520 142.630 43.980 ;
        RECT 145.450 43.520 145.680 43.980 ;
        RECT 142.430 43.500 142.620 43.520 ;
        RECT 145.475 43.475 145.665 43.520 ;
        RECT 142.790 43.240 145.290 43.470 ;
        RECT 137.700 42.680 142.090 43.160 ;
        RECT 137.700 35.080 141.190 42.680 ;
        RECT 142.820 40.610 145.280 43.240 ;
        RECT 146.650 38.080 148.400 59.245 ;
        RECT 149.900 59.110 151.905 59.280 ;
        RECT 148.810 58.750 149.510 58.800 ;
        RECT 149.900 58.750 150.730 59.110 ;
        RECT 150.905 59.080 151.905 59.110 ;
        RECT 152.130 59.030 152.310 59.360 ;
        RECT 148.810 58.030 150.730 58.750 ;
        RECT 148.810 58.000 149.510 58.030 ;
        RECT 149.900 55.130 150.730 58.030 ;
        RECT 150.900 57.020 151.890 57.250 ;
        RECT 152.110 57.070 152.340 59.030 ;
        RECT 150.900 56.790 151.905 57.020 ;
        RECT 150.900 56.580 151.890 56.790 ;
        RECT 152.130 56.740 152.310 57.070 ;
        RECT 143.120 36.295 148.400 38.080 ;
        RECT 150.470 54.710 150.730 55.130 ;
        RECT 152.110 54.780 152.340 56.740 ;
        RECT 150.905 54.710 151.905 54.730 ;
        RECT 150.470 54.540 151.905 54.710 ;
        RECT 150.470 53.520 150.730 54.540 ;
        RECT 150.905 54.500 151.905 54.540 ;
        RECT 152.140 53.520 152.310 54.780 ;
        RECT 152.620 54.440 158.270 68.530 ;
        RECT 152.620 54.360 152.880 54.440 ;
        RECT 150.470 52.340 152.310 53.520 ;
        RECT 150.470 51.170 150.730 52.340 ;
        RECT 150.470 49.210 150.750 51.170 ;
        RECT 150.950 50.900 151.960 51.750 ;
        RECT 152.140 51.190 152.310 52.340 ;
        RECT 152.670 51.500 152.980 51.570 ;
        RECT 154.780 51.500 158.270 54.440 ;
        RECT 150.470 48.880 150.730 49.210 ;
        RECT 150.940 49.160 151.950 49.460 ;
        RECT 152.140 49.190 152.390 51.190 ;
        RECT 150.940 48.930 151.955 49.160 ;
        RECT 150.470 46.920 150.750 48.880 ;
        RECT 150.940 48.610 151.950 48.930 ;
        RECT 152.140 48.880 152.310 49.190 ;
        RECT 150.470 46.590 150.730 46.920 ;
        RECT 150.470 44.630 150.750 46.590 ;
        RECT 150.950 46.360 151.960 47.210 ;
        RECT 150.470 44.300 150.730 44.630 ;
        RECT 150.960 44.580 151.970 44.900 ;
        RECT 150.955 44.350 151.970 44.580 ;
        RECT 150.470 42.340 150.750 44.300 ;
        RECT 150.960 44.050 151.970 44.350 ;
        RECT 152.140 44.630 152.390 48.880 ;
        RECT 152.140 44.310 152.310 44.630 ;
        RECT 150.470 42.010 150.730 42.340 ;
        RECT 150.940 42.290 151.950 42.620 ;
        RECT 152.140 42.340 152.390 44.310 ;
        RECT 150.940 42.060 151.955 42.290 ;
        RECT 150.470 40.050 150.750 42.010 ;
        RECT 150.940 41.770 151.950 42.060 ;
        RECT 152.140 42.030 152.310 42.340 ;
        RECT 150.470 39.720 150.730 40.050 ;
        RECT 150.940 40.000 151.950 40.330 ;
        RECT 152.140 40.050 152.390 42.030 ;
        RECT 150.940 39.770 151.955 40.000 ;
        RECT 150.470 37.760 150.750 39.720 ;
        RECT 150.940 39.480 151.950 39.770 ;
        RECT 152.140 39.740 152.310 40.050 ;
        RECT 150.970 37.950 151.980 38.010 ;
        RECT 150.470 37.750 150.730 37.760 ;
        RECT 143.120 36.290 146.810 36.295 ;
        RECT 142.630 35.080 142.920 35.130 ;
        RECT 137.700 34.990 142.920 35.080 ;
        RECT 137.700 18.750 142.890 34.990 ;
        RECT 143.190 34.730 143.400 36.290 ;
        RECT 143.580 35.010 144.580 35.160 ;
        RECT 143.560 34.780 144.580 35.010 ;
        RECT 143.170 32.770 143.400 34.730 ;
        RECT 143.580 34.650 144.580 34.780 ;
        RECT 144.720 34.730 144.930 36.290 ;
        RECT 150.950 36.270 151.990 37.950 ;
        RECT 152.140 37.760 152.390 39.740 ;
        RECT 152.140 37.745 152.310 37.760 ;
        RECT 152.670 37.740 158.270 51.500 ;
        RECT 152.640 37.410 158.270 37.740 ;
        RECT 152.640 37.300 152.960 37.410 ;
        RECT 150.290 35.260 152.160 36.270 ;
        RECT 150.290 35.040 152.130 35.260 ;
        RECT 143.190 32.440 143.400 32.770 ;
        RECT 143.570 32.720 144.570 32.880 ;
        RECT 143.560 32.490 144.570 32.720 ;
        RECT 143.170 30.480 143.400 32.440 ;
        RECT 143.570 32.370 144.570 32.490 ;
        RECT 144.720 32.770 144.950 34.730 ;
        RECT 144.720 32.440 144.930 32.770 ;
        RECT 143.190 30.150 143.400 30.480 ;
        RECT 143.580 30.430 144.580 30.580 ;
        RECT 143.560 30.200 144.580 30.430 ;
        RECT 143.170 28.190 143.400 30.150 ;
        RECT 143.580 30.070 144.580 30.200 ;
        RECT 144.720 30.480 144.950 32.440 ;
        RECT 144.720 30.150 144.930 30.480 ;
        RECT 143.190 27.860 143.400 28.190 ;
        RECT 143.170 25.900 143.400 27.860 ;
        RECT 143.550 28.140 144.550 28.250 ;
        RECT 144.720 28.190 144.950 30.150 ;
        RECT 143.550 27.910 144.560 28.140 ;
        RECT 143.550 27.740 144.550 27.910 ;
        RECT 144.720 27.860 144.930 28.190 ;
        RECT 143.190 25.570 143.400 25.900 ;
        RECT 143.580 25.850 144.580 26.000 ;
        RECT 143.560 25.620 144.580 25.850 ;
        RECT 143.170 23.610 143.400 25.570 ;
        RECT 143.580 25.490 144.580 25.620 ;
        RECT 144.720 25.900 144.950 27.860 ;
        RECT 144.720 25.570 144.930 25.900 ;
        RECT 143.190 23.280 143.400 23.610 ;
        RECT 143.570 23.560 144.570 23.710 ;
        RECT 143.560 23.330 144.570 23.560 ;
        RECT 143.170 21.320 143.400 23.280 ;
        RECT 143.570 23.200 144.570 23.330 ;
        RECT 144.720 23.610 144.950 25.570 ;
        RECT 144.720 23.280 144.930 23.610 ;
        RECT 143.190 20.990 143.400 21.320 ;
        RECT 143.570 21.270 144.570 21.410 ;
        RECT 143.560 21.040 144.570 21.270 ;
        RECT 143.170 19.030 143.400 20.990 ;
        RECT 143.570 20.900 144.570 21.040 ;
        RECT 144.720 21.320 144.950 23.280 ;
        RECT 144.720 20.990 144.930 21.320 ;
        RECT 143.190 19.000 143.400 19.030 ;
        RECT 143.550 18.980 144.550 19.120 ;
        RECT 144.720 19.030 144.950 20.990 ;
        RECT 145.690 19.300 146.860 32.850 ;
        RECT 147.370 20.090 149.060 32.880 ;
        RECT 147.070 19.390 149.060 20.090 ;
        RECT 147.070 19.300 148.320 19.390 ;
        RECT 143.550 18.750 144.560 18.980 ;
        RECT 144.720 18.970 144.930 19.030 ;
        RECT 145.690 18.930 148.320 19.300 ;
        RECT 150.290 18.965 150.520 35.040 ;
        RECT 150.730 34.720 151.760 34.790 ;
        RECT 150.725 34.490 151.760 34.720 ;
        RECT 150.730 34.410 151.760 34.490 ;
        RECT 151.930 34.440 152.130 35.040 ;
        RECT 152.580 34.820 152.770 34.920 ;
        RECT 153.240 34.820 158.270 37.410 ;
        RECT 152.580 34.440 158.270 34.820 ;
        RECT 150.690 33.930 151.720 34.010 ;
        RECT 151.930 33.980 152.160 34.440 ;
        RECT 150.690 33.700 151.725 33.930 ;
        RECT 150.690 33.630 151.720 33.700 ;
        RECT 151.930 33.650 152.130 33.980 ;
        RECT 150.700 32.830 151.730 33.210 ;
        RECT 150.710 32.060 151.740 32.440 ;
        RECT 150.700 31.270 151.730 31.650 ;
        RECT 150.700 30.480 151.730 30.860 ;
        RECT 150.710 29.670 151.740 30.050 ;
        RECT 150.700 28.890 151.730 29.270 ;
        RECT 150.710 28.090 151.740 28.470 ;
        RECT 150.710 27.300 151.740 27.680 ;
        RECT 150.700 26.520 151.730 26.900 ;
        RECT 150.700 25.730 151.730 26.110 ;
        RECT 150.710 24.940 151.740 25.320 ;
        RECT 150.700 24.150 151.730 24.530 ;
        RECT 150.700 23.370 151.730 23.750 ;
        RECT 150.700 22.580 151.730 22.960 ;
        RECT 150.700 21.790 151.730 22.170 ;
        RECT 150.720 20.980 151.750 21.360 ;
        RECT 150.720 20.200 151.750 20.580 ;
        RECT 150.700 19.420 151.730 19.800 ;
        RECT 137.700 18.660 142.920 18.750 ;
        RECT 137.700 18.085 141.190 18.660 ;
        RECT 142.630 18.610 142.920 18.660 ;
        RECT 143.550 18.610 144.550 18.750 ;
        RECT 145.690 18.500 148.220 18.930 ;
        RECT 150.690 18.920 151.720 19.000 ;
        RECT 151.930 18.965 152.160 33.650 ;
        RECT 150.690 18.690 151.725 18.920 ;
        RECT 150.690 18.620 151.720 18.690 ;
        RECT 152.580 18.520 158.310 34.440 ;
        RECT 147.220 18.190 148.220 18.500 ;
        RECT 152.410 18.450 158.310 18.520 ;
        RECT 147.420 9.410 148.020 18.190 ;
        RECT 149.660 17.930 158.310 18.450 ;
        RECT 148.440 9.410 149.040 9.440 ;
        RECT 147.380 8.810 149.040 9.410 ;
        RECT 148.440 8.780 149.040 8.810 ;
      LAYER via ;
        RECT 140.210 132.070 140.510 132.370 ;
        RECT 156.810 107.820 158.310 109.320 ;
        RECT 140.620 82.460 141.420 83.310 ;
        RECT 142.640 82.470 143.620 83.320 ;
        RECT 140.620 77.830 141.420 78.680 ;
        RECT 142.640 77.840 143.620 78.690 ;
        RECT 141.130 65.440 142.320 71.420 ;
        RECT 143.580 72.510 144.500 73.440 ;
        RECT 143.560 70.100 144.550 71.390 ;
        RECT 143.600 67.950 144.520 68.880 ;
        RECT 143.540 65.520 144.530 66.810 ;
        RECT 143.570 63.380 144.490 64.310 ;
        RECT 143.590 58.050 144.370 58.750 ;
        RECT 142.360 53.350 142.960 53.950 ;
        RECT 142.410 50.300 143.010 50.900 ;
        RECT 150.930 65.800 151.920 66.370 ;
        RECT 154.800 65.800 155.380 66.360 ;
        RECT 150.900 61.210 151.890 61.780 ;
        RECT 154.790 61.220 155.410 61.790 ;
        RECT 143.765 45.680 144.460 47.535 ;
        RECT 143.270 40.780 144.430 41.490 ;
        RECT 148.810 58.050 149.510 58.750 ;
        RECT 150.900 56.630 151.890 57.200 ;
        RECT 154.800 56.620 155.460 57.190 ;
        RECT 150.950 50.950 151.960 51.700 ;
        RECT 150.940 48.660 151.950 49.410 ;
        RECT 150.950 46.410 151.960 47.160 ;
        RECT 150.960 44.100 151.970 44.850 ;
        RECT 154.900 48.680 155.910 49.430 ;
        RECT 150.940 41.820 151.950 42.570 ;
        RECT 154.870 44.100 155.880 44.850 ;
        RECT 150.940 39.530 151.950 40.280 ;
        RECT 150.970 37.210 151.980 37.960 ;
        RECT 154.890 39.570 155.900 40.320 ;
        RECT 140.050 18.600 140.990 35.140 ;
        RECT 143.580 34.700 144.580 35.110 ;
        RECT 143.570 32.420 144.570 32.830 ;
        RECT 143.580 30.120 144.580 30.530 ;
        RECT 143.550 27.790 144.550 28.200 ;
        RECT 143.580 25.540 144.580 25.950 ;
        RECT 143.570 23.250 144.570 23.660 ;
        RECT 143.570 20.950 144.570 21.360 ;
        RECT 143.550 18.660 144.550 19.070 ;
        RECT 145.800 18.920 146.660 32.690 ;
        RECT 147.880 19.670 148.920 32.730 ;
        RECT 150.730 34.460 151.760 34.740 ;
        RECT 150.690 33.680 151.720 33.960 ;
        RECT 150.700 32.880 151.730 33.160 ;
        RECT 150.710 32.110 151.740 32.390 ;
        RECT 150.700 31.320 151.730 31.600 ;
        RECT 150.700 30.530 151.730 30.810 ;
        RECT 150.710 29.720 151.740 30.000 ;
        RECT 150.700 28.940 151.730 29.220 ;
        RECT 150.710 28.140 151.740 28.420 ;
        RECT 150.710 27.350 151.740 27.630 ;
        RECT 150.700 26.570 151.730 26.850 ;
        RECT 150.700 25.780 151.730 26.060 ;
        RECT 150.710 24.990 151.740 25.270 ;
        RECT 150.700 24.200 151.730 24.480 ;
        RECT 150.700 23.420 151.730 23.700 ;
        RECT 150.700 22.630 151.730 22.910 ;
        RECT 150.700 21.840 151.730 22.120 ;
        RECT 150.720 21.030 151.750 21.310 ;
        RECT 150.720 20.250 151.750 20.530 ;
        RECT 150.700 19.470 151.730 19.750 ;
        RECT 154.820 20.140 155.770 33.870 ;
        RECT 150.690 18.670 151.720 18.950 ;
        RECT 148.440 8.810 149.040 9.410 ;
      LAYER met2 ;
        RECT 156.810 147.935 158.310 147.960 ;
        RECT 140.210 147.630 140.510 147.640 ;
        RECT 140.175 147.350 140.545 147.630 ;
        RECT 140.210 132.040 140.510 147.350 ;
        RECT 156.790 146.485 158.330 147.935 ;
        RECT 156.810 107.790 158.310 146.485 ;
        RECT 140.610 83.310 143.670 83.320 ;
        RECT 140.570 82.470 143.670 83.310 ;
        RECT 140.570 82.460 143.650 82.470 ;
        RECT 140.570 78.670 141.470 78.680 ;
        RECT 142.590 78.670 143.670 78.690 ;
        RECT 140.570 77.830 143.670 78.670 ;
        RECT 143.530 72.510 146.330 73.440 ;
        RECT 143.580 72.490 146.330 72.510 ;
        RECT 141.080 71.390 142.370 71.420 ;
        RECT 141.080 70.100 144.600 71.390 ;
        RECT 141.080 70.070 144.560 70.100 ;
        RECT 141.080 66.790 142.370 70.070 ;
        RECT 143.550 68.875 144.570 68.880 ;
        RECT 145.380 68.875 146.330 72.490 ;
        RECT 143.550 67.950 146.330 68.875 ;
        RECT 143.585 67.925 146.330 67.950 ;
        RECT 143.490 66.790 144.580 66.810 ;
        RECT 141.080 65.520 144.580 66.790 ;
        RECT 141.080 65.470 144.570 65.520 ;
        RECT 141.080 65.440 142.370 65.470 ;
        RECT 145.380 64.335 146.330 67.925 ;
        RECT 150.930 66.370 151.920 66.420 ;
        RECT 150.880 66.360 155.390 66.370 ;
        RECT 150.880 65.800 155.430 66.360 ;
        RECT 150.930 65.750 151.920 65.800 ;
        RECT 143.545 64.310 146.330 64.335 ;
        RECT 143.520 63.385 146.330 64.310 ;
        RECT 143.520 63.380 144.540 63.385 ;
        RECT 150.900 61.780 151.890 61.830 ;
        RECT 154.740 61.780 155.460 61.790 ;
        RECT 150.850 61.220 155.460 61.780 ;
        RECT 150.850 61.210 155.170 61.220 ;
        RECT 150.900 61.200 155.170 61.210 ;
        RECT 150.900 61.160 151.890 61.200 ;
        RECT 143.540 58.050 149.560 58.750 ;
        RECT 150.900 57.200 151.890 57.250 ;
        RECT 150.850 57.190 151.890 57.200 ;
        RECT 150.850 56.640 155.510 57.190 ;
        RECT 150.850 56.630 151.940 56.640 ;
        RECT 150.900 56.580 151.890 56.630 ;
        RECT 154.750 56.620 155.510 56.640 ;
        RECT 132.385 53.950 132.935 53.970 ;
        RECT 142.360 53.950 142.960 53.980 ;
        RECT 132.360 53.350 142.960 53.950 ;
        RECT 132.385 53.330 132.935 53.350 ;
        RECT 142.360 53.320 142.960 53.350 ;
        RECT 150.900 51.690 152.010 51.700 ;
        RECT 142.410 50.900 143.010 50.930 ;
        RECT 134.480 50.300 143.010 50.900 ;
        RECT 143.735 50.415 144.505 51.125 ;
        RECT 149.270 50.950 152.010 51.690 ;
        RECT 149.270 50.930 151.990 50.950 ;
        RECT 134.480 8.455 135.080 50.300 ;
        RECT 142.410 50.270 143.010 50.300 ;
        RECT 143.765 47.535 144.475 50.415 ;
        RECT 143.715 45.680 144.510 47.535 ;
        RECT 149.270 47.150 150.220 50.930 ;
        RECT 150.890 49.370 152.000 49.410 ;
        RECT 154.850 49.370 155.960 49.430 ;
        RECT 150.890 48.700 155.960 49.370 ;
        RECT 150.890 48.660 152.000 48.700 ;
        RECT 154.850 48.680 155.960 48.700 ;
        RECT 150.900 47.150 152.010 47.160 ;
        RECT 149.270 46.450 152.010 47.150 ;
        RECT 149.270 42.550 150.220 46.450 ;
        RECT 150.900 46.410 152.010 46.450 ;
        RECT 150.910 44.830 152.020 44.850 ;
        RECT 154.820 44.830 155.930 44.850 ;
        RECT 150.910 44.160 155.930 44.830 ;
        RECT 150.910 44.100 152.020 44.160 ;
        RECT 154.820 44.100 155.930 44.160 ;
        RECT 150.890 42.550 152.000 42.570 ;
        RECT 149.270 41.850 152.000 42.550 ;
        RECT 149.270 41.490 150.220 41.850 ;
        RECT 150.890 41.820 152.000 41.850 ;
        RECT 143.220 40.780 150.220 41.490 ;
        RECT 143.280 40.730 150.220 40.780 ;
        RECT 149.260 37.960 150.220 40.730 ;
        RECT 150.900 40.260 152.000 40.280 ;
        RECT 154.840 40.260 155.950 40.320 ;
        RECT 150.900 39.590 155.950 40.260 ;
        RECT 150.900 39.530 152.000 39.590 ;
        RECT 154.840 39.570 155.950 39.590 ;
        RECT 149.260 37.260 152.030 37.960 ;
        RECT 150.920 37.210 152.030 37.260 ;
        RECT 140.000 35.110 141.040 35.140 ;
        RECT 140.000 34.730 144.630 35.110 ;
        RECT 140.000 30.510 141.040 34.730 ;
        RECT 143.530 34.700 144.630 34.730 ;
        RECT 147.810 34.890 149.140 34.910 ;
        RECT 147.810 34.780 149.360 34.890 ;
        RECT 147.810 34.450 151.810 34.780 ;
        RECT 147.810 33.190 149.360 34.450 ;
        RECT 150.640 33.650 155.850 33.980 ;
        RECT 147.810 32.860 151.780 33.190 ;
        RECT 143.520 32.810 144.620 32.830 ;
        RECT 143.520 32.790 146.140 32.810 ;
        RECT 143.520 32.690 146.670 32.790 ;
        RECT 143.520 32.430 146.710 32.690 ;
        RECT 143.520 32.420 144.620 32.430 ;
        RECT 143.530 30.510 144.630 30.530 ;
        RECT 140.000 30.130 144.630 30.510 ;
        RECT 140.000 25.920 141.040 30.130 ;
        RECT 143.530 30.120 144.630 30.130 ;
        RECT 145.730 28.210 146.710 32.430 ;
        RECT 143.530 28.200 146.710 28.210 ;
        RECT 143.500 27.830 146.710 28.200 ;
        RECT 143.500 27.790 144.600 27.830 ;
        RECT 143.530 25.920 144.630 25.950 ;
        RECT 140.000 25.540 144.630 25.920 ;
        RECT 140.000 21.340 141.040 25.540 ;
        RECT 145.730 23.660 146.710 27.830 ;
        RECT 143.520 23.280 146.710 23.660 ;
        RECT 143.520 23.250 144.620 23.280 ;
        RECT 143.520 21.340 144.620 21.360 ;
        RECT 140.000 20.960 144.620 21.340 ;
        RECT 140.000 18.600 141.040 20.960 ;
        RECT 143.520 20.950 144.620 20.960 ;
        RECT 143.500 19.050 144.600 19.070 ;
        RECT 145.730 19.050 146.710 23.280 ;
        RECT 147.810 31.620 149.360 32.860 ;
        RECT 153.080 32.410 155.850 33.650 ;
        RECT 150.680 32.390 155.850 32.410 ;
        RECT 150.660 32.110 155.850 32.390 ;
        RECT 150.680 32.080 155.850 32.110 ;
        RECT 147.810 31.600 151.760 31.620 ;
        RECT 147.810 31.320 151.780 31.600 ;
        RECT 147.810 31.290 151.760 31.320 ;
        RECT 147.810 30.020 149.360 31.290 ;
        RECT 153.080 30.840 155.850 32.080 ;
        RECT 150.680 30.810 155.850 30.840 ;
        RECT 150.650 30.530 155.850 30.810 ;
        RECT 150.680 30.510 155.850 30.530 ;
        RECT 147.810 29.690 151.790 30.020 ;
        RECT 147.810 28.450 149.360 29.690 ;
        RECT 153.080 29.250 155.850 30.510 ;
        RECT 150.630 28.920 155.850 29.250 ;
        RECT 147.810 28.120 151.790 28.450 ;
        RECT 147.810 26.880 149.360 28.120 ;
        RECT 153.080 27.650 155.850 28.920 ;
        RECT 150.690 27.630 155.850 27.650 ;
        RECT 150.660 27.350 155.850 27.630 ;
        RECT 150.690 27.320 155.850 27.350 ;
        RECT 147.810 26.850 151.770 26.880 ;
        RECT 147.810 26.570 151.780 26.850 ;
        RECT 147.810 26.550 151.770 26.570 ;
        RECT 147.810 25.310 149.360 26.550 ;
        RECT 153.080 26.090 155.850 27.320 ;
        RECT 150.680 26.060 155.850 26.090 ;
        RECT 150.650 25.780 155.850 26.060 ;
        RECT 150.680 25.760 155.850 25.780 ;
        RECT 147.810 24.980 151.790 25.310 ;
        RECT 147.810 23.730 149.360 24.980 ;
        RECT 153.080 24.500 155.850 25.760 ;
        RECT 150.670 24.480 155.850 24.500 ;
        RECT 150.650 24.200 155.850 24.480 ;
        RECT 150.670 24.170 155.850 24.200 ;
        RECT 147.810 23.700 151.750 23.730 ;
        RECT 147.810 23.420 151.780 23.700 ;
        RECT 147.810 23.400 151.750 23.420 ;
        RECT 147.810 22.130 149.360 23.400 ;
        RECT 153.080 22.930 155.850 24.170 ;
        RECT 150.680 22.910 155.850 22.930 ;
        RECT 150.650 22.630 155.850 22.910 ;
        RECT 150.680 22.600 155.850 22.630 ;
        RECT 147.810 22.120 151.770 22.130 ;
        RECT 147.810 21.840 151.780 22.120 ;
        RECT 147.810 21.800 151.770 21.840 ;
        RECT 147.810 20.560 149.360 21.800 ;
        RECT 153.080 21.340 155.850 22.600 ;
        RECT 150.680 21.310 155.850 21.340 ;
        RECT 150.670 21.030 155.850 21.310 ;
        RECT 150.680 21.010 155.850 21.030 ;
        RECT 147.810 20.530 151.750 20.560 ;
        RECT 147.810 20.250 151.800 20.530 ;
        RECT 147.810 20.230 151.750 20.250 ;
        RECT 147.810 19.490 149.360 20.230 ;
        RECT 153.080 19.780 155.850 21.010 ;
        RECT 150.690 19.750 155.850 19.780 ;
        RECT 143.500 18.920 146.710 19.050 ;
        RECT 148.500 18.970 149.360 19.490 ;
        RECT 150.650 19.470 155.850 19.750 ;
        RECT 150.690 19.450 155.850 19.470 ;
        RECT 153.080 19.400 155.850 19.450 ;
        RECT 143.500 18.670 146.670 18.920 ;
        RECT 143.500 18.660 144.600 18.670 ;
        RECT 145.730 18.610 146.670 18.670 ;
        RECT 148.500 18.640 151.780 18.970 ;
        RECT 148.500 18.140 149.360 18.640 ;
        RECT 151.075 9.410 151.625 9.430 ;
        RECT 148.410 8.810 151.650 9.410 ;
        RECT 151.075 8.790 151.625 8.810 ;
        RECT 134.460 7.905 135.100 8.455 ;
        RECT 134.480 7.880 135.080 7.905 ;
      LAYER via2 ;
        RECT 140.220 147.350 140.500 147.630 ;
        RECT 156.835 146.485 158.285 147.935 ;
        RECT 132.385 53.375 132.935 53.925 ;
        RECT 151.075 8.835 151.625 9.385 ;
        RECT 134.505 7.905 135.055 8.455 ;
      LAYER met3 ;
        RECT 15.905 214.660 17.395 214.685 ;
        RECT 15.900 213.160 158.310 214.660 ;
        RECT 15.905 213.135 17.395 213.160 ;
        RECT 140.170 156.490 140.550 156.810 ;
        RECT 140.210 147.655 140.510 156.490 ;
        RECT 140.195 147.325 140.525 147.655 ;
        RECT 156.810 146.460 158.310 213.160 ;
        RECT 119.905 53.950 120.495 53.975 ;
        RECT 119.900 53.350 132.960 53.950 ;
        RECT 119.905 53.325 120.495 53.350 ;
        RECT 151.050 8.810 157.160 9.410 ;
        RECT 134.480 6.015 135.080 8.480 ;
        RECT 156.560 6.715 157.160 8.810 ;
        RECT 156.535 6.125 157.185 6.715 ;
        RECT 156.560 6.120 157.160 6.125 ;
        RECT 134.455 5.425 135.105 6.015 ;
        RECT 134.480 5.420 135.080 5.425 ;
      LAYER via3 ;
        RECT 15.905 213.165 17.395 214.655 ;
        RECT 140.200 156.490 140.520 156.810 ;
        RECT 119.905 53.355 120.495 53.945 ;
        RECT 156.565 6.125 157.155 6.715 ;
        RECT 134.485 5.425 135.075 6.015 ;
      LAYER met4 ;
        RECT 3.990 219.750 4.290 224.760 ;
        RECT 7.670 219.750 7.970 224.760 ;
        RECT 11.350 219.750 11.650 224.760 ;
        RECT 15.030 219.750 15.330 224.760 ;
        RECT 18.710 219.750 19.010 224.760 ;
        RECT 22.390 219.750 22.690 224.760 ;
        RECT 26.070 219.750 26.370 224.760 ;
        RECT 29.750 219.750 30.050 224.760 ;
        RECT 33.430 219.750 33.730 224.760 ;
        RECT 37.110 219.750 37.410 224.760 ;
        RECT 40.790 219.750 41.090 224.760 ;
        RECT 44.470 219.750 44.770 224.760 ;
        RECT 48.150 219.750 48.450 224.760 ;
        RECT 3.990 219.450 49.000 219.750 ;
        RECT 51.830 219.720 52.130 224.760 ;
        RECT 55.510 219.720 55.810 224.760 ;
        RECT 59.190 219.720 59.490 224.760 ;
        RECT 62.870 219.720 63.170 224.760 ;
        RECT 66.550 219.720 66.850 224.760 ;
        RECT 70.230 219.720 70.530 224.760 ;
        RECT 73.910 219.720 74.210 224.760 ;
        RECT 77.590 219.720 77.890 224.760 ;
        RECT 81.270 219.720 81.570 224.760 ;
        RECT 84.950 219.720 85.250 224.760 ;
        RECT 88.630 219.720 88.930 224.760 ;
        RECT 50.500 219.420 140.510 219.720 ;
        RECT 2.500 213.160 17.400 214.660 ;
        RECT 140.210 156.815 140.510 219.420 ;
        RECT 140.195 156.485 140.525 156.815 ;
        RECT 112.400 53.350 120.500 53.950 ;
        RECT 112.400 1.000 113.000 53.350 ;
        RECT 134.480 1.000 135.080 6.020 ;
        RECT 156.560 1.000 157.160 6.720 ;
  END
END tt_um_argunda_tiny_opamp
END LIBRARY

