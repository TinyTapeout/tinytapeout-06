VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_lisa
  CLASS BLOCK ;
  FOREIGN tt_um_lisa ;
  ORIGIN 0.000 0.000 ;
  SIZE 1030.400 BY 225.760 ;
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 258.680 11.880 260.280 144.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 105.080 11.880 106.680 144.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 1026.680 2.480 1028.280 223.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 873.080 2.480 874.680 223.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 719.480 2.480 721.080 223.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 565.880 2.480 567.480 223.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 412.280 2.480 413.880 223.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 258.680 144.120 260.280 223.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 105.080 144.120 106.680 223.280 ;
    END
  END VGND
  PIN VPWR
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 335.480 11.880 337.080 144.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 181.880 11.880 183.480 144.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 28.280 11.880 29.880 144.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 949.880 2.480 951.480 223.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 796.280 2.480 797.880 223.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 642.680 2.480 644.280 223.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 489.080 2.480 490.680 223.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 335.480 144.120 337.080 223.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 181.880 144.120 183.480 223.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 28.280 144.120 29.880 223.280 ;
    END
  END VPWR
  PIN clk
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met4 ;
        RECT 154.870 224.760 155.170 225.760 ;
    END
  END clk
  PIN ena
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met4 ;
        RECT 158.550 224.760 158.850 225.760 ;
    END
  END ena
  PIN rst_n
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 151.190 224.760 151.490 225.760 ;
    END
  END rst_n
  PIN ui_in[0]
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 147.510 224.760 147.810 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met4 ;
        RECT 140.150 224.760 140.450 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met4 ;
        RECT 136.470 224.760 136.770 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met4 ;
        RECT 129.110 224.760 129.410 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met4 ;
        RECT 125.430 224.760 125.730 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 118.070 224.760 118.370 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met4 ;
        RECT 114.390 224.760 114.690 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met4 ;
        RECT 107.030 224.760 107.330 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met4 ;
        RECT 103.350 224.760 103.650 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met4 ;
        RECT 95.990 224.760 96.290 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met4 ;
        RECT 92.310 224.760 92.610 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 29.750 224.760 30.050 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 26.070 224.760 26.370 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 22.390 224.760 22.690 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 18.710 224.760 19.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 15.030 224.760 15.330 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 11.350 224.760 11.650 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 7.670 224.760 7.970 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 3.990 224.760 4.290 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 59.190 224.760 59.490 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 51.830 224.760 52.130 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 48.150 224.760 48.450 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 40.790 224.760 41.090 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 37.110 224.760 37.410 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 84.950 224.760 85.250 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 81.270 224.760 81.570 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 73.910 224.760 74.210 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 70.230 224.760 70.530 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 62.870 224.760 63.170 225.760 ;
    END
  END uo_out[7]
  OBS
      LAYER nwell ;
        RECT 2.570 221.625 1027.830 223.230 ;
        RECT 2.570 216.185 1027.830 219.015 ;
        RECT 2.570 210.745 1027.830 213.575 ;
        RECT 2.570 205.305 1027.830 208.135 ;
        RECT 2.570 199.865 1027.830 202.695 ;
        RECT 2.570 194.425 1027.830 197.255 ;
        RECT 2.570 188.985 1027.830 191.815 ;
        RECT 2.570 183.545 1027.830 186.375 ;
        RECT 2.570 178.105 1027.830 180.935 ;
        RECT 2.570 172.665 1027.830 175.495 ;
        RECT 2.570 167.225 1027.830 170.055 ;
        RECT 2.570 161.785 1027.830 164.615 ;
        RECT 2.570 157.570 1027.830 159.175 ;
      LAYER li1 ;
        RECT 2.760 2.635 1027.640 223.125 ;
      LAYER met1 ;
        RECT 2.760 0.040 1028.280 224.020 ;
      LAYER met2 ;
        RECT 2.860 0.010 1028.250 224.925 ;
      LAYER met3 ;
        RECT 3.745 0.175 1028.270 224.905 ;
      LAYER met4 ;
        RECT 4.690 224.360 7.270 224.905 ;
        RECT 8.370 224.360 10.950 224.905 ;
        RECT 12.050 224.360 14.630 224.905 ;
        RECT 15.730 224.360 18.310 224.905 ;
        RECT 19.410 224.360 21.990 224.905 ;
        RECT 23.090 224.360 25.670 224.905 ;
        RECT 26.770 224.360 29.350 224.905 ;
        RECT 30.450 224.360 33.030 224.905 ;
        RECT 34.130 224.360 36.710 224.905 ;
        RECT 37.810 224.360 40.390 224.905 ;
        RECT 41.490 224.360 44.070 224.905 ;
        RECT 45.170 224.360 47.750 224.905 ;
        RECT 48.850 224.360 51.430 224.905 ;
        RECT 52.530 224.360 55.110 224.905 ;
        RECT 56.210 224.360 58.790 224.905 ;
        RECT 59.890 224.360 62.470 224.905 ;
        RECT 63.570 224.360 66.150 224.905 ;
        RECT 67.250 224.360 69.830 224.905 ;
        RECT 70.930 224.360 73.510 224.905 ;
        RECT 74.610 224.360 77.190 224.905 ;
        RECT 78.290 224.360 80.870 224.905 ;
        RECT 81.970 224.360 84.550 224.905 ;
        RECT 85.650 224.360 88.230 224.905 ;
        RECT 89.330 224.360 91.910 224.905 ;
        RECT 93.010 224.360 95.590 224.905 ;
        RECT 96.690 224.360 99.270 224.905 ;
        RECT 100.370 224.360 102.950 224.905 ;
        RECT 104.050 224.360 106.630 224.905 ;
        RECT 107.730 224.360 110.310 224.905 ;
        RECT 111.410 224.360 113.990 224.905 ;
        RECT 115.090 224.360 117.670 224.905 ;
        RECT 118.770 224.360 121.350 224.905 ;
        RECT 122.450 224.360 125.030 224.905 ;
        RECT 126.130 224.360 128.710 224.905 ;
        RECT 129.810 224.360 132.390 224.905 ;
        RECT 133.490 224.360 136.070 224.905 ;
        RECT 137.170 224.360 139.750 224.905 ;
        RECT 140.850 224.360 143.430 224.905 ;
        RECT 144.530 224.360 147.110 224.905 ;
        RECT 148.210 224.360 150.790 224.905 ;
        RECT 151.890 224.360 154.470 224.905 ;
        RECT 155.570 224.360 158.150 224.905 ;
        RECT 159.250 224.360 1000.665 224.905 ;
        RECT 3.975 223.680 1000.665 224.360 ;
        RECT 3.975 11.480 27.880 223.680 ;
        RECT 30.280 11.480 104.680 223.680 ;
        RECT 107.080 11.480 181.480 223.680 ;
        RECT 183.880 11.480 258.280 223.680 ;
        RECT 260.680 11.480 335.080 223.680 ;
        RECT 337.480 11.480 411.880 223.680 ;
        RECT 3.975 2.080 411.880 11.480 ;
        RECT 414.280 2.080 488.680 223.680 ;
        RECT 491.080 2.080 565.480 223.680 ;
        RECT 567.880 2.080 642.280 223.680 ;
        RECT 644.680 2.080 719.080 223.680 ;
        RECT 721.480 2.080 795.880 223.680 ;
        RECT 798.280 2.080 872.680 223.680 ;
        RECT 875.080 2.080 949.480 223.680 ;
        RECT 951.880 2.080 1000.665 223.680 ;
        RECT 3.975 0.855 1000.665 2.080 ;
  END
END tt_um_lisa
END LIBRARY

