VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_rejunity_current_cmp
  CLASS BLOCK ;
  FOREIGN tt_um_rejunity_current_cmp ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 154.870 224.760 155.170 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 158.550 224.760 158.850 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 151.190 224.760 151.490 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.639000 ;
    PORT
      LAYER met4 ;
        RECT 156.560 0.000 157.160 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.781000 ;
    PORT
      LAYER met4 ;
        RECT 134.480 0.000 135.080 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 112.400 0.000 113.000 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 90.320 0.000 90.920 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 68.240 0.000 68.840 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 46.160 0.000 46.760 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 24.080 0.000 24.680 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 2.000 0.000 2.600 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 147.510 224.760 147.810 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 140.150 224.760 140.450 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 136.470 224.760 136.770 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 129.110 224.760 129.410 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 125.430 224.760 125.730 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.070 224.760 118.370 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 114.390 224.760 114.690 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.030 224.760 107.330 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 103.350 224.760 103.650 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 95.990 224.760 96.290 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 92.310 224.760 92.610 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 12.974000 ;
    PORT
      LAYER met4 ;
        RECT 29.750 224.760 30.050 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 12.974000 ;
    PORT
      LAYER met4 ;
        RECT 26.070 224.760 26.370 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 12.974000 ;
    PORT
      LAYER met4 ;
        RECT 22.390 224.760 22.690 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 12.974000 ;
    PORT
      LAYER met4 ;
        RECT 18.710 224.760 19.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 12.974000 ;
    PORT
      LAYER met4 ;
        RECT 15.030 224.760 15.330 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 12.974000 ;
    PORT
      LAYER met4 ;
        RECT 11.350 224.760 11.650 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 12.974000 ;
    PORT
      LAYER met4 ;
        RECT 7.670 224.760 7.970 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 12.974000 ;
    PORT
      LAYER met4 ;
        RECT 3.990 224.760 4.290 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 12.974000 ;
    PORT
      LAYER met4 ;
        RECT 59.190 224.760 59.490 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 12.974000 ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 12.974000 ;
    PORT
      LAYER met4 ;
        RECT 51.830 224.760 52.130 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 12.974000 ;
    PORT
      LAYER met4 ;
        RECT 48.150 224.760 48.450 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 12.974000 ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 12.974000 ;
    PORT
      LAYER met4 ;
        RECT 40.790 224.760 41.090 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 12.974000 ;
    PORT
      LAYER met4 ;
        RECT 37.110 224.760 37.410 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 12.974000 ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 12.974000 ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 12.974000 ;
    PORT
      LAYER met4 ;
        RECT 84.950 224.760 85.250 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 12.974000 ;
    PORT
      LAYER met4 ;
        RECT 81.270 224.760 81.570 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 12.974000 ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 12.974000 ;
    PORT
      LAYER met4 ;
        RECT 73.910 224.760 74.210 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 12.974000 ;
    PORT
      LAYER met4 ;
        RECT 70.230 224.760 70.530 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 12.974000 ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 12.974000 ;
    PORT
      LAYER met4 ;
        RECT 62.870 224.760 63.170 225.760 ;
    END
  END uo_out[7]
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 2.500 220.760 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 49.000 5.000 50.500 220.760 ;
    END
  END VGND
  OBS
      LAYER nwell ;
        RECT 108.300 209.050 131.800 210.950 ;
        RECT 118.050 204.850 123.300 206.750 ;
        RECT 64.350 194.850 68.000 196.750 ;
        RECT 108.300 196.100 131.800 198.000 ;
      LAYER li1 ;
        RECT 105.700 210.450 133.950 210.850 ;
        RECT 109.000 209.250 109.300 210.450 ;
        RECT 109.650 209.050 109.850 210.250 ;
        RECT 110.200 209.250 110.500 210.450 ;
        RECT 110.850 209.050 111.050 210.250 ;
        RECT 111.400 209.250 111.700 210.450 ;
        RECT 112.050 209.050 112.250 210.250 ;
        RECT 112.600 209.250 112.900 210.450 ;
        RECT 113.250 209.050 113.450 210.250 ;
        RECT 113.800 209.250 114.100 210.450 ;
        RECT 114.450 209.050 114.650 210.250 ;
        RECT 115.000 209.250 115.300 210.450 ;
        RECT 115.650 209.050 115.850 210.250 ;
        RECT 116.200 209.250 116.500 210.450 ;
        RECT 116.850 209.050 117.050 210.250 ;
        RECT 117.400 209.250 117.700 210.450 ;
        RECT 118.050 209.050 118.250 210.250 ;
        RECT 118.900 209.250 119.300 210.450 ;
        RECT 108.900 208.650 119.450 209.050 ;
        RECT 105.750 208.000 107.750 208.400 ;
        RECT 109.050 208.250 109.450 208.450 ;
        RECT 107.350 207.400 107.750 208.000 ;
        RECT 109.000 207.400 109.300 208.000 ;
        RECT 109.650 207.600 109.850 208.650 ;
        RECT 110.250 208.250 110.650 208.450 ;
        RECT 110.200 207.400 110.500 208.000 ;
        RECT 110.850 207.600 111.050 208.650 ;
        RECT 111.450 208.250 111.850 208.450 ;
        RECT 111.400 207.400 111.700 208.000 ;
        RECT 112.050 207.600 112.250 208.650 ;
        RECT 112.650 208.250 113.050 208.450 ;
        RECT 112.600 207.400 112.900 208.000 ;
        RECT 113.250 207.600 113.450 208.650 ;
        RECT 113.850 208.250 114.250 208.450 ;
        RECT 113.800 207.400 114.100 208.000 ;
        RECT 114.450 207.600 114.650 208.650 ;
        RECT 115.050 208.250 115.450 208.450 ;
        RECT 115.000 207.400 115.300 208.000 ;
        RECT 115.650 207.600 115.850 208.650 ;
        RECT 116.250 208.250 116.650 208.450 ;
        RECT 116.200 207.400 116.500 208.000 ;
        RECT 116.850 207.600 117.050 208.650 ;
        RECT 118.050 208.550 119.450 208.650 ;
        RECT 117.450 208.250 117.850 208.450 ;
        RECT 117.400 207.400 117.700 208.000 ;
        RECT 118.050 207.600 118.250 208.550 ;
        RECT 119.650 208.000 120.050 210.250 ;
        RECT 122.000 209.250 122.300 210.450 ;
        RECT 122.050 208.750 122.450 209.050 ;
        RECT 121.100 208.550 121.650 208.650 ;
        RECT 122.650 208.550 122.850 210.250 ;
        RECT 123.200 209.250 123.500 210.450 ;
        RECT 123.250 208.750 123.650 209.050 ;
        RECT 123.850 208.550 124.050 210.250 ;
        RECT 124.400 209.250 124.700 210.450 ;
        RECT 124.450 208.750 124.850 209.050 ;
        RECT 125.050 208.550 125.250 210.250 ;
        RECT 125.600 209.250 125.900 210.450 ;
        RECT 125.650 208.750 126.050 209.050 ;
        RECT 126.250 208.550 126.450 210.250 ;
        RECT 126.800 209.250 127.100 210.450 ;
        RECT 126.850 208.750 127.250 209.050 ;
        RECT 127.450 208.550 127.650 210.250 ;
        RECT 128.000 209.250 128.300 210.450 ;
        RECT 128.050 208.750 128.450 209.050 ;
        RECT 128.650 208.550 128.850 210.250 ;
        RECT 129.200 209.250 129.500 210.450 ;
        RECT 129.250 208.750 129.650 209.050 ;
        RECT 129.850 208.550 130.050 210.250 ;
        RECT 130.400 209.250 130.700 210.450 ;
        RECT 130.450 208.750 130.850 209.050 ;
        RECT 131.050 208.550 131.250 210.250 ;
        RECT 121.100 208.200 131.250 208.550 ;
        RECT 119.650 207.600 120.900 208.000 ;
        RECT 121.250 207.400 121.650 208.000 ;
        RECT 122.100 207.400 122.300 208.000 ;
        RECT 122.650 207.600 122.850 208.200 ;
        RECT 123.200 207.400 123.500 208.000 ;
        RECT 123.850 207.600 124.050 208.200 ;
        RECT 124.500 207.400 124.700 208.000 ;
        RECT 125.050 207.600 125.250 208.200 ;
        RECT 125.600 207.400 125.900 208.000 ;
        RECT 126.250 207.600 126.450 208.200 ;
        RECT 126.900 207.400 127.100 208.000 ;
        RECT 127.450 207.600 127.650 208.200 ;
        RECT 128.000 207.400 128.300 208.000 ;
        RECT 128.650 207.600 128.850 208.200 ;
        RECT 129.300 207.400 129.500 208.000 ;
        RECT 129.850 207.600 130.050 208.200 ;
        RECT 130.400 207.400 130.700 208.000 ;
        RECT 131.050 207.600 131.250 208.200 ;
        RECT 107.350 207.000 132.700 207.400 ;
        RECT 105.700 206.250 131.700 206.650 ;
        RECT 118.350 203.350 118.550 206.050 ;
        RECT 118.750 203.550 118.950 206.250 ;
        RECT 119.300 204.800 119.500 206.050 ;
        RECT 120.300 205.050 120.600 206.250 ;
        RECT 120.950 204.800 121.250 206.050 ;
        RECT 121.600 205.050 121.900 206.250 ;
        RECT 119.300 204.600 120.700 204.800 ;
        RECT 120.950 204.600 122.000 204.800 ;
        RECT 122.250 204.600 122.550 206.050 ;
        RECT 119.300 203.550 119.500 204.600 ;
        RECT 120.950 204.400 121.250 204.600 ;
        RECT 119.700 204.200 121.250 204.400 ;
        RECT 120.300 203.350 120.600 203.950 ;
        RECT 120.950 203.550 121.250 204.200 ;
        RECT 122.250 204.350 131.600 204.600 ;
        RECT 121.600 203.350 121.900 203.950 ;
        RECT 122.250 203.550 122.550 204.350 ;
        RECT 132.300 203.350 132.700 207.000 ;
        RECT 105.700 202.950 132.700 203.350 ;
        RECT 105.700 197.500 133.950 197.900 ;
        RECT 63.540 196.250 67.750 196.650 ;
        RECT 109.000 196.300 109.300 197.500 ;
        RECT 64.650 193.350 64.850 196.050 ;
        RECT 65.050 193.550 65.250 196.250 ;
        RECT 65.600 194.800 65.800 196.050 ;
        RECT 66.600 195.050 66.900 196.250 ;
        RECT 109.650 196.100 109.850 197.300 ;
        RECT 110.200 196.300 110.500 197.500 ;
        RECT 110.850 196.100 111.050 197.300 ;
        RECT 111.400 196.300 111.700 197.500 ;
        RECT 112.050 196.100 112.250 197.300 ;
        RECT 112.600 196.300 112.900 197.500 ;
        RECT 113.250 196.100 113.450 197.300 ;
        RECT 113.800 196.300 114.100 197.500 ;
        RECT 114.450 196.100 114.650 197.300 ;
        RECT 115.000 196.300 115.300 197.500 ;
        RECT 115.650 196.100 115.850 197.300 ;
        RECT 116.200 196.300 116.500 197.500 ;
        RECT 116.850 196.100 117.050 197.300 ;
        RECT 117.400 196.300 117.700 197.500 ;
        RECT 118.050 196.100 118.250 197.300 ;
        RECT 118.900 196.300 119.300 197.500 ;
        RECT 65.600 194.600 67.000 194.800 ;
        RECT 67.250 194.600 67.550 196.050 ;
        RECT 108.900 195.700 119.450 196.100 ;
        RECT 71.050 194.600 71.300 195.450 ;
        RECT 109.050 195.300 109.450 195.500 ;
        RECT 65.600 193.550 65.800 194.600 ;
        RECT 67.250 194.400 68.090 194.600 ;
        RECT 70.700 194.400 71.300 194.600 ;
        RECT 109.000 194.450 109.300 195.050 ;
        RECT 109.650 194.650 109.850 195.700 ;
        RECT 110.250 195.300 110.650 195.500 ;
        RECT 110.200 194.450 110.500 195.050 ;
        RECT 110.850 194.650 111.050 195.700 ;
        RECT 111.450 195.300 111.850 195.500 ;
        RECT 111.400 194.450 111.700 195.050 ;
        RECT 112.050 194.650 112.250 195.700 ;
        RECT 112.650 195.300 113.050 195.500 ;
        RECT 112.600 194.450 112.900 195.050 ;
        RECT 113.250 194.650 113.450 195.700 ;
        RECT 113.850 195.300 114.250 195.500 ;
        RECT 113.800 194.450 114.100 195.050 ;
        RECT 114.450 194.650 114.650 195.700 ;
        RECT 115.050 195.300 115.450 195.500 ;
        RECT 115.000 194.450 115.300 195.050 ;
        RECT 115.650 194.650 115.850 195.700 ;
        RECT 116.250 195.300 116.650 195.500 ;
        RECT 116.200 194.450 116.500 195.050 ;
        RECT 116.850 194.650 117.050 195.700 ;
        RECT 118.050 195.600 119.450 195.700 ;
        RECT 117.450 195.300 117.850 195.500 ;
        RECT 117.400 194.450 117.700 195.050 ;
        RECT 118.050 194.650 118.250 195.600 ;
        RECT 119.650 195.050 120.050 197.300 ;
        RECT 122.000 196.300 122.300 197.500 ;
        RECT 122.050 195.800 122.450 196.100 ;
        RECT 121.100 195.600 121.650 195.700 ;
        RECT 122.650 195.600 122.850 197.300 ;
        RECT 123.200 196.300 123.500 197.500 ;
        RECT 123.250 195.800 123.650 196.100 ;
        RECT 123.850 195.600 124.050 197.300 ;
        RECT 124.400 196.300 124.700 197.500 ;
        RECT 124.450 195.800 124.850 196.100 ;
        RECT 125.050 195.600 125.250 197.300 ;
        RECT 125.600 196.300 125.900 197.500 ;
        RECT 125.650 195.800 126.050 196.100 ;
        RECT 126.250 195.600 126.450 197.300 ;
        RECT 126.800 196.300 127.100 197.500 ;
        RECT 126.850 195.800 127.250 196.100 ;
        RECT 127.450 195.600 127.650 197.300 ;
        RECT 128.000 196.300 128.300 197.500 ;
        RECT 128.050 195.800 128.450 196.100 ;
        RECT 128.650 195.600 128.850 197.300 ;
        RECT 129.200 196.300 129.500 197.500 ;
        RECT 129.250 195.800 129.650 196.100 ;
        RECT 129.850 195.600 130.050 197.300 ;
        RECT 130.400 196.300 130.700 197.500 ;
        RECT 130.450 195.800 130.850 196.100 ;
        RECT 131.050 195.600 131.250 197.300 ;
        RECT 121.100 195.250 131.250 195.600 ;
        RECT 119.650 194.650 120.900 195.050 ;
        RECT 121.250 194.450 121.650 195.050 ;
        RECT 122.100 194.450 122.300 195.050 ;
        RECT 122.650 194.650 122.850 195.250 ;
        RECT 123.200 194.450 123.500 195.050 ;
        RECT 123.850 194.650 124.050 195.250 ;
        RECT 124.500 194.450 124.700 195.050 ;
        RECT 125.050 194.650 125.250 195.250 ;
        RECT 125.600 194.450 125.900 195.050 ;
        RECT 126.250 194.650 126.450 195.250 ;
        RECT 126.900 194.450 127.100 195.050 ;
        RECT 127.450 194.650 127.650 195.250 ;
        RECT 128.000 194.450 128.300 195.050 ;
        RECT 128.650 194.650 128.850 195.250 ;
        RECT 129.300 194.450 129.500 195.050 ;
        RECT 129.850 194.650 130.050 195.250 ;
        RECT 130.400 194.450 130.700 195.050 ;
        RECT 131.050 194.650 131.250 195.250 ;
        RECT 66.000 194.200 67.550 194.400 ;
        RECT 66.600 193.350 66.900 193.950 ;
        RECT 67.250 193.550 67.550 194.200 ;
        RECT 105.700 194.050 132.700 194.450 ;
        RECT 63.540 192.950 67.750 193.350 ;
      LAYER met1 ;
        RECT 92.150 220.050 92.650 220.550 ;
        RECT 95.850 220.050 96.350 220.550 ;
        RECT 99.550 220.050 100.050 220.550 ;
        RECT 103.250 220.050 103.750 220.550 ;
        RECT 106.950 220.050 107.450 220.550 ;
        RECT 110.650 220.050 111.150 220.550 ;
        RECT 114.350 220.050 114.850 220.550 ;
        RECT 117.950 220.050 118.450 220.550 ;
        RECT 121.750 220.050 122.450 220.550 ;
        RECT 125.450 220.050 125.950 220.550 ;
        RECT 129.150 220.050 129.650 220.550 ;
        RECT 132.850 220.050 133.350 220.550 ;
        RECT 136.550 220.050 137.050 220.550 ;
        RECT 140.250 220.050 140.750 220.550 ;
        RECT 143.950 220.050 144.450 220.550 ;
        RECT 147.650 220.050 148.150 220.550 ;
        RECT 92.350 218.450 92.650 220.050 ;
        RECT 92.350 213.250 92.750 218.450 ;
        RECT 96.050 218.400 96.350 220.050 ;
        RECT 96.000 214.150 96.400 218.400 ;
        RECT 99.750 218.300 100.050 220.050 ;
        RECT 99.700 214.950 100.100 218.300 ;
        RECT 103.450 218.250 103.750 220.050 ;
        RECT 107.150 218.250 107.450 220.050 ;
        RECT 110.850 218.400 111.150 220.050 ;
        RECT 103.400 215.800 103.800 218.250 ;
        RECT 107.100 216.750 107.500 218.250 ;
        RECT 110.800 217.600 111.200 218.400 ;
        RECT 114.550 218.300 114.850 220.050 ;
        RECT 118.150 218.300 118.450 220.050 ;
        RECT 114.550 217.900 116.650 218.300 ;
        RECT 110.800 217.200 115.450 217.600 ;
        RECT 107.100 216.350 114.250 216.750 ;
        RECT 103.400 215.400 113.050 215.800 ;
        RECT 99.700 214.550 111.850 214.950 ;
        RECT 96.000 213.750 110.650 214.150 ;
        RECT 92.350 212.850 109.450 213.250 ;
        RECT 104.400 210.150 106.400 211.150 ;
        RECT 104.400 207.650 106.400 208.650 ;
        RECT 104.400 205.950 106.400 206.950 ;
        RECT 104.350 202.600 106.350 203.600 ;
        RECT 104.400 197.200 106.400 198.200 ;
        RECT 65.945 195.365 66.355 196.870 ;
        RECT 65.950 194.500 66.350 195.365 ;
        RECT 70.840 195.330 72.050 195.600 ;
        RECT 70.850 195.000 72.050 195.330 ;
        RECT 109.050 195.200 109.450 212.850 ;
        RECT 110.250 195.200 110.650 213.750 ;
        RECT 111.450 195.200 111.850 214.550 ;
        RECT 112.650 195.200 113.050 215.400 ;
        RECT 113.850 195.200 114.250 216.350 ;
        RECT 115.050 195.200 115.450 217.200 ;
        RECT 116.250 195.200 116.650 217.900 ;
        RECT 117.450 217.900 118.450 218.300 ;
        RECT 117.450 195.200 117.850 217.900 ;
        RECT 119.650 207.805 120.050 208.000 ;
        RECT 119.645 205.365 120.055 207.805 ;
        RECT 119.650 204.500 120.050 205.365 ;
        RECT 122.050 195.750 122.450 220.050 ;
        RECT 125.650 218.300 125.950 220.050 ;
        RECT 129.350 218.300 129.650 220.050 ;
        RECT 133.050 218.300 133.350 220.050 ;
        RECT 136.750 218.350 137.050 220.050 ;
        RECT 123.250 217.900 125.950 218.300 ;
        RECT 123.250 195.750 123.650 217.900 ;
        RECT 129.250 217.600 129.650 218.300 ;
        RECT 124.450 217.200 129.650 217.600 ;
        RECT 124.450 195.750 124.850 217.200 ;
        RECT 133.000 216.750 133.400 218.300 ;
        RECT 125.650 216.350 133.400 216.750 ;
        RECT 125.650 195.750 126.050 216.350 ;
        RECT 136.700 215.850 137.100 218.350 ;
        RECT 140.450 218.300 140.750 220.050 ;
        RECT 126.850 215.450 137.100 215.850 ;
        RECT 126.850 195.750 127.250 215.450 ;
        RECT 140.350 214.850 140.750 218.300 ;
        RECT 128.050 214.450 140.750 214.850 ;
        RECT 144.150 218.500 144.450 220.050 ;
        RECT 147.850 218.600 148.150 220.050 ;
        RECT 128.050 195.750 128.450 214.450 ;
        RECT 144.150 214.200 144.550 218.500 ;
        RECT 129.250 213.800 144.550 214.200 ;
        RECT 129.250 195.750 129.650 213.800 ;
        RECT 147.850 213.300 148.250 218.600 ;
        RECT 130.450 212.900 148.250 213.300 ;
        RECT 130.450 195.750 130.850 212.900 ;
        RECT 133.250 210.150 135.250 211.150 ;
        RECT 131.000 205.950 133.000 206.950 ;
        RECT 131.200 204.150 132.350 204.750 ;
        RECT 132.050 201.650 133.050 203.650 ;
        RECT 133.250 197.200 135.250 198.200 ;
        RECT 119.650 194.855 120.050 195.050 ;
        RECT 104.350 193.700 106.350 194.700 ;
        RECT 66.350 191.800 70.050 192.400 ;
        RECT 119.645 188.650 120.055 194.855 ;
        RECT 132.050 192.750 133.050 194.750 ;
        RECT 119.550 188.050 120.150 188.650 ;
      LAYER met2 ;
        RECT 92.200 220.600 92.600 221.000 ;
        RECT 95.900 220.600 96.300 221.000 ;
        RECT 99.600 220.600 100.000 221.000 ;
        RECT 103.300 220.600 103.700 221.000 ;
        RECT 107.000 220.600 107.400 221.000 ;
        RECT 110.700 220.600 111.100 221.000 ;
        RECT 114.400 220.600 114.800 221.000 ;
        RECT 118.000 220.600 118.400 221.000 ;
        RECT 121.800 220.600 122.200 221.000 ;
        RECT 125.500 220.600 125.900 221.000 ;
        RECT 129.200 220.600 129.600 221.000 ;
        RECT 132.900 220.600 133.300 221.000 ;
        RECT 136.600 220.600 137.000 221.000 ;
        RECT 140.300 220.600 140.700 221.000 ;
        RECT 144.000 220.600 144.400 221.000 ;
        RECT 147.700 220.600 148.100 221.000 ;
        RECT 92.150 220.050 92.650 220.550 ;
        RECT 95.850 220.050 96.350 220.550 ;
        RECT 99.550 220.050 100.050 220.550 ;
        RECT 103.250 220.050 103.750 220.550 ;
        RECT 106.950 220.050 107.450 220.550 ;
        RECT 110.650 220.050 111.150 220.550 ;
        RECT 114.350 220.050 114.850 220.550 ;
        RECT 117.950 220.050 118.450 220.550 ;
        RECT 121.750 220.050 122.250 220.550 ;
        RECT 125.450 220.050 125.950 220.550 ;
        RECT 129.150 220.050 129.650 220.550 ;
        RECT 132.850 220.050 133.350 220.550 ;
        RECT 136.550 220.050 137.050 220.550 ;
        RECT 140.250 220.050 140.750 220.550 ;
        RECT 143.950 220.050 144.450 220.550 ;
        RECT 147.650 220.050 148.150 220.550 ;
        RECT 103.400 210.150 105.400 211.150 ;
        RECT 134.250 210.150 136.250 211.150 ;
        RECT 103.400 207.650 105.400 208.650 ;
        RECT 103.400 205.950 105.400 206.950 ;
        RECT 132.000 205.950 134.000 206.950 ;
        RECT 131.750 204.150 132.950 204.750 ;
        RECT 103.350 202.600 105.350 203.600 ;
        RECT 132.050 200.650 133.050 202.650 ;
        RECT 103.400 197.200 105.400 198.200 ;
        RECT 134.250 197.200 136.250 198.200 ;
        RECT 71.450 195.000 72.650 195.600 ;
        RECT 103.350 193.700 105.350 194.700 ;
        RECT 69.450 191.800 70.650 192.400 ;
        RECT 132.050 191.750 133.050 193.750 ;
        RECT 119.550 188.050 120.750 188.650 ;
      LAYER met3 ;
        RECT 92.150 220.550 92.650 221.550 ;
        RECT 95.850 220.550 96.350 221.550 ;
        RECT 99.550 220.550 100.050 221.550 ;
        RECT 103.250 220.550 103.750 221.550 ;
        RECT 106.950 220.550 107.450 221.550 ;
        RECT 110.650 220.550 111.150 221.550 ;
        RECT 114.350 220.550 114.850 221.550 ;
        RECT 117.950 220.550 118.450 221.550 ;
        RECT 121.750 220.550 122.250 221.550 ;
        RECT 125.450 220.550 125.950 221.550 ;
        RECT 129.150 220.550 129.650 221.550 ;
        RECT 132.850 220.550 133.350 221.550 ;
        RECT 136.550 220.550 137.050 221.550 ;
        RECT 140.250 220.550 140.750 221.550 ;
        RECT 143.950 220.550 144.450 221.550 ;
        RECT 147.650 220.550 148.150 221.550 ;
        RECT 101.950 211.550 136.550 212.850 ;
        RECT 46.400 211.350 136.550 211.550 ;
        RECT 46.400 210.050 104.400 211.350 ;
        RECT 46.400 207.350 47.900 210.050 ;
        RECT 102.400 207.650 104.400 208.650 ;
        RECT 44.490 205.850 104.400 207.350 ;
        RECT 135.050 207.250 136.550 211.350 ;
        RECT 132.700 206.950 136.550 207.250 ;
        RECT 98.650 198.600 100.150 205.850 ;
        RECT 132.800 205.700 136.550 206.950 ;
        RECT 132.350 204.150 133.550 204.750 ;
        RECT 102.350 202.600 104.350 203.600 ;
        RECT 132.050 199.650 133.050 201.650 ;
        RECT 98.650 197.100 104.400 198.600 ;
        RECT 135.000 197.225 136.550 205.700 ;
        RECT 135.050 197.200 136.550 197.225 ;
        RECT 72.050 195.000 73.250 195.600 ;
        RECT 102.400 193.700 104.350 194.700 ;
        RECT 70.050 191.800 71.250 192.400 ;
        RECT 132.050 190.750 133.050 192.750 ;
        RECT 120.150 188.050 121.350 188.650 ;
      LAYER met4 ;
        RECT 3.990 222.450 4.290 224.760 ;
        RECT 7.670 222.450 7.970 224.760 ;
        RECT 11.350 222.450 11.650 224.760 ;
        RECT 15.030 222.450 15.330 224.760 ;
        RECT 18.710 222.450 19.010 224.760 ;
        RECT 22.390 222.450 22.690 224.760 ;
        RECT 26.070 222.450 26.370 224.760 ;
        RECT 29.750 222.450 30.050 224.760 ;
        RECT 33.430 222.450 33.730 224.760 ;
        RECT 37.110 222.450 37.410 224.760 ;
        RECT 40.790 222.450 41.090 224.760 ;
        RECT 44.470 222.450 44.770 224.760 ;
        RECT 48.150 222.450 48.450 224.760 ;
        RECT 51.830 222.450 52.130 224.760 ;
        RECT 55.510 222.450 55.810 224.760 ;
        RECT 59.190 222.450 59.490 224.760 ;
        RECT 62.870 222.450 63.170 224.760 ;
        RECT 66.550 222.450 66.850 224.760 ;
        RECT 70.230 222.450 70.530 224.760 ;
        RECT 73.910 222.450 74.210 224.760 ;
        RECT 77.590 222.450 77.890 224.760 ;
        RECT 81.270 222.450 81.570 224.760 ;
        RECT 84.950 222.450 85.250 224.760 ;
        RECT 88.630 222.450 88.930 224.760 ;
        RECT 3.990 222.150 88.950 222.450 ;
        RECT 49.600 220.760 49.900 222.150 ;
        RECT 92.310 221.550 92.610 224.760 ;
        RECT 95.990 221.550 96.290 224.760 ;
        RECT 99.670 221.550 99.970 224.760 ;
        RECT 103.350 221.550 103.650 224.760 ;
        RECT 107.030 221.550 107.330 224.760 ;
        RECT 110.710 221.550 111.010 224.760 ;
        RECT 114.390 221.550 114.690 224.760 ;
        RECT 118.070 221.550 118.370 224.760 ;
        RECT 121.750 221.550 122.050 224.760 ;
        RECT 125.430 221.800 125.730 224.760 ;
        RECT 129.110 221.800 129.410 224.760 ;
        RECT 132.790 221.800 133.090 224.760 ;
        RECT 136.470 221.800 136.770 224.760 ;
        RECT 140.150 221.800 140.450 224.760 ;
        RECT 143.830 221.800 144.130 224.760 ;
        RECT 147.510 221.800 147.810 224.760 ;
        RECT 125.430 221.550 125.750 221.800 ;
        RECT 129.110 221.600 129.450 221.800 ;
        RECT 132.790 221.600 133.150 221.800 ;
        RECT 129.150 221.550 129.450 221.600 ;
        RECT 132.850 221.550 133.150 221.600 ;
        RECT 136.470 221.550 136.850 221.800 ;
        RECT 140.150 221.550 140.550 221.800 ;
        RECT 143.830 221.550 144.250 221.800 ;
        RECT 147.510 221.550 147.950 221.800 ;
        RECT 92.150 221.050 92.650 221.550 ;
        RECT 95.850 221.050 96.350 221.550 ;
        RECT 99.550 221.050 100.050 221.550 ;
        RECT 103.250 221.050 103.750 221.550 ;
        RECT 106.950 221.050 107.450 221.550 ;
        RECT 110.650 221.050 111.150 221.550 ;
        RECT 114.350 221.050 114.850 221.550 ;
        RECT 117.950 221.050 118.450 221.550 ;
        RECT 121.750 221.050 122.250 221.550 ;
        RECT 125.450 221.050 125.950 221.550 ;
        RECT 129.150 221.050 129.650 221.550 ;
        RECT 132.850 221.050 133.350 221.550 ;
        RECT 136.470 221.350 137.050 221.550 ;
        RECT 140.150 221.400 140.750 221.550 ;
        RECT 136.550 221.050 137.050 221.350 ;
        RECT 140.250 221.050 140.750 221.400 ;
        RECT 143.830 221.150 144.450 221.550 ;
        RECT 147.510 221.150 148.150 221.550 ;
        RECT 143.950 221.050 144.450 221.150 ;
        RECT 147.650 221.050 148.150 221.150 ;
        RECT 50.500 207.540 103.400 209.040 ;
        RECT 2.500 205.850 45.990 207.350 ;
        RECT 132.950 204.710 133.600 204.750 ;
        RECT 132.950 204.170 157.130 204.710 ;
        RECT 132.950 204.150 133.600 204.170 ;
        RECT 50.500 202.490 103.350 203.990 ;
        RECT 100.900 200.700 102.400 202.490 ;
        RECT 100.900 200.650 133.150 200.700 ;
        RECT 100.900 199.200 133.160 200.650 ;
        RECT 72.650 195.560 73.300 195.600 ;
        RECT 72.650 195.020 74.170 195.560 ;
        RECT 100.900 195.090 102.400 199.200 ;
        RECT 72.650 195.000 73.300 195.020 ;
        RECT 100.900 193.590 103.350 195.090 ;
        RECT 70.650 192.340 72.750 192.400 ;
        RECT 70.650 191.800 74.170 192.340 ;
        RECT 72.740 191.740 74.170 191.800 ;
        RECT 100.900 191.800 102.400 193.590 ;
        RECT 100.900 191.750 133.150 191.800 ;
        RECT 100.900 190.300 133.160 191.750 ;
        RECT 120.750 188.050 135.100 188.650 ;
        RECT 134.500 173.750 135.100 188.050 ;
        RECT 134.480 171.700 135.100 173.750 ;
        RECT 134.480 1.000 135.080 171.700 ;
        RECT 156.590 171.390 157.130 204.170 ;
        RECT 156.595 1.000 157.125 171.390 ;
  END
END tt_um_rejunity_current_cmp
END LIBRARY

