VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_lk_ans_top
  CLASS BLOCK ;
  FOREIGN tt_um_lk_ans_top ;
  ORIGIN 0.000 0.000 ;
  SIZE 334.880 BY 225.760 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 95.080 2.480 96.680 223.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 248.680 2.480 250.280 223.280 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 18.280 2.480 19.880 223.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 171.880 2.480 173.480 223.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 325.480 2.480 327.080 223.280 ;
    END
  END VPWR
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met4 ;
        RECT 154.870 224.760 155.170 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 158.550 224.760 158.850 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 151.190 224.760 151.490 225.760 ;
    END
  END rst_n
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met4 ;
        RECT 147.510 224.760 147.810 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met4 ;
        RECT 140.150 224.760 140.450 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met4 ;
        RECT 136.470 224.760 136.770 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 129.110 224.760 129.410 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 125.430 224.760 125.730 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met4 ;
        RECT 118.070 224.760 118.370 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met4 ;
        RECT 114.390 224.760 114.690 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met4 ;
        RECT 107.030 224.760 107.330 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 103.350 224.760 103.650 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 95.990 224.760 96.290 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 92.310 224.760 92.610 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 29.750 224.760 30.050 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 26.070 224.760 26.370 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 22.390 224.760 22.690 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 18.710 224.760 19.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 15.030 224.760 15.330 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 11.350 224.760 11.650 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 7.670 224.760 7.970 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 3.990 224.760 4.290 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 59.190 224.760 59.490 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 51.830 224.760 52.130 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 48.150 224.760 48.450 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met4 ;
        RECT 40.790 224.760 41.090 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 37.110 224.760 37.410 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met4 ;
        RECT 84.950 224.760 85.250 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met4 ;
        RECT 81.270 224.760 81.570 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 73.910 224.760 74.210 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 70.230 224.760 70.530 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 62.870 224.760 63.170 225.760 ;
    END
  END uo_out[7]
  OBS
      LAYER nwell ;
        RECT 2.570 221.625 332.310 223.230 ;
        RECT 2.570 216.185 332.310 219.015 ;
        RECT 2.570 210.745 332.310 213.575 ;
        RECT 2.570 205.305 332.310 208.135 ;
        RECT 2.570 199.865 332.310 202.695 ;
        RECT 2.570 194.425 332.310 197.255 ;
        RECT 2.570 188.985 332.310 191.815 ;
        RECT 2.570 183.545 332.310 186.375 ;
        RECT 2.570 178.105 332.310 180.935 ;
        RECT 2.570 172.665 332.310 175.495 ;
        RECT 2.570 167.225 332.310 170.055 ;
        RECT 2.570 161.785 332.310 164.615 ;
        RECT 2.570 156.345 332.310 159.175 ;
        RECT 2.570 150.905 332.310 153.735 ;
        RECT 2.570 145.465 332.310 148.295 ;
        RECT 2.570 140.025 332.310 142.855 ;
        RECT 2.570 134.585 332.310 137.415 ;
        RECT 2.570 129.145 332.310 131.975 ;
        RECT 2.570 123.705 332.310 126.535 ;
        RECT 2.570 118.265 332.310 121.095 ;
        RECT 2.570 112.825 332.310 115.655 ;
        RECT 2.570 107.385 332.310 110.215 ;
        RECT 2.570 101.945 332.310 104.775 ;
        RECT 2.570 96.505 332.310 99.335 ;
        RECT 2.570 91.065 332.310 93.895 ;
        RECT 2.570 85.625 332.310 88.455 ;
        RECT 2.570 80.185 332.310 83.015 ;
        RECT 2.570 74.745 332.310 77.575 ;
        RECT 2.570 69.305 332.310 72.135 ;
        RECT 2.570 63.865 332.310 66.695 ;
        RECT 2.570 58.425 332.310 61.255 ;
        RECT 2.570 52.985 332.310 55.815 ;
        RECT 2.570 47.545 332.310 50.375 ;
        RECT 2.570 42.105 332.310 44.935 ;
        RECT 2.570 36.665 332.310 39.495 ;
        RECT 2.570 31.225 332.310 34.055 ;
        RECT 2.570 25.785 332.310 28.615 ;
        RECT 2.570 20.345 332.310 23.175 ;
        RECT 2.570 14.905 332.310 17.735 ;
        RECT 2.570 9.465 332.310 12.295 ;
        RECT 2.570 4.025 332.310 6.855 ;
      LAYER li1 ;
        RECT 2.760 2.635 332.120 223.125 ;
      LAYER met1 ;
        RECT 2.760 2.080 332.120 223.680 ;
      LAYER met2 ;
        RECT 4.230 2.050 330.640 224.245 ;
      LAYER met3 ;
        RECT 3.950 2.555 327.070 224.225 ;
      LAYER met4 ;
        RECT 4.690 224.360 7.270 224.760 ;
        RECT 8.370 224.360 10.950 224.760 ;
        RECT 12.050 224.360 14.630 224.760 ;
        RECT 15.730 224.360 18.310 224.760 ;
        RECT 19.410 224.360 21.990 224.760 ;
        RECT 23.090 224.360 25.670 224.760 ;
        RECT 26.770 224.360 29.350 224.760 ;
        RECT 30.450 224.360 33.030 224.760 ;
        RECT 34.130 224.360 36.710 224.760 ;
        RECT 37.810 224.360 40.390 224.760 ;
        RECT 41.490 224.360 44.070 224.760 ;
        RECT 45.170 224.360 47.750 224.760 ;
        RECT 48.850 224.360 51.430 224.760 ;
        RECT 52.530 224.360 55.110 224.760 ;
        RECT 56.210 224.360 58.790 224.760 ;
        RECT 59.890 224.360 62.470 224.760 ;
        RECT 63.570 224.360 66.150 224.760 ;
        RECT 67.250 224.360 69.830 224.760 ;
        RECT 70.930 224.360 73.510 224.760 ;
        RECT 74.610 224.360 77.190 224.760 ;
        RECT 78.290 224.360 80.870 224.760 ;
        RECT 81.970 224.360 84.550 224.760 ;
        RECT 85.650 224.360 88.230 224.760 ;
        RECT 89.330 224.360 91.910 224.760 ;
        RECT 93.010 224.360 95.590 224.760 ;
        RECT 96.690 224.360 99.270 224.760 ;
        RECT 100.370 224.360 102.950 224.760 ;
        RECT 104.050 224.360 106.630 224.760 ;
        RECT 107.730 224.360 110.310 224.760 ;
        RECT 111.410 224.360 113.990 224.760 ;
        RECT 115.090 224.360 117.670 224.760 ;
        RECT 118.770 224.360 121.350 224.760 ;
        RECT 122.450 224.360 125.030 224.760 ;
        RECT 126.130 224.360 128.710 224.760 ;
        RECT 129.810 224.360 132.390 224.760 ;
        RECT 133.490 224.360 136.070 224.760 ;
        RECT 137.170 224.360 139.750 224.760 ;
        RECT 140.850 224.360 143.430 224.760 ;
        RECT 144.530 224.360 147.110 224.760 ;
        RECT 148.210 224.360 150.790 224.760 ;
        RECT 151.890 224.360 154.470 224.760 ;
        RECT 155.570 224.360 158.150 224.760 ;
        RECT 159.250 224.360 244.425 224.760 ;
        RECT 3.975 223.680 244.425 224.360 ;
        RECT 3.975 40.975 17.880 223.680 ;
        RECT 20.280 40.975 94.680 223.680 ;
        RECT 97.080 40.975 171.480 223.680 ;
        RECT 173.880 40.975 244.425 223.680 ;
  END
END tt_um_lk_ans_top
END LIBRARY

