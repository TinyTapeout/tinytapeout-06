VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_nurirfansyah_alits01
  CLASS BLOCK ;
  FOREIGN tt_um_nurirfansyah_alits01 ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 154.870 224.760 155.170 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 158.550 224.760 158.850 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 151.190 224.760 151.490 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.250000 ;
    PORT
      LAYER met4 ;
        RECT 156.560 0.000 157.160 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 5.000000 ;
    PORT
      LAYER met4 ;
        RECT 134.480 0.000 135.080 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 10.000000 ;
    PORT
      LAYER met4 ;
        RECT 112.400 0.000 113.000 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 90.320 0.000 90.920 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 68.240 0.000 68.840 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 46.160 0.000 46.760 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 24.080 0.000 24.680 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 2.000 0.000 2.600 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 147.510 224.760 147.810 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 140.150 224.760 140.450 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 136.470 224.760 136.770 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 129.110 224.760 129.410 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 125.430 224.760 125.730 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.070 224.760 118.370 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 114.390 224.760 114.690 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.030 224.760 107.330 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 103.350 224.760 103.650 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 95.990 224.760 96.290 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 92.310 224.760 92.610 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 19.000000 ;
    PORT
      LAYER met4 ;
        RECT 29.750 224.760 30.050 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 19.000000 ;
    PORT
      LAYER met4 ;
        RECT 26.070 224.760 26.370 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 19.000000 ;
    PORT
      LAYER met4 ;
        RECT 22.390 224.760 22.690 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 19.000000 ;
    PORT
      LAYER met4 ;
        RECT 18.710 224.760 19.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 19.000000 ;
    PORT
      LAYER met4 ;
        RECT 15.030 224.760 15.330 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 19.000000 ;
    PORT
      LAYER met4 ;
        RECT 11.350 224.760 11.650 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 19.000000 ;
    PORT
      LAYER met4 ;
        RECT 7.670 224.760 7.970 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 19.000000 ;
    PORT
      LAYER met4 ;
        RECT 3.990 224.760 4.290 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 19.000000 ;
    PORT
      LAYER met4 ;
        RECT 59.190 224.760 59.490 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 19.000000 ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 19.000000 ;
    PORT
      LAYER met4 ;
        RECT 51.830 224.760 52.130 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 19.000000 ;
    PORT
      LAYER met4 ;
        RECT 48.150 224.760 48.450 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 19.000000 ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 19.000000 ;
    PORT
      LAYER met4 ;
        RECT 40.790 224.760 41.090 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 19.000000 ;
    PORT
      LAYER met4 ;
        RECT 37.110 224.760 37.410 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 19.000000 ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.250000 ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.250000 ;
    PORT
      LAYER met4 ;
        RECT 84.950 224.760 85.250 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.250000 ;
    PORT
      LAYER met4 ;
        RECT 81.270 224.760 81.570 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.250000 ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.250000 ;
    PORT
      LAYER met4 ;
        RECT 73.910 224.760 74.210 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 19.000000 ;
    PORT
      LAYER met4 ;
        RECT 70.230 224.760 70.530 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 19.000000 ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 19.000000 ;
    PORT
      LAYER met4 ;
        RECT 62.870 224.760 63.170 225.760 ;
    END
  END uo_out[7]
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 2.500 220.760 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 49.000 5.000 50.500 220.760 ;
    END
  END VGND
  OBS
      LAYER nwell ;
        RECT 79.250 199.550 108.500 202.200 ;
        RECT 118.590 31.340 147.840 33.990 ;
      LAYER li1 ;
        RECT 79.250 202.350 108.500 202.700 ;
        RECT 79.750 199.750 79.950 202.350 ;
        RECT 79.450 199.150 80.000 199.550 ;
        RECT 80.200 198.950 80.400 201.750 ;
        RECT 79.550 198.600 80.400 198.950 ;
        RECT 79.450 198.000 80.000 198.400 ;
        RECT 79.750 196.400 79.950 197.800 ;
        RECT 80.200 196.800 80.400 198.600 ;
        RECT 81.100 198.950 81.300 201.750 ;
        RECT 82.400 199.750 82.600 202.350 ;
        RECT 82.850 199.750 83.050 202.350 ;
        RECT 83.150 198.950 83.550 199.500 ;
        RECT 81.100 198.600 81.900 198.950 ;
        RECT 81.100 196.800 81.300 198.600 ;
        RECT 82.400 198.550 83.550 198.950 ;
        RECT 83.150 198.050 83.550 198.550 ;
        RECT 83.750 198.950 83.950 201.750 ;
        RECT 84.650 199.750 84.850 202.350 ;
        RECT 85.600 199.750 85.800 202.350 ;
        RECT 85.300 199.150 85.850 199.550 ;
        RECT 86.050 198.950 86.250 201.750 ;
        RECT 83.750 198.550 84.750 198.950 ;
        RECT 85.400 198.600 86.250 198.950 ;
        RECT 82.400 196.400 82.600 197.800 ;
        RECT 82.850 196.400 83.050 197.800 ;
        RECT 83.750 196.800 83.950 198.550 ;
        RECT 85.300 198.000 85.850 198.400 ;
        RECT 84.650 196.400 84.850 197.800 ;
        RECT 85.600 196.400 85.800 197.800 ;
        RECT 86.050 196.800 86.250 198.600 ;
        RECT 86.950 198.950 87.150 201.750 ;
        RECT 88.250 199.750 88.450 202.350 ;
        RECT 88.700 199.750 88.900 202.350 ;
        RECT 89.000 198.950 89.400 199.500 ;
        RECT 86.950 198.600 87.750 198.950 ;
        RECT 86.950 196.800 87.150 198.600 ;
        RECT 88.250 198.550 89.400 198.950 ;
        RECT 89.000 198.050 89.400 198.550 ;
        RECT 89.600 198.950 89.800 201.750 ;
        RECT 90.500 199.750 90.700 202.350 ;
        RECT 91.450 199.750 91.650 202.350 ;
        RECT 91.150 199.150 91.700 199.550 ;
        RECT 91.900 198.950 92.100 201.750 ;
        RECT 89.600 198.550 90.600 198.950 ;
        RECT 91.250 198.600 92.100 198.950 ;
        RECT 88.250 196.400 88.450 197.800 ;
        RECT 88.700 196.400 88.900 197.800 ;
        RECT 89.600 196.800 89.800 198.550 ;
        RECT 91.150 198.000 91.700 198.400 ;
        RECT 90.500 196.400 90.700 197.800 ;
        RECT 91.450 196.400 91.650 197.800 ;
        RECT 91.900 196.800 92.100 198.600 ;
        RECT 92.800 198.950 93.000 201.750 ;
        RECT 94.100 199.750 94.300 202.350 ;
        RECT 94.550 199.750 94.750 202.350 ;
        RECT 94.850 198.950 95.250 199.500 ;
        RECT 92.800 198.600 93.600 198.950 ;
        RECT 92.800 196.800 93.000 198.600 ;
        RECT 94.100 198.550 95.250 198.950 ;
        RECT 94.850 198.050 95.250 198.550 ;
        RECT 95.450 198.950 95.650 201.750 ;
        RECT 96.350 199.750 96.550 202.350 ;
        RECT 97.300 199.750 97.500 202.350 ;
        RECT 97.000 199.150 97.550 199.550 ;
        RECT 97.750 198.950 97.950 201.750 ;
        RECT 95.450 198.550 96.450 198.950 ;
        RECT 97.100 198.600 97.950 198.950 ;
        RECT 94.100 196.400 94.300 197.800 ;
        RECT 94.550 196.400 94.750 197.800 ;
        RECT 95.450 196.800 95.650 198.550 ;
        RECT 97.000 198.000 97.550 198.400 ;
        RECT 96.350 196.400 96.550 197.800 ;
        RECT 97.300 196.400 97.500 197.800 ;
        RECT 97.750 196.800 97.950 198.600 ;
        RECT 98.650 198.950 98.850 201.750 ;
        RECT 99.950 199.750 100.150 202.350 ;
        RECT 100.400 199.750 100.600 202.350 ;
        RECT 100.700 198.950 101.100 199.500 ;
        RECT 98.650 198.600 99.450 198.950 ;
        RECT 98.650 196.800 98.850 198.600 ;
        RECT 99.950 198.550 101.100 198.950 ;
        RECT 100.700 198.050 101.100 198.550 ;
        RECT 101.300 198.950 101.500 201.750 ;
        RECT 102.200 199.750 102.400 202.350 ;
        RECT 103.150 199.750 103.350 202.350 ;
        RECT 102.850 199.150 103.400 199.550 ;
        RECT 103.600 198.950 103.800 201.750 ;
        RECT 101.300 198.550 102.300 198.950 ;
        RECT 102.950 198.600 103.800 198.950 ;
        RECT 99.950 196.400 100.150 197.800 ;
        RECT 100.400 196.400 100.600 197.800 ;
        RECT 101.300 196.800 101.500 198.550 ;
        RECT 102.850 198.000 103.400 198.400 ;
        RECT 102.200 196.400 102.400 197.800 ;
        RECT 103.150 196.400 103.350 197.800 ;
        RECT 103.600 196.800 103.800 198.600 ;
        RECT 104.500 198.950 104.700 201.750 ;
        RECT 105.800 199.750 106.000 202.350 ;
        RECT 106.250 199.750 106.450 202.350 ;
        RECT 106.550 198.950 106.950 199.500 ;
        RECT 104.500 198.600 105.300 198.950 ;
        RECT 104.500 196.800 104.700 198.600 ;
        RECT 105.800 198.550 106.950 198.950 ;
        RECT 106.550 198.050 106.950 198.550 ;
        RECT 107.150 198.950 107.350 201.750 ;
        RECT 108.050 199.750 108.250 202.350 ;
        RECT 107.150 198.550 108.150 198.950 ;
        RECT 105.800 196.400 106.000 197.800 ;
        RECT 106.250 196.400 106.450 197.800 ;
        RECT 107.150 196.800 107.350 198.550 ;
        RECT 108.050 196.400 108.250 197.800 ;
        RECT 79.250 196.050 108.500 196.400 ;
        RECT 118.590 34.140 147.840 34.490 ;
        RECT 119.090 31.540 119.290 34.140 ;
        RECT 118.790 30.940 119.340 31.340 ;
        RECT 119.540 30.740 119.740 33.540 ;
        RECT 118.890 30.390 119.740 30.740 ;
        RECT 118.790 29.790 119.340 30.190 ;
        RECT 119.090 28.190 119.290 29.590 ;
        RECT 119.540 28.590 119.740 30.390 ;
        RECT 120.440 30.740 120.640 33.540 ;
        RECT 121.740 31.540 121.940 34.140 ;
        RECT 122.190 31.540 122.390 34.140 ;
        RECT 122.490 30.740 122.890 31.290 ;
        RECT 120.440 30.390 121.240 30.740 ;
        RECT 120.440 28.590 120.640 30.390 ;
        RECT 121.740 30.340 122.890 30.740 ;
        RECT 122.490 29.840 122.890 30.340 ;
        RECT 123.090 30.740 123.290 33.540 ;
        RECT 123.990 31.540 124.190 34.140 ;
        RECT 124.940 31.540 125.140 34.140 ;
        RECT 124.640 30.940 125.190 31.340 ;
        RECT 125.390 30.740 125.590 33.540 ;
        RECT 123.090 30.340 124.090 30.740 ;
        RECT 124.740 30.390 125.590 30.740 ;
        RECT 121.740 28.190 121.940 29.590 ;
        RECT 122.190 28.190 122.390 29.590 ;
        RECT 123.090 28.590 123.290 30.340 ;
        RECT 124.640 29.790 125.190 30.190 ;
        RECT 123.990 28.190 124.190 29.590 ;
        RECT 124.940 28.190 125.140 29.590 ;
        RECT 125.390 28.590 125.590 30.390 ;
        RECT 126.290 30.740 126.490 33.540 ;
        RECT 127.590 31.540 127.790 34.140 ;
        RECT 128.040 31.540 128.240 34.140 ;
        RECT 128.340 30.740 128.740 31.290 ;
        RECT 126.290 30.390 127.090 30.740 ;
        RECT 126.290 28.590 126.490 30.390 ;
        RECT 127.590 30.340 128.740 30.740 ;
        RECT 128.340 29.840 128.740 30.340 ;
        RECT 128.940 30.740 129.140 33.540 ;
        RECT 129.840 31.540 130.040 34.140 ;
        RECT 130.790 31.540 130.990 34.140 ;
        RECT 130.490 30.940 131.040 31.340 ;
        RECT 131.240 30.740 131.440 33.540 ;
        RECT 128.940 30.340 129.940 30.740 ;
        RECT 130.590 30.390 131.440 30.740 ;
        RECT 127.590 28.190 127.790 29.590 ;
        RECT 128.040 28.190 128.240 29.590 ;
        RECT 128.940 28.590 129.140 30.340 ;
        RECT 130.490 29.790 131.040 30.190 ;
        RECT 129.840 28.190 130.040 29.590 ;
        RECT 130.790 28.190 130.990 29.590 ;
        RECT 131.240 28.590 131.440 30.390 ;
        RECT 132.140 30.740 132.340 33.540 ;
        RECT 133.440 31.540 133.640 34.140 ;
        RECT 133.890 31.540 134.090 34.140 ;
        RECT 134.190 30.740 134.590 31.290 ;
        RECT 132.140 30.390 132.940 30.740 ;
        RECT 132.140 28.590 132.340 30.390 ;
        RECT 133.440 30.340 134.590 30.740 ;
        RECT 134.190 29.840 134.590 30.340 ;
        RECT 134.790 30.740 134.990 33.540 ;
        RECT 135.690 31.540 135.890 34.140 ;
        RECT 136.640 31.540 136.840 34.140 ;
        RECT 136.340 30.940 136.890 31.340 ;
        RECT 137.090 30.740 137.290 33.540 ;
        RECT 134.790 30.340 135.790 30.740 ;
        RECT 136.440 30.390 137.290 30.740 ;
        RECT 133.440 28.190 133.640 29.590 ;
        RECT 133.890 28.190 134.090 29.590 ;
        RECT 134.790 28.590 134.990 30.340 ;
        RECT 136.340 29.790 136.890 30.190 ;
        RECT 135.690 28.190 135.890 29.590 ;
        RECT 136.640 28.190 136.840 29.590 ;
        RECT 137.090 28.590 137.290 30.390 ;
        RECT 137.990 30.740 138.190 33.540 ;
        RECT 139.290 31.540 139.490 34.140 ;
        RECT 139.740 31.540 139.940 34.140 ;
        RECT 140.040 30.740 140.440 31.290 ;
        RECT 137.990 30.390 138.790 30.740 ;
        RECT 137.990 28.590 138.190 30.390 ;
        RECT 139.290 30.340 140.440 30.740 ;
        RECT 140.040 29.840 140.440 30.340 ;
        RECT 140.640 30.740 140.840 33.540 ;
        RECT 141.540 31.540 141.740 34.140 ;
        RECT 142.490 31.540 142.690 34.140 ;
        RECT 142.190 30.940 142.740 31.340 ;
        RECT 142.940 30.740 143.140 33.540 ;
        RECT 140.640 30.340 141.640 30.740 ;
        RECT 142.290 30.390 143.140 30.740 ;
        RECT 139.290 28.190 139.490 29.590 ;
        RECT 139.740 28.190 139.940 29.590 ;
        RECT 140.640 28.590 140.840 30.340 ;
        RECT 142.190 29.790 142.740 30.190 ;
        RECT 141.540 28.190 141.740 29.590 ;
        RECT 142.490 28.190 142.690 29.590 ;
        RECT 142.940 28.590 143.140 30.390 ;
        RECT 143.840 30.740 144.040 33.540 ;
        RECT 145.140 31.540 145.340 34.140 ;
        RECT 145.590 31.540 145.790 34.140 ;
        RECT 145.890 30.740 146.290 31.290 ;
        RECT 143.840 30.390 144.640 30.740 ;
        RECT 143.840 28.590 144.040 30.390 ;
        RECT 145.140 30.340 146.290 30.740 ;
        RECT 145.890 29.840 146.290 30.340 ;
        RECT 146.490 30.740 146.690 33.540 ;
        RECT 147.390 31.540 147.590 34.140 ;
        RECT 146.490 30.340 147.490 30.740 ;
        RECT 145.140 28.190 145.340 29.590 ;
        RECT 145.590 28.190 145.790 29.590 ;
        RECT 146.490 28.590 146.690 30.340 ;
        RECT 147.390 28.190 147.590 29.590 ;
        RECT 118.590 27.840 147.840 28.190 ;
      LAYER met1 ;
        RECT 0.850 202.500 108.500 203.300 ;
        RECT 0.850 201.450 2.600 202.500 ;
        RECT 79.250 202.300 108.500 202.500 ;
        RECT 79.400 199.500 80.050 200.000 ;
        RECT 85.250 199.500 85.900 200.000 ;
        RECT 91.100 199.500 91.750 200.000 ;
        RECT 96.950 199.500 97.600 200.000 ;
        RECT 102.800 199.500 103.450 200.000 ;
        RECT 79.450 199.150 80.000 199.500 ;
        RECT 85.300 199.150 85.850 199.500 ;
        RECT 91.150 199.150 91.700 199.500 ;
        RECT 97.000 199.150 97.550 199.500 ;
        RECT 102.850 199.150 103.400 199.500 ;
        RECT 78.700 198.950 79.250 199.050 ;
        RECT 81.900 198.950 82.950 199.050 ;
        RECT 78.700 198.600 80.200 198.950 ;
        RECT 81.250 198.600 82.950 198.950 ;
        RECT 78.700 198.500 79.250 198.600 ;
        RECT 81.900 198.450 82.950 198.600 ;
        RECT 83.950 198.950 84.850 199.100 ;
        RECT 87.750 198.950 88.800 199.050 ;
        RECT 83.950 198.600 86.050 198.950 ;
        RECT 87.100 198.600 88.800 198.950 ;
        RECT 83.950 198.400 84.850 198.600 ;
        RECT 87.750 198.450 88.800 198.600 ;
        RECT 89.750 198.950 90.650 199.100 ;
        RECT 93.600 198.950 94.650 199.050 ;
        RECT 89.750 198.600 91.900 198.950 ;
        RECT 92.950 198.600 94.650 198.950 ;
        RECT 89.750 198.400 90.650 198.600 ;
        RECT 93.600 198.450 94.650 198.600 ;
        RECT 95.650 198.950 96.550 199.100 ;
        RECT 99.450 198.950 100.500 199.050 ;
        RECT 95.650 198.600 97.750 198.950 ;
        RECT 98.800 198.600 100.500 198.950 ;
        RECT 95.650 198.400 96.550 198.600 ;
        RECT 99.450 198.450 100.500 198.600 ;
        RECT 101.450 198.950 102.350 199.100 ;
        RECT 105.300 198.950 106.350 199.050 ;
        RECT 101.450 198.600 103.600 198.950 ;
        RECT 104.650 198.600 106.350 198.950 ;
        RECT 101.450 198.400 102.350 198.600 ;
        RECT 105.300 198.450 106.350 198.600 ;
        RECT 107.600 198.450 108.200 199.050 ;
        RECT 79.450 198.000 80.000 198.400 ;
        RECT 85.300 198.000 85.850 198.400 ;
        RECT 91.150 198.000 91.700 198.400 ;
        RECT 97.000 198.000 97.550 198.400 ;
        RECT 102.850 198.000 103.400 198.400 ;
        RECT 79.400 197.500 80.050 198.000 ;
        RECT 85.250 197.500 85.900 198.000 ;
        RECT 91.100 197.500 91.750 198.000 ;
        RECT 96.950 197.500 97.600 198.000 ;
        RECT 102.800 197.500 103.450 198.000 ;
        RECT 79.250 196.400 108.500 196.450 ;
        RECT 48.900 195.700 108.500 196.400 ;
        RECT 48.900 194.550 50.600 195.700 ;
        RECT 0.950 34.150 147.850 34.850 ;
        RECT 118.590 34.090 147.840 34.150 ;
        RECT 118.740 31.290 119.390 31.790 ;
        RECT 124.590 31.290 125.240 31.790 ;
        RECT 130.440 31.290 131.090 31.790 ;
        RECT 136.290 31.290 136.940 31.790 ;
        RECT 142.140 31.290 142.790 31.790 ;
        RECT 118.790 30.940 119.340 31.290 ;
        RECT 124.640 30.940 125.190 31.290 ;
        RECT 130.490 30.940 131.040 31.290 ;
        RECT 136.340 30.940 136.890 31.290 ;
        RECT 142.190 30.940 142.740 31.290 ;
        RECT 118.040 30.740 118.590 30.840 ;
        RECT 121.240 30.740 122.290 30.840 ;
        RECT 118.040 30.390 119.540 30.740 ;
        RECT 120.590 30.390 122.290 30.740 ;
        RECT 118.040 30.290 118.590 30.390 ;
        RECT 121.240 30.240 122.290 30.390 ;
        RECT 123.540 30.740 124.140 30.840 ;
        RECT 127.090 30.740 128.140 30.840 ;
        RECT 123.540 30.390 125.390 30.740 ;
        RECT 126.440 30.390 128.140 30.740 ;
        RECT 123.540 30.240 124.140 30.390 ;
        RECT 127.090 30.240 128.140 30.390 ;
        RECT 129.390 30.740 129.990 30.840 ;
        RECT 132.940 30.740 133.990 30.840 ;
        RECT 129.390 30.390 131.240 30.740 ;
        RECT 132.290 30.390 133.990 30.740 ;
        RECT 129.390 30.240 129.990 30.390 ;
        RECT 132.940 30.240 133.990 30.390 ;
        RECT 135.240 30.740 135.840 30.840 ;
        RECT 138.790 30.740 139.840 30.840 ;
        RECT 135.240 30.390 137.090 30.740 ;
        RECT 138.140 30.390 139.840 30.740 ;
        RECT 135.240 30.240 135.840 30.390 ;
        RECT 138.790 30.240 139.840 30.390 ;
        RECT 141.090 30.740 141.690 30.840 ;
        RECT 144.640 30.740 145.690 30.840 ;
        RECT 141.090 30.390 142.940 30.740 ;
        RECT 143.990 30.390 145.690 30.740 ;
        RECT 141.090 30.240 141.690 30.390 ;
        RECT 144.640 30.240 145.690 30.390 ;
        RECT 146.940 30.240 147.540 30.840 ;
        RECT 118.790 29.790 119.340 30.190 ;
        RECT 124.640 29.790 125.190 30.190 ;
        RECT 130.490 29.790 131.040 30.190 ;
        RECT 136.340 29.790 136.890 30.190 ;
        RECT 142.190 29.790 142.740 30.190 ;
        RECT 118.740 29.290 119.390 29.790 ;
        RECT 124.590 29.290 125.240 29.790 ;
        RECT 130.440 29.290 131.090 29.790 ;
        RECT 136.290 29.290 136.940 29.790 ;
        RECT 142.140 29.290 142.790 29.790 ;
        RECT 118.590 28.200 147.840 28.240 ;
        RECT 48.600 27.300 148.500 28.200 ;
      LAYER met2 ;
        RECT 0.850 201.450 2.600 203.300 ;
        RECT 75.100 199.950 75.700 200.000 ;
        RECT 79.400 199.950 80.050 200.000 ;
        RECT 75.100 199.900 80.050 199.950 ;
        RECT 85.250 199.900 85.900 200.000 ;
        RECT 91.100 199.900 91.750 200.000 ;
        RECT 96.950 199.900 97.600 200.000 ;
        RECT 102.800 199.900 103.450 200.000 ;
        RECT 75.100 199.550 107.850 199.900 ;
        RECT 48.900 194.550 50.600 196.400 ;
        RECT 75.100 187.800 75.700 199.550 ;
        RECT 79.400 199.500 80.050 199.550 ;
        RECT 85.250 199.500 85.900 199.550 ;
        RECT 91.100 199.500 91.750 199.550 ;
        RECT 96.950 199.500 97.600 199.550 ;
        RECT 102.800 199.500 103.450 199.550 ;
        RECT 78.150 198.300 79.250 199.100 ;
        RECT 83.950 198.400 84.850 199.100 ;
        RECT 89.750 198.400 90.650 199.100 ;
        RECT 95.650 198.400 96.550 199.100 ;
        RECT 101.450 198.400 102.350 199.100 ;
        RECT 107.600 198.950 108.350 199.050 ;
        RECT 107.550 198.600 108.350 198.950 ;
        RECT 107.600 198.450 108.350 198.600 ;
        RECT 79.400 197.900 80.050 198.000 ;
        RECT 76.800 197.850 80.050 197.900 ;
        RECT 85.250 197.850 85.900 198.000 ;
        RECT 91.100 197.850 91.750 198.000 ;
        RECT 96.950 197.850 97.600 198.000 ;
        RECT 102.800 197.850 103.450 198.000 ;
        RECT 76.800 197.500 103.450 197.850 ;
        RECT 76.800 192.400 77.400 197.500 ;
        RECT 107.750 196.800 108.350 198.450 ;
        RECT 78.050 196.300 108.350 196.800 ;
        RECT 78.050 196.100 79.350 196.300 ;
        RECT 76.800 191.600 117.000 192.400 ;
        RECT 75.100 187.000 113.000 187.800 ;
        RECT 0.950 34.850 2.550 35.550 ;
        RECT 0.950 34.150 4.850 34.850 ;
        RECT 0.950 33.500 2.550 34.150 ;
        RECT 112.050 31.690 119.400 31.800 ;
        RECT 124.590 31.690 125.240 31.790 ;
        RECT 130.440 31.690 131.090 31.790 ;
        RECT 136.290 31.690 136.940 31.790 ;
        RECT 142.140 31.690 142.790 31.790 ;
        RECT 112.050 31.340 147.190 31.690 ;
        RECT 112.050 31.300 119.400 31.340 ;
        RECT 48.600 28.200 50.750 31.300 ;
        RECT 112.050 30.850 113.300 31.300 ;
        RECT 118.740 31.290 119.390 31.300 ;
        RECT 124.590 31.290 125.240 31.340 ;
        RECT 130.440 31.290 131.090 31.340 ;
        RECT 136.290 31.290 136.940 31.340 ;
        RECT 142.140 31.290 142.790 31.340 ;
        RECT 118.040 30.740 118.590 30.840 ;
        RECT 146.900 30.740 157.200 30.850 ;
        RECT 118.040 30.390 157.200 30.740 ;
        RECT 118.040 30.290 118.590 30.390 ;
        RECT 146.900 30.250 157.200 30.390 ;
        RECT 146.900 30.150 148.300 30.250 ;
        RECT 115.600 29.640 120.050 29.800 ;
        RECT 124.590 29.640 125.240 29.790 ;
        RECT 130.440 29.640 131.090 29.790 ;
        RECT 136.290 29.640 136.940 29.790 ;
        RECT 142.140 29.640 142.790 29.790 ;
        RECT 156.250 29.700 157.200 30.250 ;
        RECT 115.600 29.300 142.790 29.640 ;
        RECT 115.600 28.900 116.850 29.300 ;
        RECT 118.740 29.290 142.790 29.300 ;
        RECT 48.600 27.300 57.600 28.200 ;
        RECT 48.600 25.300 50.750 27.300 ;
      LAYER met3 ;
        RECT 88.500 221.850 108.350 222.450 ;
        RECT 84.950 220.600 102.150 221.250 ;
        RECT 81.200 219.100 96.350 219.750 ;
        RECT 77.450 217.150 90.450 217.700 ;
        RECT 73.750 214.850 84.650 215.550 ;
        RECT 0.850 201.450 2.600 203.300 ;
        RECT 84.150 199.100 84.650 214.850 ;
        RECT 89.950 199.100 90.450 217.150 ;
        RECT 95.850 199.100 96.350 219.100 ;
        RECT 101.650 199.100 102.150 220.600 ;
        RECT 78.150 198.300 79.250 199.100 ;
        RECT 83.950 198.400 84.850 199.100 ;
        RECT 89.750 198.400 90.650 199.100 ;
        RECT 95.650 198.400 96.550 199.100 ;
        RECT 101.450 198.400 102.350 199.100 ;
        RECT 107.850 199.050 108.350 221.850 ;
        RECT 107.750 198.450 108.350 199.050 ;
        RECT 78.150 196.800 78.650 198.300 ;
        RECT 107.850 197.950 108.350 198.450 ;
        RECT 48.900 194.550 50.600 196.400 ;
        RECT 78.050 196.100 79.350 196.800 ;
        RECT 1.000 33.350 2.500 35.700 ;
        RECT 48.900 25.150 50.600 31.350 ;
        RECT 112.000 1.550 113.100 187.900 ;
        RECT 115.650 12.950 116.700 192.450 ;
        RECT 115.650 12.200 135.100 12.950 ;
        RECT 115.850 12.150 135.100 12.200 ;
        RECT 134.350 2.900 135.100 12.150 ;
        RECT 156.450 3.100 157.100 31.000 ;
        RECT 134.350 1.550 135.200 2.900 ;
        RECT 156.450 1.650 157.300 3.100 ;
      LAYER met4 ;
        RECT 3.990 223.500 4.290 224.760 ;
        RECT 7.670 223.500 7.970 224.760 ;
        RECT 11.350 223.500 11.650 224.760 ;
        RECT 15.030 223.500 15.330 224.760 ;
        RECT 18.710 223.500 19.010 224.760 ;
        RECT 22.390 223.500 22.690 224.760 ;
        RECT 26.070 223.500 26.370 224.760 ;
        RECT 29.750 223.500 30.050 224.760 ;
        RECT 33.430 223.500 33.730 224.760 ;
        RECT 37.110 223.500 37.410 224.760 ;
        RECT 40.790 223.500 41.090 224.760 ;
        RECT 44.470 223.500 44.770 224.760 ;
        RECT 48.150 223.500 48.450 224.760 ;
        RECT 51.830 223.500 52.130 224.760 ;
        RECT 55.510 223.500 55.810 224.760 ;
        RECT 59.190 223.500 59.490 224.760 ;
        RECT 62.870 223.500 63.170 224.760 ;
        RECT 66.550 223.500 66.850 224.760 ;
        RECT 70.230 223.500 70.530 224.760 ;
        RECT 73.910 223.650 74.210 224.760 ;
        RECT 77.590 223.800 77.890 224.760 ;
        RECT 3.600 222.600 70.530 223.500 ;
        RECT 49.300 220.760 50.200 222.600 ;
        RECT 73.750 214.800 74.400 223.650 ;
        RECT 77.500 217.800 78.000 223.800 ;
        RECT 81.270 223.650 81.570 224.760 ;
        RECT 84.950 223.650 85.250 224.760 ;
        RECT 88.630 223.700 88.930 224.760 ;
        RECT 81.200 219.100 81.900 223.650 ;
        RECT 84.950 220.600 85.750 223.650 ;
        RECT 88.500 221.850 89.300 223.700 ;
        RECT 77.500 217.150 78.150 217.800 ;
        RECT 112.250 1.550 113.100 2.750 ;
        RECT 134.350 1.550 135.200 2.750 ;
        RECT 156.450 1.650 157.300 2.850 ;
        RECT 112.400 1.000 113.000 1.550 ;
        RECT 134.480 1.000 135.080 1.550 ;
        RECT 156.560 1.000 157.160 1.650 ;
  END
END tt_um_nurirfansyah_alits01
END LIBRARY

