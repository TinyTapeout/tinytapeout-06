VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_argunda_tiny_opamp
  CLASS BLOCK ;
  FOREIGN tt_um_argunda_tiny_opamp ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 154.870 224.760 155.170 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 158.550 224.760 158.850 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 151.190 224.760 151.490 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.350000 ;
    PORT
      LAYER met4 ;
        RECT 156.560 0.000 157.160 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.250000 ;
    PORT
      LAYER met4 ;
        RECT 134.480 0.000 135.080 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.250000 ;
    PORT
      LAYER met4 ;
        RECT 112.400 0.000 113.000 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.350000 ;
    PORT
      LAYER met4 ;
        RECT 90.320 0.000 90.920 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.250000 ;
    PORT
      LAYER met4 ;
        RECT 68.240 0.000 68.840 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.250000 ;
    PORT
      LAYER met4 ;
        RECT 46.160 0.000 46.760 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 24.080 0.000 24.680 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 2.000 0.000 2.600 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 147.510 224.760 147.810 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 140.150 224.760 140.450 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 136.470 224.760 136.770 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 129.110 224.760 129.410 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 125.430 224.760 125.730 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.070 224.760 118.370 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 114.390 224.760 114.690 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.030 224.760 107.330 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 103.350 224.760 103.650 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 95.990 224.760 96.290 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 92.310 224.760 92.610 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 44.755798 ;
    PORT
      LAYER met4 ;
        RECT 29.750 224.760 30.050 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 44.755798 ;
    PORT
      LAYER met4 ;
        RECT 26.070 224.760 26.370 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 44.755798 ;
    PORT
      LAYER met4 ;
        RECT 22.390 224.760 22.690 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 44.755798 ;
    PORT
      LAYER met4 ;
        RECT 18.710 224.760 19.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 44.755798 ;
    PORT
      LAYER met4 ;
        RECT 15.030 224.760 15.330 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 44.755798 ;
    PORT
      LAYER met4 ;
        RECT 11.350 224.760 11.650 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 44.755798 ;
    PORT
      LAYER met4 ;
        RECT 7.670 224.760 7.970 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 44.755798 ;
    PORT
      LAYER met4 ;
        RECT 3.990 224.760 4.290 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 44.755798 ;
    PORT
      LAYER met4 ;
        RECT 59.190 224.760 59.490 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 44.755798 ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 44.755798 ;
    PORT
      LAYER met4 ;
        RECT 51.830 224.760 52.130 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 44.755798 ;
    PORT
      LAYER met4 ;
        RECT 48.150 224.760 48.450 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 44.755798 ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 44.755798 ;
    PORT
      LAYER met4 ;
        RECT 40.790 224.760 41.090 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 44.755798 ;
    PORT
      LAYER met4 ;
        RECT 37.110 224.760 37.410 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 44.755798 ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 44.755798 ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 44.755798 ;
    PORT
      LAYER met4 ;
        RECT 84.950 224.760 85.250 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 44.755798 ;
    PORT
      LAYER met4 ;
        RECT 81.270 224.760 81.570 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 44.755798 ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 44.755798 ;
    PORT
      LAYER met4 ;
        RECT 73.910 224.760 74.210 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 44.755798 ;
    PORT
      LAYER met4 ;
        RECT 70.230 224.760 70.530 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 44.755798 ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 44.755798 ;
    PORT
      LAYER met4 ;
        RECT 62.870 224.760 63.170 225.760 ;
    END
  END uo_out[7]
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 2.500 220.760 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 155.860 4.920 157.360 220.680 ;
    END
  END VGND
  OBS
      LAYER nwell ;
        RECT 60.880 34.830 66.730 50.240 ;
      LAYER pwell ;
        RECT 61.590 29.860 65.980 34.460 ;
        RECT 54.850 24.420 65.680 27.520 ;
        RECT 72.510 25.370 75.610 43.070 ;
      LAYER nwell ;
        RECT 77.650 32.760 80.840 50.230 ;
      LAYER pwell ;
        RECT 99.400 41.360 101.410 49.980 ;
        RECT 94.790 37.040 105.620 40.140 ;
      LAYER nwell ;
        RECT 123.110 34.430 128.960 49.840 ;
      LAYER pwell ;
        RECT 123.820 29.460 128.210 34.060 ;
        RECT 117.080 24.020 127.910 27.120 ;
        RECT 134.740 24.970 137.840 42.670 ;
      LAYER nwell ;
        RECT 139.880 32.360 143.070 49.830 ;
      LAYER li1 ;
        RECT 54.840 49.890 84.840 52.430 ;
        RECT 94.360 50.340 106.510 51.780 ;
        RECT 54.840 35.180 61.230 49.890 ;
        RECT 61.955 49.320 62.995 49.490 ;
        RECT 61.570 47.260 61.740 49.260 ;
        RECT 63.210 47.260 63.380 49.260 ;
        RECT 61.955 47.030 62.995 47.200 ;
        RECT 61.570 44.970 61.740 46.970 ;
        RECT 63.210 44.970 63.380 46.970 ;
        RECT 61.955 44.740 62.995 44.910 ;
        RECT 61.570 42.680 61.740 44.680 ;
        RECT 63.210 42.680 63.380 44.680 ;
        RECT 61.955 42.450 62.995 42.620 ;
        RECT 61.570 40.390 61.740 42.390 ;
        RECT 63.210 40.390 63.380 42.390 ;
        RECT 61.955 40.160 62.995 40.330 ;
        RECT 61.570 38.100 61.740 40.100 ;
        RECT 63.210 38.100 63.380 40.100 ;
        RECT 61.955 37.870 62.995 38.040 ;
        RECT 61.570 35.810 61.740 37.810 ;
        RECT 63.210 35.810 63.380 37.810 ;
        RECT 61.955 35.580 62.995 35.750 ;
        RECT 63.720 35.180 63.890 49.890 ;
        RECT 66.380 49.880 84.840 49.890 ;
        RECT 64.615 49.320 65.655 49.490 ;
        RECT 64.230 47.260 64.400 49.260 ;
        RECT 65.870 47.260 66.040 49.260 ;
        RECT 64.615 47.030 65.655 47.200 ;
        RECT 64.230 44.970 64.400 46.970 ;
        RECT 65.870 44.970 66.040 46.970 ;
        RECT 64.615 44.740 65.655 44.910 ;
        RECT 64.230 42.680 64.400 44.680 ;
        RECT 65.870 42.680 66.040 44.680 ;
        RECT 66.380 43.690 78.000 49.880 ;
        RECT 78.725 49.310 79.765 49.480 ;
        RECT 78.340 48.750 78.510 49.250 ;
        RECT 79.980 48.750 80.150 49.250 ;
        RECT 78.725 48.520 79.765 48.690 ;
        RECT 78.340 47.960 78.510 48.460 ;
        RECT 79.980 47.960 80.150 48.460 ;
        RECT 78.725 47.730 79.765 47.900 ;
        RECT 78.340 47.170 78.510 47.670 ;
        RECT 79.980 47.170 80.150 47.670 ;
        RECT 78.725 46.940 79.765 47.110 ;
        RECT 78.340 46.380 78.510 46.880 ;
        RECT 79.980 46.380 80.150 46.880 ;
        RECT 78.725 46.150 79.765 46.320 ;
        RECT 78.340 45.590 78.510 46.090 ;
        RECT 79.980 45.590 80.150 46.090 ;
        RECT 78.725 45.360 79.765 45.530 ;
        RECT 78.340 44.800 78.510 45.300 ;
        RECT 79.980 44.800 80.150 45.300 ;
        RECT 78.725 44.570 79.765 44.740 ;
        RECT 78.340 44.010 78.510 44.510 ;
        RECT 79.980 44.010 80.150 44.510 ;
        RECT 78.725 43.780 79.765 43.950 ;
        RECT 64.615 42.450 65.655 42.620 ;
        RECT 64.230 40.390 64.400 42.390 ;
        RECT 65.870 40.390 66.040 42.390 ;
        RECT 64.615 40.160 65.655 40.330 ;
        RECT 64.230 38.100 64.400 40.100 ;
        RECT 65.870 38.100 66.040 40.100 ;
        RECT 64.615 37.870 65.655 38.040 ;
        RECT 64.230 35.810 64.400 37.810 ;
        RECT 65.870 35.810 66.040 37.810 ;
        RECT 64.615 35.580 65.655 35.750 ;
        RECT 66.380 35.180 71.810 43.690 ;
        RECT 54.840 34.810 71.810 35.180 ;
        RECT 72.690 42.720 75.430 42.890 ;
        RECT 54.840 34.800 71.660 34.810 ;
        RECT 72.690 34.280 72.860 42.720 ;
        RECT 73.540 42.150 74.580 42.320 ;
        RECT 73.200 40.090 73.370 42.090 ;
        RECT 74.750 40.090 74.920 42.090 ;
        RECT 73.540 39.860 74.580 40.030 ;
        RECT 73.200 37.800 73.370 39.800 ;
        RECT 74.750 37.800 74.920 39.800 ;
        RECT 73.540 37.570 74.580 37.740 ;
        RECT 73.200 35.510 73.370 37.510 ;
        RECT 74.750 35.510 74.920 37.510 ;
        RECT 73.540 35.280 74.580 35.450 ;
        RECT 54.840 34.110 72.860 34.280 ;
        RECT 54.840 30.210 61.940 34.110 ;
        RECT 62.570 33.600 63.070 33.770 ;
        RECT 62.340 30.890 62.510 33.430 ;
        RECT 63.130 30.890 63.300 33.430 ;
        RECT 62.570 30.550 63.070 30.720 ;
        RECT 63.700 30.210 63.870 34.110 ;
        RECT 64.500 33.600 65.000 33.770 ;
        RECT 64.270 30.890 64.440 33.430 ;
        RECT 65.060 30.890 65.230 33.430 ;
        RECT 64.500 30.550 65.000 30.720 ;
        RECT 65.630 30.210 72.860 34.110 ;
        RECT 73.200 33.220 73.370 35.220 ;
        RECT 74.750 33.220 74.920 35.220 ;
        RECT 73.540 32.990 74.580 33.160 ;
        RECT 73.200 30.930 73.370 32.930 ;
        RECT 74.750 30.930 74.920 32.930 ;
        RECT 75.260 31.730 75.430 42.720 ;
        RECT 76.330 33.220 78.000 43.690 ;
        RECT 78.340 43.220 78.510 43.720 ;
        RECT 79.980 43.220 80.150 43.720 ;
        RECT 78.725 42.990 79.765 43.160 ;
        RECT 78.340 42.430 78.510 42.930 ;
        RECT 79.980 42.430 80.150 42.930 ;
        RECT 78.725 42.200 79.765 42.370 ;
        RECT 78.340 41.640 78.510 42.140 ;
        RECT 79.980 41.640 80.150 42.140 ;
        RECT 78.725 41.410 79.765 41.580 ;
        RECT 78.340 40.850 78.510 41.350 ;
        RECT 79.980 40.850 80.150 41.350 ;
        RECT 78.725 40.620 79.765 40.790 ;
        RECT 78.340 40.060 78.510 40.560 ;
        RECT 79.980 40.060 80.150 40.560 ;
        RECT 78.725 39.830 79.765 40.000 ;
        RECT 78.340 39.270 78.510 39.770 ;
        RECT 79.980 39.270 80.150 39.770 ;
        RECT 78.725 39.040 79.765 39.210 ;
        RECT 78.340 38.480 78.510 38.980 ;
        RECT 79.980 38.480 80.150 38.980 ;
        RECT 78.725 38.250 79.765 38.420 ;
        RECT 78.340 37.690 78.510 38.190 ;
        RECT 79.980 37.690 80.150 38.190 ;
        RECT 78.725 37.460 79.765 37.630 ;
        RECT 78.340 36.900 78.510 37.400 ;
        RECT 79.980 36.900 80.150 37.400 ;
        RECT 78.725 36.670 79.765 36.840 ;
        RECT 78.340 36.110 78.510 36.610 ;
        RECT 79.980 36.110 80.150 36.610 ;
        RECT 78.725 35.880 79.765 36.050 ;
        RECT 78.340 35.320 78.510 35.820 ;
        RECT 79.980 35.320 80.150 35.820 ;
        RECT 78.725 35.090 79.765 35.260 ;
        RECT 78.340 34.530 78.510 35.030 ;
        RECT 79.980 34.530 80.150 35.030 ;
        RECT 78.725 34.300 79.765 34.470 ;
        RECT 78.340 33.740 78.510 34.240 ;
        RECT 79.980 33.740 80.150 34.240 ;
        RECT 78.725 33.510 79.765 33.680 ;
        RECT 80.490 33.220 84.840 49.880 ;
        RECT 94.380 49.800 99.650 49.870 ;
        RECT 101.120 49.800 106.490 49.810 ;
        RECT 94.380 49.630 106.490 49.800 ;
        RECT 94.380 41.710 99.750 49.630 ;
        RECT 100.230 46.990 100.580 49.150 ;
        RECT 100.230 42.190 100.580 44.350 ;
        RECT 101.060 41.710 106.490 49.630 ;
        RECT 94.380 39.790 106.490 41.710 ;
        RECT 94.380 37.390 95.140 39.790 ;
        RECT 95.770 39.280 97.770 39.450 ;
        RECT 98.060 39.280 100.060 39.450 ;
        RECT 100.350 39.280 102.350 39.450 ;
        RECT 102.640 39.280 104.640 39.450 ;
        RECT 95.540 38.070 95.710 39.110 ;
        RECT 97.830 38.070 98.000 39.110 ;
        RECT 100.120 38.070 100.290 39.110 ;
        RECT 102.410 38.070 102.580 39.110 ;
        RECT 104.700 38.070 104.870 39.110 ;
        RECT 95.770 37.730 97.770 37.900 ;
        RECT 98.060 37.730 100.060 37.900 ;
        RECT 100.350 37.730 102.350 37.900 ;
        RECT 102.640 37.730 104.640 37.900 ;
        RECT 105.270 37.390 106.490 39.790 ;
        RECT 94.380 36.810 106.490 37.390 ;
        RECT 94.360 35.380 106.490 36.810 ;
        RECT 94.340 34.100 106.490 35.380 ;
        RECT 117.070 49.490 147.070 52.030 ;
        RECT 117.070 34.780 123.460 49.490 ;
        RECT 124.185 48.920 125.225 49.090 ;
        RECT 123.800 46.860 123.970 48.860 ;
        RECT 125.440 46.860 125.610 48.860 ;
        RECT 124.185 46.630 125.225 46.800 ;
        RECT 123.800 44.570 123.970 46.570 ;
        RECT 125.440 44.570 125.610 46.570 ;
        RECT 124.185 44.340 125.225 44.510 ;
        RECT 123.800 42.280 123.970 44.280 ;
        RECT 125.440 42.280 125.610 44.280 ;
        RECT 124.185 42.050 125.225 42.220 ;
        RECT 123.800 39.990 123.970 41.990 ;
        RECT 125.440 39.990 125.610 41.990 ;
        RECT 124.185 39.760 125.225 39.930 ;
        RECT 123.800 37.700 123.970 39.700 ;
        RECT 125.440 37.700 125.610 39.700 ;
        RECT 124.185 37.470 125.225 37.640 ;
        RECT 123.800 35.410 123.970 37.410 ;
        RECT 125.440 35.410 125.610 37.410 ;
        RECT 124.185 35.180 125.225 35.350 ;
        RECT 125.950 34.780 126.120 49.490 ;
        RECT 128.610 49.480 147.070 49.490 ;
        RECT 126.845 48.920 127.885 49.090 ;
        RECT 126.460 46.860 126.630 48.860 ;
        RECT 128.100 46.860 128.270 48.860 ;
        RECT 126.845 46.630 127.885 46.800 ;
        RECT 126.460 44.570 126.630 46.570 ;
        RECT 128.100 44.570 128.270 46.570 ;
        RECT 126.845 44.340 127.885 44.510 ;
        RECT 126.460 42.280 126.630 44.280 ;
        RECT 128.100 42.280 128.270 44.280 ;
        RECT 128.610 43.290 140.230 49.480 ;
        RECT 140.955 48.910 141.995 49.080 ;
        RECT 140.570 48.350 140.740 48.850 ;
        RECT 142.210 48.350 142.380 48.850 ;
        RECT 140.955 48.120 141.995 48.290 ;
        RECT 140.570 47.560 140.740 48.060 ;
        RECT 142.210 47.560 142.380 48.060 ;
        RECT 140.955 47.330 141.995 47.500 ;
        RECT 140.570 46.770 140.740 47.270 ;
        RECT 142.210 46.770 142.380 47.270 ;
        RECT 140.955 46.540 141.995 46.710 ;
        RECT 140.570 45.980 140.740 46.480 ;
        RECT 142.210 45.980 142.380 46.480 ;
        RECT 140.955 45.750 141.995 45.920 ;
        RECT 140.570 45.190 140.740 45.690 ;
        RECT 142.210 45.190 142.380 45.690 ;
        RECT 140.955 44.960 141.995 45.130 ;
        RECT 140.570 44.400 140.740 44.900 ;
        RECT 142.210 44.400 142.380 44.900 ;
        RECT 140.955 44.170 141.995 44.340 ;
        RECT 140.570 43.610 140.740 44.110 ;
        RECT 142.210 43.610 142.380 44.110 ;
        RECT 140.955 43.380 141.995 43.550 ;
        RECT 126.845 42.050 127.885 42.220 ;
        RECT 126.460 39.990 126.630 41.990 ;
        RECT 128.100 39.990 128.270 41.990 ;
        RECT 126.845 39.760 127.885 39.930 ;
        RECT 126.460 37.700 126.630 39.700 ;
        RECT 128.100 37.700 128.270 39.700 ;
        RECT 126.845 37.470 127.885 37.640 ;
        RECT 126.460 35.410 126.630 37.410 ;
        RECT 128.100 35.410 128.270 37.410 ;
        RECT 126.845 35.180 127.885 35.350 ;
        RECT 128.610 34.780 134.040 43.290 ;
        RECT 117.070 34.410 134.040 34.780 ;
        RECT 134.920 42.320 137.660 42.490 ;
        RECT 117.070 34.400 133.890 34.410 ;
        RECT 134.920 33.880 135.090 42.320 ;
        RECT 135.770 41.750 136.810 41.920 ;
        RECT 135.430 39.690 135.600 41.690 ;
        RECT 136.980 39.690 137.150 41.690 ;
        RECT 135.770 39.460 136.810 39.630 ;
        RECT 135.430 37.400 135.600 39.400 ;
        RECT 136.980 37.400 137.150 39.400 ;
        RECT 135.770 37.170 136.810 37.340 ;
        RECT 135.430 35.110 135.600 37.110 ;
        RECT 136.980 35.110 137.150 37.110 ;
        RECT 135.770 34.880 136.810 35.050 ;
        RECT 76.330 32.690 84.840 33.220 ;
        RECT 117.070 33.710 135.090 33.880 ;
        RECT 73.540 30.700 74.580 30.870 ;
        RECT 54.840 27.170 72.860 30.210 ;
        RECT 73.200 28.640 73.370 30.640 ;
        RECT 74.750 28.640 74.920 30.640 ;
        RECT 73.540 28.410 74.580 28.580 ;
        RECT 54.840 24.770 55.200 27.170 ;
        RECT 55.830 26.660 57.830 26.830 ;
        RECT 58.120 26.660 60.120 26.830 ;
        RECT 60.410 26.660 62.410 26.830 ;
        RECT 62.700 26.660 64.700 26.830 ;
        RECT 55.600 25.450 55.770 26.490 ;
        RECT 57.890 25.450 58.060 26.490 ;
        RECT 60.180 25.450 60.350 26.490 ;
        RECT 62.470 25.450 62.640 26.490 ;
        RECT 64.760 25.450 64.930 26.490 ;
        RECT 65.330 25.720 72.860 27.170 ;
        RECT 73.200 26.350 73.370 28.350 ;
        RECT 74.750 26.350 74.920 28.350 ;
        RECT 73.540 26.120 74.580 26.290 ;
        RECT 75.260 25.720 84.840 31.730 ;
        RECT 55.830 25.110 57.830 25.280 ;
        RECT 58.120 25.110 60.120 25.280 ;
        RECT 60.410 25.110 62.410 25.280 ;
        RECT 62.700 25.110 64.700 25.280 ;
        RECT 65.330 24.770 84.840 25.720 ;
        RECT 54.840 22.450 84.840 24.770 ;
        RECT 117.070 29.810 124.170 33.710 ;
        RECT 124.800 33.200 125.300 33.370 ;
        RECT 124.570 30.490 124.740 33.030 ;
        RECT 125.360 30.490 125.530 33.030 ;
        RECT 124.800 30.150 125.300 30.320 ;
        RECT 125.930 29.810 126.100 33.710 ;
        RECT 126.730 33.200 127.230 33.370 ;
        RECT 126.500 30.490 126.670 33.030 ;
        RECT 127.290 30.490 127.460 33.030 ;
        RECT 126.730 30.150 127.230 30.320 ;
        RECT 127.860 29.810 135.090 33.710 ;
        RECT 135.430 32.820 135.600 34.820 ;
        RECT 136.980 32.820 137.150 34.820 ;
        RECT 135.770 32.590 136.810 32.760 ;
        RECT 135.430 30.530 135.600 32.530 ;
        RECT 136.980 30.530 137.150 32.530 ;
        RECT 137.490 31.330 137.660 42.320 ;
        RECT 138.560 32.820 140.230 43.290 ;
        RECT 140.570 42.820 140.740 43.320 ;
        RECT 142.210 42.820 142.380 43.320 ;
        RECT 140.955 42.590 141.995 42.760 ;
        RECT 140.570 42.030 140.740 42.530 ;
        RECT 142.210 42.030 142.380 42.530 ;
        RECT 140.955 41.800 141.995 41.970 ;
        RECT 140.570 41.240 140.740 41.740 ;
        RECT 142.210 41.240 142.380 41.740 ;
        RECT 140.955 41.010 141.995 41.180 ;
        RECT 140.570 40.450 140.740 40.950 ;
        RECT 142.210 40.450 142.380 40.950 ;
        RECT 140.955 40.220 141.995 40.390 ;
        RECT 140.570 39.660 140.740 40.160 ;
        RECT 142.210 39.660 142.380 40.160 ;
        RECT 140.955 39.430 141.995 39.600 ;
        RECT 140.570 38.870 140.740 39.370 ;
        RECT 142.210 38.870 142.380 39.370 ;
        RECT 140.955 38.640 141.995 38.810 ;
        RECT 140.570 38.080 140.740 38.580 ;
        RECT 142.210 38.080 142.380 38.580 ;
        RECT 140.955 37.850 141.995 38.020 ;
        RECT 140.570 37.290 140.740 37.790 ;
        RECT 142.210 37.290 142.380 37.790 ;
        RECT 140.955 37.060 141.995 37.230 ;
        RECT 140.570 36.500 140.740 37.000 ;
        RECT 142.210 36.500 142.380 37.000 ;
        RECT 140.955 36.270 141.995 36.440 ;
        RECT 140.570 35.710 140.740 36.210 ;
        RECT 142.210 35.710 142.380 36.210 ;
        RECT 140.955 35.480 141.995 35.650 ;
        RECT 140.570 34.920 140.740 35.420 ;
        RECT 142.210 34.920 142.380 35.420 ;
        RECT 140.955 34.690 141.995 34.860 ;
        RECT 140.570 34.130 140.740 34.630 ;
        RECT 142.210 34.130 142.380 34.630 ;
        RECT 140.955 33.900 141.995 34.070 ;
        RECT 140.570 33.340 140.740 33.840 ;
        RECT 142.210 33.340 142.380 33.840 ;
        RECT 140.955 33.110 141.995 33.280 ;
        RECT 142.720 32.820 147.070 49.480 ;
        RECT 138.560 32.290 147.070 32.820 ;
        RECT 135.770 30.300 136.810 30.470 ;
        RECT 117.070 26.770 135.090 29.810 ;
        RECT 135.430 28.240 135.600 30.240 ;
        RECT 136.980 28.240 137.150 30.240 ;
        RECT 135.770 28.010 136.810 28.180 ;
        RECT 117.070 24.370 117.430 26.770 ;
        RECT 118.060 26.260 120.060 26.430 ;
        RECT 120.350 26.260 122.350 26.430 ;
        RECT 122.640 26.260 124.640 26.430 ;
        RECT 124.930 26.260 126.930 26.430 ;
        RECT 117.830 25.050 118.000 26.090 ;
        RECT 120.120 25.050 120.290 26.090 ;
        RECT 122.410 25.050 122.580 26.090 ;
        RECT 124.700 25.050 124.870 26.090 ;
        RECT 126.990 25.050 127.160 26.090 ;
        RECT 127.560 25.320 135.090 26.770 ;
        RECT 135.430 25.950 135.600 27.950 ;
        RECT 136.980 25.950 137.150 27.950 ;
        RECT 135.770 25.720 136.810 25.890 ;
        RECT 137.490 25.320 147.070 31.330 ;
        RECT 118.060 24.710 120.060 24.880 ;
        RECT 120.350 24.710 122.350 24.880 ;
        RECT 122.640 24.710 124.640 24.880 ;
        RECT 124.930 24.710 126.930 24.880 ;
        RECT 127.560 24.370 147.070 25.320 ;
        RECT 54.840 22.430 84.290 22.450 ;
        RECT 117.070 22.050 147.070 24.370 ;
        RECT 117.070 22.030 146.520 22.050 ;
      LAYER mcon ;
        RECT 56.100 51.140 84.500 52.080 ;
        RECT 55.040 50.560 84.500 51.140 ;
        RECT 55.040 46.070 60.510 50.560 ;
        RECT 62.035 49.320 62.915 49.490 ;
        RECT 61.570 47.340 61.740 49.180 ;
        RECT 63.210 47.340 63.380 49.180 ;
        RECT 62.035 47.030 62.915 47.200 ;
        RECT 61.570 45.050 61.740 46.890 ;
        RECT 63.210 45.050 63.380 46.890 ;
        RECT 62.035 44.740 62.915 44.910 ;
        RECT 61.570 42.760 61.740 44.600 ;
        RECT 63.210 42.760 63.380 44.600 ;
        RECT 62.035 42.450 62.915 42.620 ;
        RECT 61.570 40.470 61.740 42.310 ;
        RECT 63.210 40.470 63.380 42.310 ;
        RECT 62.035 40.160 62.915 40.330 ;
        RECT 61.570 38.180 61.740 40.020 ;
        RECT 63.210 38.180 63.380 40.020 ;
        RECT 62.035 37.870 62.915 38.040 ;
        RECT 61.570 35.890 61.740 37.730 ;
        RECT 63.210 35.890 63.380 37.730 ;
        RECT 62.035 35.580 62.915 35.750 ;
        RECT 64.695 49.320 65.575 49.490 ;
        RECT 64.230 47.340 64.400 49.180 ;
        RECT 65.870 47.340 66.040 49.180 ;
        RECT 67.030 48.190 77.340 50.560 ;
        RECT 96.080 50.740 105.390 51.570 ;
        RECT 118.330 50.740 146.730 51.680 ;
        RECT 78.805 49.310 79.685 49.480 ;
        RECT 78.340 48.830 78.510 49.170 ;
        RECT 79.980 48.830 80.150 49.170 ;
        RECT 78.805 48.520 79.685 48.690 ;
        RECT 64.695 47.030 65.575 47.200 ;
        RECT 64.230 45.050 64.400 46.890 ;
        RECT 65.870 45.050 66.040 46.890 ;
        RECT 64.695 44.740 65.575 44.910 ;
        RECT 64.230 42.760 64.400 44.600 ;
        RECT 65.870 42.760 66.040 44.600 ;
        RECT 78.340 48.040 78.510 48.380 ;
        RECT 79.980 48.040 80.150 48.380 ;
        RECT 78.805 47.730 79.685 47.900 ;
        RECT 78.340 47.250 78.510 47.590 ;
        RECT 79.980 47.250 80.150 47.590 ;
        RECT 78.805 46.940 79.685 47.110 ;
        RECT 78.340 46.460 78.510 46.800 ;
        RECT 79.980 46.460 80.150 46.800 ;
        RECT 78.805 46.150 79.685 46.320 ;
        RECT 78.340 45.670 78.510 46.010 ;
        RECT 79.980 45.670 80.150 46.010 ;
        RECT 78.805 45.360 79.685 45.530 ;
        RECT 78.340 44.880 78.510 45.220 ;
        RECT 79.980 44.880 80.150 45.220 ;
        RECT 78.805 44.570 79.685 44.740 ;
        RECT 78.340 44.090 78.510 44.430 ;
        RECT 79.980 44.090 80.150 44.430 ;
        RECT 78.805 43.780 79.685 43.950 ;
        RECT 64.695 42.450 65.575 42.620 ;
        RECT 64.230 40.470 64.400 42.310 ;
        RECT 65.870 40.470 66.040 42.310 ;
        RECT 64.695 40.160 65.575 40.330 ;
        RECT 64.230 38.180 64.400 40.020 ;
        RECT 65.870 38.180 66.040 40.020 ;
        RECT 64.695 37.870 65.575 38.040 ;
        RECT 64.230 35.890 64.400 37.730 ;
        RECT 65.870 35.890 66.040 37.730 ;
        RECT 64.695 35.580 65.575 35.750 ;
        RECT 73.620 42.150 74.500 42.320 ;
        RECT 73.200 40.170 73.370 42.010 ;
        RECT 74.750 40.170 74.920 42.010 ;
        RECT 73.620 39.860 74.500 40.030 ;
        RECT 73.200 37.880 73.370 39.720 ;
        RECT 74.750 37.880 74.920 39.720 ;
        RECT 73.620 37.570 74.500 37.740 ;
        RECT 73.200 35.590 73.370 37.430 ;
        RECT 74.750 35.590 74.920 37.430 ;
        RECT 73.620 35.280 74.500 35.450 ;
        RECT 62.650 33.600 62.990 33.770 ;
        RECT 62.340 30.970 62.510 33.350 ;
        RECT 63.130 30.970 63.300 33.350 ;
        RECT 62.650 30.550 62.990 30.720 ;
        RECT 64.580 33.600 64.920 33.770 ;
        RECT 64.270 30.970 64.440 33.350 ;
        RECT 65.060 30.970 65.230 33.350 ;
        RECT 64.580 30.550 64.920 30.720 ;
        RECT 73.200 33.300 73.370 35.140 ;
        RECT 74.750 33.300 74.920 35.140 ;
        RECT 73.620 32.990 74.500 33.160 ;
        RECT 73.200 31.010 73.370 32.850 ;
        RECT 74.750 31.010 74.920 32.850 ;
        RECT 78.340 43.300 78.510 43.640 ;
        RECT 79.980 43.300 80.150 43.640 ;
        RECT 78.805 42.990 79.685 43.160 ;
        RECT 78.340 42.510 78.510 42.850 ;
        RECT 79.980 42.510 80.150 42.850 ;
        RECT 78.805 42.200 79.685 42.370 ;
        RECT 78.340 41.720 78.510 42.060 ;
        RECT 79.980 41.720 80.150 42.060 ;
        RECT 78.805 41.410 79.685 41.580 ;
        RECT 78.340 40.930 78.510 41.270 ;
        RECT 79.980 40.930 80.150 41.270 ;
        RECT 78.805 40.620 79.685 40.790 ;
        RECT 78.340 40.140 78.510 40.480 ;
        RECT 79.980 40.140 80.150 40.480 ;
        RECT 78.805 39.830 79.685 40.000 ;
        RECT 78.340 39.350 78.510 39.690 ;
        RECT 79.980 39.350 80.150 39.690 ;
        RECT 78.805 39.040 79.685 39.210 ;
        RECT 78.340 38.560 78.510 38.900 ;
        RECT 79.980 38.560 80.150 38.900 ;
        RECT 78.805 38.250 79.685 38.420 ;
        RECT 78.340 37.770 78.510 38.110 ;
        RECT 79.980 37.770 80.150 38.110 ;
        RECT 78.805 37.460 79.685 37.630 ;
        RECT 78.340 36.980 78.510 37.320 ;
        RECT 79.980 36.980 80.150 37.320 ;
        RECT 78.805 36.670 79.685 36.840 ;
        RECT 78.340 36.190 78.510 36.530 ;
        RECT 79.980 36.190 80.150 36.530 ;
        RECT 78.805 35.880 79.685 36.050 ;
        RECT 78.340 35.400 78.510 35.740 ;
        RECT 79.980 35.400 80.150 35.740 ;
        RECT 78.805 35.090 79.685 35.260 ;
        RECT 78.340 34.610 78.510 34.950 ;
        RECT 79.980 34.610 80.150 34.950 ;
        RECT 78.805 34.300 79.685 34.470 ;
        RECT 78.340 33.820 78.510 34.160 ;
        RECT 79.980 33.820 80.150 34.160 ;
        RECT 78.805 33.510 79.685 33.680 ;
        RECT 100.310 47.075 100.500 49.060 ;
        RECT 100.310 42.280 100.500 44.265 ;
        RECT 95.850 39.280 97.690 39.450 ;
        RECT 98.140 39.280 99.980 39.450 ;
        RECT 100.430 39.280 102.270 39.450 ;
        RECT 102.720 39.280 104.560 39.450 ;
        RECT 95.540 38.150 95.710 39.030 ;
        RECT 97.830 38.150 98.000 39.030 ;
        RECT 100.120 38.150 100.290 39.030 ;
        RECT 102.410 38.150 102.580 39.030 ;
        RECT 104.700 38.150 104.870 39.030 ;
        RECT 95.850 37.730 97.690 37.900 ;
        RECT 98.140 37.730 99.980 37.900 ;
        RECT 100.430 37.730 102.270 37.900 ;
        RECT 102.720 37.730 104.560 37.900 ;
        RECT 95.250 34.630 105.560 36.550 ;
        RECT 117.270 50.160 146.730 50.740 ;
        RECT 117.270 45.670 122.740 50.160 ;
        RECT 124.265 48.920 125.145 49.090 ;
        RECT 123.800 46.940 123.970 48.780 ;
        RECT 125.440 46.940 125.610 48.780 ;
        RECT 124.265 46.630 125.145 46.800 ;
        RECT 123.800 44.650 123.970 46.490 ;
        RECT 125.440 44.650 125.610 46.490 ;
        RECT 124.265 44.340 125.145 44.510 ;
        RECT 123.800 42.360 123.970 44.200 ;
        RECT 125.440 42.360 125.610 44.200 ;
        RECT 124.265 42.050 125.145 42.220 ;
        RECT 123.800 40.070 123.970 41.910 ;
        RECT 125.440 40.070 125.610 41.910 ;
        RECT 124.265 39.760 125.145 39.930 ;
        RECT 123.800 37.780 123.970 39.620 ;
        RECT 125.440 37.780 125.610 39.620 ;
        RECT 124.265 37.470 125.145 37.640 ;
        RECT 123.800 35.490 123.970 37.330 ;
        RECT 125.440 35.490 125.610 37.330 ;
        RECT 124.265 35.180 125.145 35.350 ;
        RECT 126.925 48.920 127.805 49.090 ;
        RECT 126.460 46.940 126.630 48.780 ;
        RECT 128.100 46.940 128.270 48.780 ;
        RECT 129.260 47.790 139.570 50.160 ;
        RECT 141.035 48.910 141.915 49.080 ;
        RECT 140.570 48.430 140.740 48.770 ;
        RECT 142.210 48.430 142.380 48.770 ;
        RECT 141.035 48.120 141.915 48.290 ;
        RECT 126.925 46.630 127.805 46.800 ;
        RECT 126.460 44.650 126.630 46.490 ;
        RECT 128.100 44.650 128.270 46.490 ;
        RECT 126.925 44.340 127.805 44.510 ;
        RECT 126.460 42.360 126.630 44.200 ;
        RECT 128.100 42.360 128.270 44.200 ;
        RECT 140.570 47.640 140.740 47.980 ;
        RECT 142.210 47.640 142.380 47.980 ;
        RECT 141.035 47.330 141.915 47.500 ;
        RECT 140.570 46.850 140.740 47.190 ;
        RECT 142.210 46.850 142.380 47.190 ;
        RECT 141.035 46.540 141.915 46.710 ;
        RECT 140.570 46.060 140.740 46.400 ;
        RECT 142.210 46.060 142.380 46.400 ;
        RECT 141.035 45.750 141.915 45.920 ;
        RECT 140.570 45.270 140.740 45.610 ;
        RECT 142.210 45.270 142.380 45.610 ;
        RECT 141.035 44.960 141.915 45.130 ;
        RECT 140.570 44.480 140.740 44.820 ;
        RECT 142.210 44.480 142.380 44.820 ;
        RECT 141.035 44.170 141.915 44.340 ;
        RECT 140.570 43.690 140.740 44.030 ;
        RECT 142.210 43.690 142.380 44.030 ;
        RECT 141.035 43.380 141.915 43.550 ;
        RECT 126.925 42.050 127.805 42.220 ;
        RECT 126.460 40.070 126.630 41.910 ;
        RECT 128.100 40.070 128.270 41.910 ;
        RECT 126.925 39.760 127.805 39.930 ;
        RECT 126.460 37.780 126.630 39.620 ;
        RECT 128.100 37.780 128.270 39.620 ;
        RECT 126.925 37.470 127.805 37.640 ;
        RECT 126.460 35.490 126.630 37.330 ;
        RECT 128.100 35.490 128.270 37.330 ;
        RECT 126.925 35.180 127.805 35.350 ;
        RECT 135.850 41.750 136.730 41.920 ;
        RECT 135.430 39.770 135.600 41.610 ;
        RECT 136.980 39.770 137.150 41.610 ;
        RECT 135.850 39.460 136.730 39.630 ;
        RECT 135.430 37.480 135.600 39.320 ;
        RECT 136.980 37.480 137.150 39.320 ;
        RECT 135.850 37.170 136.730 37.340 ;
        RECT 135.430 35.190 135.600 37.030 ;
        RECT 136.980 35.190 137.150 37.030 ;
        RECT 135.850 34.880 136.730 35.050 ;
        RECT 73.620 30.700 74.500 30.870 ;
        RECT 73.200 28.720 73.370 30.560 ;
        RECT 74.750 28.720 74.920 30.560 ;
        RECT 73.620 28.410 74.500 28.580 ;
        RECT 55.910 26.660 57.750 26.830 ;
        RECT 58.200 26.660 60.040 26.830 ;
        RECT 60.490 26.660 62.330 26.830 ;
        RECT 62.780 26.660 64.620 26.830 ;
        RECT 55.600 25.530 55.770 26.410 ;
        RECT 57.890 25.530 58.060 26.410 ;
        RECT 60.180 25.530 60.350 26.410 ;
        RECT 62.470 25.530 62.640 26.410 ;
        RECT 64.760 25.530 64.930 26.410 ;
        RECT 73.200 26.430 73.370 28.270 ;
        RECT 74.750 26.430 74.920 28.270 ;
        RECT 73.620 26.120 74.500 26.290 ;
        RECT 55.910 25.110 57.750 25.280 ;
        RECT 58.200 25.110 60.040 25.280 ;
        RECT 60.490 25.110 62.330 25.280 ;
        RECT 62.780 25.110 64.620 25.280 ;
        RECT 70.540 24.250 84.430 25.350 ;
        RECT 56.040 22.730 84.440 24.250 ;
        RECT 124.880 33.200 125.220 33.370 ;
        RECT 124.570 30.570 124.740 32.950 ;
        RECT 125.360 30.570 125.530 32.950 ;
        RECT 124.880 30.150 125.220 30.320 ;
        RECT 126.810 33.200 127.150 33.370 ;
        RECT 126.500 30.570 126.670 32.950 ;
        RECT 127.290 30.570 127.460 32.950 ;
        RECT 126.810 30.150 127.150 30.320 ;
        RECT 135.430 32.900 135.600 34.740 ;
        RECT 136.980 32.900 137.150 34.740 ;
        RECT 135.850 32.590 136.730 32.760 ;
        RECT 135.430 30.610 135.600 32.450 ;
        RECT 136.980 30.610 137.150 32.450 ;
        RECT 140.570 42.900 140.740 43.240 ;
        RECT 142.210 42.900 142.380 43.240 ;
        RECT 141.035 42.590 141.915 42.760 ;
        RECT 140.570 42.110 140.740 42.450 ;
        RECT 142.210 42.110 142.380 42.450 ;
        RECT 141.035 41.800 141.915 41.970 ;
        RECT 140.570 41.320 140.740 41.660 ;
        RECT 142.210 41.320 142.380 41.660 ;
        RECT 141.035 41.010 141.915 41.180 ;
        RECT 140.570 40.530 140.740 40.870 ;
        RECT 142.210 40.530 142.380 40.870 ;
        RECT 141.035 40.220 141.915 40.390 ;
        RECT 140.570 39.740 140.740 40.080 ;
        RECT 142.210 39.740 142.380 40.080 ;
        RECT 141.035 39.430 141.915 39.600 ;
        RECT 140.570 38.950 140.740 39.290 ;
        RECT 142.210 38.950 142.380 39.290 ;
        RECT 141.035 38.640 141.915 38.810 ;
        RECT 140.570 38.160 140.740 38.500 ;
        RECT 142.210 38.160 142.380 38.500 ;
        RECT 141.035 37.850 141.915 38.020 ;
        RECT 140.570 37.370 140.740 37.710 ;
        RECT 142.210 37.370 142.380 37.710 ;
        RECT 141.035 37.060 141.915 37.230 ;
        RECT 140.570 36.580 140.740 36.920 ;
        RECT 142.210 36.580 142.380 36.920 ;
        RECT 141.035 36.270 141.915 36.440 ;
        RECT 140.570 35.790 140.740 36.130 ;
        RECT 142.210 35.790 142.380 36.130 ;
        RECT 141.035 35.480 141.915 35.650 ;
        RECT 140.570 35.000 140.740 35.340 ;
        RECT 142.210 35.000 142.380 35.340 ;
        RECT 141.035 34.690 141.915 34.860 ;
        RECT 140.570 34.210 140.740 34.550 ;
        RECT 142.210 34.210 142.380 34.550 ;
        RECT 141.035 33.900 141.915 34.070 ;
        RECT 140.570 33.420 140.740 33.760 ;
        RECT 142.210 33.420 142.380 33.760 ;
        RECT 141.035 33.110 141.915 33.280 ;
        RECT 135.850 30.300 136.730 30.470 ;
        RECT 135.430 28.320 135.600 30.160 ;
        RECT 136.980 28.320 137.150 30.160 ;
        RECT 135.850 28.010 136.730 28.180 ;
        RECT 118.140 26.260 119.980 26.430 ;
        RECT 120.430 26.260 122.270 26.430 ;
        RECT 122.720 26.260 124.560 26.430 ;
        RECT 125.010 26.260 126.850 26.430 ;
        RECT 117.830 25.130 118.000 26.010 ;
        RECT 120.120 25.130 120.290 26.010 ;
        RECT 122.410 25.130 122.580 26.010 ;
        RECT 124.700 25.130 124.870 26.010 ;
        RECT 126.990 25.130 127.160 26.010 ;
        RECT 135.430 26.030 135.600 27.870 ;
        RECT 136.980 26.030 137.150 27.870 ;
        RECT 135.850 25.720 136.730 25.890 ;
        RECT 118.140 24.710 119.980 24.880 ;
        RECT 120.430 24.710 122.270 24.880 ;
        RECT 122.720 24.710 124.560 24.880 ;
        RECT 125.010 24.710 126.850 24.880 ;
        RECT 132.770 23.850 146.660 24.950 ;
        RECT 118.270 22.330 146.670 23.850 ;
      LAYER met1 ;
        RECT 54.810 56.250 77.300 59.710 ;
        RECT 54.810 52.430 77.350 56.250 ;
        RECT 54.810 50.390 84.840 52.430 ;
        RECT 95.020 51.750 105.690 60.270 ;
        RECT 117.080 52.030 134.980 58.630 ;
        RECT 94.700 50.580 105.900 51.750 ;
        RECT 54.840 50.350 84.840 50.390 ;
        RECT 54.840 50.340 77.780 50.350 ;
        RECT 54.840 37.380 60.790 50.340 ;
        RECT 61.530 49.540 63.410 50.340 ;
        RECT 61.910 49.290 63.030 49.540 ;
        RECT 64.200 49.490 66.080 50.340 ;
        RECT 64.630 49.300 65.640 49.490 ;
        RECT 64.635 49.290 65.635 49.300 ;
        RECT 63.210 49.240 64.390 49.270 ;
        RECT 61.540 49.030 61.770 49.240 ;
        RECT 61.540 49.020 61.780 49.030 ;
        RECT 61.530 48.370 61.780 49.020 ;
        RECT 63.180 48.370 64.430 49.240 ;
        RECT 65.840 48.370 66.070 49.240 ;
        RECT 61.530 48.190 66.070 48.370 ;
        RECT 61.530 48.110 61.780 48.190 ;
        RECT 61.530 47.230 61.770 48.110 ;
        RECT 63.180 47.280 64.430 48.190 ;
        RECT 65.840 47.280 66.070 48.190 ;
        RECT 66.710 47.690 77.780 50.340 ;
        RECT 78.310 49.875 80.180 50.105 ;
        RECT 80.950 49.890 84.840 50.350 ;
        RECT 78.310 48.770 78.540 49.875 ;
        RECT 78.710 49.160 79.800 49.640 ;
        RECT 78.330 48.440 78.520 48.770 ;
        RECT 78.310 47.980 78.540 48.440 ;
        RECT 78.710 48.380 79.800 48.860 ;
        RECT 79.950 48.770 80.180 49.875 ;
        RECT 79.970 48.440 80.160 48.770 ;
        RECT 78.330 47.650 78.520 47.980 ;
        RECT 78.310 47.460 78.540 47.650 ;
        RECT 78.700 47.580 79.790 48.060 ;
        RECT 79.950 47.980 80.180 48.440 ;
        RECT 79.970 47.650 80.160 47.980 ;
        RECT 78.060 47.410 78.540 47.460 ;
        RECT 77.890 47.310 78.540 47.410 ;
        RECT 63.180 47.230 64.390 47.280 ;
        RECT 61.530 47.000 64.390 47.230 ;
        RECT 61.530 46.200 61.770 47.000 ;
        RECT 63.180 46.950 64.390 47.000 ;
        RECT 63.180 46.200 64.430 46.950 ;
        RECT 64.580 46.910 65.690 47.280 ;
        RECT 77.490 47.190 78.540 47.310 ;
        RECT 65.840 46.200 66.070 46.950 ;
        RECT 77.490 46.870 78.520 47.190 ;
        RECT 77.890 46.860 78.520 46.870 ;
        RECT 77.890 46.710 78.540 46.860 ;
        RECT 78.700 46.800 79.790 47.280 ;
        RECT 79.950 47.190 80.180 47.650 ;
        RECT 80.960 47.560 83.000 49.890 ;
        RECT 79.970 46.860 80.160 47.190 ;
        RECT 99.970 47.000 100.980 50.580 ;
        RECT 117.070 49.950 147.070 52.030 ;
        RECT 117.070 49.940 140.010 49.950 ;
        RECT 78.310 46.400 78.540 46.710 ;
        RECT 61.530 46.020 66.070 46.200 ;
        RECT 78.330 46.070 78.520 46.400 ;
        RECT 61.530 45.850 61.780 46.020 ;
        RECT 61.530 44.960 61.770 45.850 ;
        RECT 61.530 44.710 61.780 44.960 ;
        RECT 61.530 43.850 61.770 44.710 ;
        RECT 61.950 44.650 62.990 45.010 ;
        RECT 63.180 44.990 64.430 46.020 ;
        RECT 63.190 44.660 64.390 44.990 ;
        RECT 61.530 43.810 61.780 43.850 ;
        RECT 63.180 43.810 64.430 44.660 ;
        RECT 64.630 44.630 65.640 45.030 ;
        RECT 65.840 44.990 66.070 46.020 ;
        RECT 78.310 45.610 78.540 46.070 ;
        RECT 78.690 46.010 79.780 46.490 ;
        RECT 79.950 46.400 80.180 46.860 ;
        RECT 79.970 46.070 80.160 46.400 ;
        RECT 78.330 45.280 78.520 45.610 ;
        RECT 78.310 44.820 78.540 45.280 ;
        RECT 78.700 45.210 79.790 45.690 ;
        RECT 79.950 45.610 80.180 46.070 ;
        RECT 79.970 45.280 80.160 45.610 ;
        RECT 65.840 43.810 66.070 44.660 ;
        RECT 78.330 44.490 78.520 44.820 ;
        RECT 78.310 44.030 78.540 44.490 ;
        RECT 78.720 44.420 79.810 44.900 ;
        RECT 79.950 44.820 80.180 45.280 ;
        RECT 79.970 44.490 80.160 44.820 ;
        RECT 61.530 43.630 66.070 43.810 ;
        RECT 78.330 43.700 78.520 44.030 ;
        RECT 61.530 43.550 61.780 43.630 ;
        RECT 61.530 42.640 61.770 43.550 ;
        RECT 63.180 42.700 64.430 43.630 ;
        RECT 61.975 42.640 62.975 42.650 ;
        RECT 63.180 42.640 64.390 42.700 ;
        RECT 61.530 42.410 64.390 42.640 ;
        RECT 61.530 41.620 61.770 42.410 ;
        RECT 63.180 42.370 64.390 42.410 ;
        RECT 61.530 41.600 61.780 41.620 ;
        RECT 63.180 41.600 64.430 42.370 ;
        RECT 64.580 42.350 65.690 42.720 ;
        RECT 65.840 42.700 66.070 43.630 ;
        RECT 78.310 43.240 78.540 43.700 ;
        RECT 78.710 43.640 79.800 44.120 ;
        RECT 79.950 44.030 80.180 44.490 ;
        RECT 79.970 43.700 80.160 44.030 ;
        RECT 78.330 42.910 78.520 43.240 ;
        RECT 78.310 42.450 78.540 42.910 ;
        RECT 78.720 42.840 79.810 43.320 ;
        RECT 79.950 43.240 80.180 43.700 ;
        RECT 99.930 43.470 100.870 44.560 ;
        RECT 106.985 43.470 108.715 43.500 ;
        RECT 79.970 42.910 80.160 43.240 ;
        RECT 65.840 41.600 66.070 42.370 ;
        RECT 61.530 41.420 66.070 41.600 ;
        RECT 61.530 41.320 61.780 41.420 ;
        RECT 61.530 40.370 61.770 41.320 ;
        RECT 61.530 40.120 61.780 40.370 ;
        RECT 61.530 39.340 61.770 40.120 ;
        RECT 61.960 40.080 63.000 40.440 ;
        RECT 63.180 40.410 64.430 41.420 ;
        RECT 63.190 40.080 64.390 40.410 ;
        RECT 64.620 40.360 65.630 40.460 ;
        RECT 65.840 40.410 66.070 41.420 ;
        RECT 73.170 41.260 73.400 42.070 ;
        RECT 73.560 42.040 74.570 42.400 ;
        RECT 78.330 42.120 78.520 42.450 ;
        RECT 74.720 41.260 74.950 42.070 ;
        RECT 78.310 41.660 78.540 42.120 ;
        RECT 78.710 42.060 79.800 42.540 ;
        RECT 79.950 42.450 80.180 42.910 ;
        RECT 79.970 42.120 80.160 42.450 ;
        RECT 78.330 41.330 78.520 41.660 ;
        RECT 73.170 40.970 74.950 41.260 ;
        RECT 64.620 40.130 65.635 40.360 ;
        RECT 62.020 40.060 62.930 40.080 ;
        RECT 61.530 39.160 61.780 39.340 ;
        RECT 63.180 39.160 64.430 40.080 ;
        RECT 64.620 40.060 65.630 40.130 ;
        RECT 73.170 40.110 73.400 40.970 ;
        RECT 65.840 39.160 66.070 40.080 ;
        RECT 73.190 39.780 73.360 40.110 ;
        RECT 61.530 38.980 66.070 39.160 ;
        RECT 61.530 38.070 61.770 38.980 ;
        RECT 63.180 38.120 64.430 38.980 ;
        RECT 63.180 38.070 64.390 38.120 ;
        RECT 61.530 37.840 64.390 38.070 ;
        RECT 61.530 36.930 61.770 37.840 ;
        RECT 63.180 37.790 64.390 37.840 ;
        RECT 61.530 36.900 61.780 36.930 ;
        RECT 63.180 36.900 64.430 37.790 ;
        RECT 64.580 37.770 65.690 38.140 ;
        RECT 65.840 38.120 66.070 38.980 ;
        RECT 73.170 38.930 73.400 39.780 ;
        RECT 73.540 39.750 74.580 40.140 ;
        RECT 74.720 40.110 74.950 40.970 ;
        RECT 78.310 40.870 78.540 41.330 ;
        RECT 78.720 41.260 79.810 41.740 ;
        RECT 79.950 41.660 80.180 42.120 ;
        RECT 99.930 41.740 108.715 43.470 ;
        RECT 79.970 41.330 80.160 41.660 ;
        RECT 78.330 40.540 78.520 40.870 ;
        RECT 74.760 39.780 74.900 40.110 ;
        RECT 78.310 40.080 78.540 40.540 ;
        RECT 78.710 40.480 79.800 40.960 ;
        RECT 79.950 40.870 80.180 41.330 ;
        RECT 79.970 40.540 80.160 40.870 ;
        RECT 99.930 40.710 100.870 41.740 ;
        RECT 106.985 41.710 108.715 41.740 ;
        RECT 74.720 38.930 74.950 39.780 ;
        RECT 78.330 39.750 78.520 40.080 ;
        RECT 78.310 39.290 78.540 39.750 ;
        RECT 78.700 39.680 79.790 40.160 ;
        RECT 79.950 40.080 80.180 40.540 ;
        RECT 97.370 40.160 103.120 40.710 ;
        RECT 97.340 40.150 103.120 40.160 ;
        RECT 79.970 39.750 80.160 40.080 ;
        RECT 97.340 39.810 103.160 40.150 ;
        RECT 78.330 38.960 78.520 39.290 ;
        RECT 73.170 38.640 74.950 38.930 ;
        RECT 73.170 37.820 73.400 38.640 ;
        RECT 65.840 36.900 66.070 37.790 ;
        RECT 73.190 37.490 73.360 37.820 ;
        RECT 73.550 37.490 74.560 37.850 ;
        RECT 74.720 37.820 74.950 38.640 ;
        RECT 78.310 38.500 78.540 38.960 ;
        RECT 78.710 38.900 79.800 39.380 ;
        RECT 79.950 39.290 80.180 39.750 ;
        RECT 97.340 39.480 98.600 39.810 ;
        RECT 101.900 39.480 103.160 39.810 ;
        RECT 79.970 38.960 80.160 39.290 ;
        RECT 95.790 39.250 100.040 39.480 ;
        RECT 100.370 39.250 104.620 39.480 ;
        RECT 78.330 38.170 78.520 38.500 ;
        RECT 74.760 37.490 74.900 37.820 ;
        RECT 78.310 37.710 78.540 38.170 ;
        RECT 78.710 38.100 79.800 38.580 ;
        RECT 79.950 38.500 80.180 38.960 ;
        RECT 79.970 38.170 80.160 38.500 ;
        RECT 61.530 36.720 66.070 36.900 ;
        RECT 61.530 36.630 61.780 36.720 ;
        RECT 61.530 35.920 61.770 36.630 ;
        RECT 61.530 35.020 61.780 35.920 ;
        RECT 62.020 35.840 62.930 35.850 ;
        RECT 61.980 35.780 62.990 35.840 ;
        RECT 61.975 35.550 62.990 35.780 ;
        RECT 61.980 35.540 62.990 35.550 ;
        RECT 63.180 35.830 64.430 36.720 ;
        RECT 63.180 35.640 64.390 35.830 ;
        RECT 64.640 35.780 65.640 35.840 ;
        RECT 65.840 35.830 66.070 36.720 ;
        RECT 73.170 36.660 73.400 37.490 ;
        RECT 74.720 36.660 74.950 37.490 ;
        RECT 78.330 37.380 78.520 37.710 ;
        RECT 78.310 36.920 78.540 37.380 ;
        RECT 78.710 37.310 79.800 37.790 ;
        RECT 79.950 37.710 80.180 38.170 ;
        RECT 95.060 38.110 96.160 39.110 ;
        RECT 95.510 38.090 95.740 38.110 ;
        RECT 96.620 37.930 99.110 39.250 ;
        RECT 100.090 39.070 100.320 39.090 ;
        RECT 99.640 38.070 100.740 39.070 ;
        RECT 101.220 37.930 103.740 39.250 ;
        RECT 104.190 38.090 105.290 39.090 ;
        RECT 95.790 37.780 100.040 37.930 ;
        RECT 79.970 37.380 80.160 37.710 ;
        RECT 95.790 37.700 97.750 37.780 ;
        RECT 98.080 37.700 100.040 37.780 ;
        RECT 100.370 37.820 104.620 37.930 ;
        RECT 100.370 37.700 102.330 37.820 ;
        RECT 102.660 37.700 104.620 37.820 ;
        RECT 73.170 36.370 74.950 36.660 ;
        RECT 78.330 36.590 78.520 36.920 ;
        RECT 62.020 35.500 62.930 35.540 ;
        RECT 63.180 35.020 63.430 35.640 ;
        RECT 64.635 35.550 65.640 35.780 ;
        RECT 64.640 35.490 65.640 35.550 ;
        RECT 73.170 35.530 73.400 36.370 ;
        RECT 64.670 35.470 65.600 35.490 ;
        RECT 73.190 35.210 73.350 35.530 ;
        RECT 73.190 35.200 73.390 35.210 ;
        RECT 61.530 34.680 63.700 35.020 ;
        RECT 64.710 34.690 65.840 35.110 ;
        RECT 62.570 33.570 63.070 33.860 ;
        RECT 61.940 30.910 62.540 33.420 ;
        RECT 62.680 30.750 62.960 33.570 ;
        RECT 63.310 33.420 63.700 34.680 ;
        RECT 64.500 33.550 65.010 33.850 ;
        RECT 63.100 30.910 63.700 33.420 ;
        RECT 63.870 33.030 64.470 33.410 ;
        RECT 63.840 31.040 64.470 33.030 ;
        RECT 63.870 30.910 64.470 31.040 ;
        RECT 64.610 30.750 64.890 33.550 ;
        RECT 65.250 33.410 65.630 34.690 ;
        RECT 73.170 34.340 73.400 35.200 ;
        RECT 73.540 35.110 74.580 35.620 ;
        RECT 74.720 35.530 74.950 36.370 ;
        RECT 78.310 36.130 78.540 36.590 ;
        RECT 78.720 36.520 79.810 37.000 ;
        RECT 79.950 36.920 80.180 37.380 ;
        RECT 79.970 36.590 80.160 36.920 ;
        RECT 78.330 35.800 78.520 36.130 ;
        RECT 74.760 35.200 74.900 35.530 ;
        RECT 78.310 35.340 78.540 35.800 ;
        RECT 78.710 35.730 79.800 36.210 ;
        RECT 79.950 36.130 80.180 36.590 ;
        RECT 79.970 35.800 80.160 36.130 ;
        RECT 74.720 34.340 74.950 35.200 ;
        RECT 78.330 35.010 78.520 35.340 ;
        RECT 78.310 34.550 78.540 35.010 ;
        RECT 78.720 34.950 79.810 35.430 ;
        RECT 79.950 35.340 80.180 35.800 ;
        RECT 94.870 35.440 106.020 37.020 ;
        RECT 117.070 36.980 123.020 49.940 ;
        RECT 123.760 49.140 125.640 49.940 ;
        RECT 124.140 48.890 125.260 49.140 ;
        RECT 126.430 49.090 128.310 49.940 ;
        RECT 126.860 48.900 127.870 49.090 ;
        RECT 126.865 48.890 127.865 48.900 ;
        RECT 125.440 48.840 126.620 48.870 ;
        RECT 123.770 48.630 124.000 48.840 ;
        RECT 123.770 48.620 124.010 48.630 ;
        RECT 123.760 47.970 124.010 48.620 ;
        RECT 125.410 47.970 126.660 48.840 ;
        RECT 128.070 47.970 128.300 48.840 ;
        RECT 123.760 47.790 128.300 47.970 ;
        RECT 123.760 47.710 124.010 47.790 ;
        RECT 123.760 46.830 124.000 47.710 ;
        RECT 125.410 46.880 126.660 47.790 ;
        RECT 128.070 46.880 128.300 47.790 ;
        RECT 128.940 47.290 140.010 49.940 ;
        RECT 140.540 49.475 142.410 49.705 ;
        RECT 143.180 49.490 147.070 49.950 ;
        RECT 140.540 48.370 140.770 49.475 ;
        RECT 140.940 48.760 142.030 49.240 ;
        RECT 140.560 48.040 140.750 48.370 ;
        RECT 140.540 47.580 140.770 48.040 ;
        RECT 140.940 47.980 142.030 48.460 ;
        RECT 142.180 48.370 142.410 49.475 ;
        RECT 142.200 48.040 142.390 48.370 ;
        RECT 140.560 47.250 140.750 47.580 ;
        RECT 140.540 47.060 140.770 47.250 ;
        RECT 140.930 47.180 142.020 47.660 ;
        RECT 142.180 47.580 142.410 48.040 ;
        RECT 142.200 47.250 142.390 47.580 ;
        RECT 140.290 47.010 140.770 47.060 ;
        RECT 140.120 46.910 140.770 47.010 ;
        RECT 125.410 46.830 126.620 46.880 ;
        RECT 123.760 46.600 126.620 46.830 ;
        RECT 123.760 45.800 124.000 46.600 ;
        RECT 125.410 46.550 126.620 46.600 ;
        RECT 125.410 45.800 126.660 46.550 ;
        RECT 126.810 46.510 127.920 46.880 ;
        RECT 139.720 46.790 140.770 46.910 ;
        RECT 128.070 45.800 128.300 46.550 ;
        RECT 139.720 46.470 140.750 46.790 ;
        RECT 140.120 46.460 140.750 46.470 ;
        RECT 140.120 46.310 140.770 46.460 ;
        RECT 140.930 46.400 142.020 46.880 ;
        RECT 142.180 46.790 142.410 47.250 ;
        RECT 143.190 47.160 145.230 49.490 ;
        RECT 142.200 46.460 142.390 46.790 ;
        RECT 140.540 46.000 140.770 46.310 ;
        RECT 123.760 45.620 128.300 45.800 ;
        RECT 140.560 45.670 140.750 46.000 ;
        RECT 123.760 45.450 124.010 45.620 ;
        RECT 123.760 44.560 124.000 45.450 ;
        RECT 123.760 44.310 124.010 44.560 ;
        RECT 123.760 43.450 124.000 44.310 ;
        RECT 124.180 44.250 125.220 44.610 ;
        RECT 125.410 44.590 126.660 45.620 ;
        RECT 125.420 44.260 126.620 44.590 ;
        RECT 123.760 43.410 124.010 43.450 ;
        RECT 125.410 43.410 126.660 44.260 ;
        RECT 126.860 44.230 127.870 44.630 ;
        RECT 128.070 44.590 128.300 45.620 ;
        RECT 140.540 45.210 140.770 45.670 ;
        RECT 140.920 45.610 142.010 46.090 ;
        RECT 142.180 46.000 142.410 46.460 ;
        RECT 142.200 45.670 142.390 46.000 ;
        RECT 140.560 44.880 140.750 45.210 ;
        RECT 140.540 44.420 140.770 44.880 ;
        RECT 140.930 44.810 142.020 45.290 ;
        RECT 142.180 45.210 142.410 45.670 ;
        RECT 142.200 44.880 142.390 45.210 ;
        RECT 128.070 43.410 128.300 44.260 ;
        RECT 140.560 44.090 140.750 44.420 ;
        RECT 140.540 43.630 140.770 44.090 ;
        RECT 140.950 44.020 142.040 44.500 ;
        RECT 142.180 44.420 142.410 44.880 ;
        RECT 142.200 44.090 142.390 44.420 ;
        RECT 123.760 43.230 128.300 43.410 ;
        RECT 140.560 43.300 140.750 43.630 ;
        RECT 123.760 43.150 124.010 43.230 ;
        RECT 123.760 42.240 124.000 43.150 ;
        RECT 125.410 42.300 126.660 43.230 ;
        RECT 124.205 42.240 125.205 42.250 ;
        RECT 125.410 42.240 126.620 42.300 ;
        RECT 123.760 42.010 126.620 42.240 ;
        RECT 123.760 41.220 124.000 42.010 ;
        RECT 125.410 41.970 126.620 42.010 ;
        RECT 123.760 41.200 124.010 41.220 ;
        RECT 125.410 41.200 126.660 41.970 ;
        RECT 126.810 41.950 127.920 42.320 ;
        RECT 128.070 42.300 128.300 43.230 ;
        RECT 140.540 42.840 140.770 43.300 ;
        RECT 140.940 43.240 142.030 43.720 ;
        RECT 142.180 43.630 142.410 44.090 ;
        RECT 142.200 43.300 142.390 43.630 ;
        RECT 140.560 42.510 140.750 42.840 ;
        RECT 140.540 42.050 140.770 42.510 ;
        RECT 140.950 42.440 142.040 42.920 ;
        RECT 142.180 42.840 142.410 43.300 ;
        RECT 142.200 42.510 142.390 42.840 ;
        RECT 128.070 41.200 128.300 41.970 ;
        RECT 123.760 41.020 128.300 41.200 ;
        RECT 123.760 40.920 124.010 41.020 ;
        RECT 123.760 39.970 124.000 40.920 ;
        RECT 123.760 39.720 124.010 39.970 ;
        RECT 123.760 38.940 124.000 39.720 ;
        RECT 124.190 39.680 125.230 40.040 ;
        RECT 125.410 40.010 126.660 41.020 ;
        RECT 125.420 39.680 126.620 40.010 ;
        RECT 126.850 39.960 127.860 40.060 ;
        RECT 128.070 40.010 128.300 41.020 ;
        RECT 135.400 40.860 135.630 41.670 ;
        RECT 135.790 41.640 136.800 42.000 ;
        RECT 140.560 41.720 140.750 42.050 ;
        RECT 136.950 40.860 137.180 41.670 ;
        RECT 140.540 41.260 140.770 41.720 ;
        RECT 140.940 41.660 142.030 42.140 ;
        RECT 142.180 42.050 142.410 42.510 ;
        RECT 142.200 41.720 142.390 42.050 ;
        RECT 140.560 40.930 140.750 41.260 ;
        RECT 135.400 40.570 137.180 40.860 ;
        RECT 126.850 39.730 127.865 39.960 ;
        RECT 124.250 39.660 125.160 39.680 ;
        RECT 123.760 38.760 124.010 38.940 ;
        RECT 125.410 38.760 126.660 39.680 ;
        RECT 126.850 39.660 127.860 39.730 ;
        RECT 135.400 39.710 135.630 40.570 ;
        RECT 128.070 38.760 128.300 39.680 ;
        RECT 135.420 39.380 135.590 39.710 ;
        RECT 123.760 38.580 128.300 38.760 ;
        RECT 123.760 37.670 124.000 38.580 ;
        RECT 125.410 37.720 126.660 38.580 ;
        RECT 125.410 37.670 126.620 37.720 ;
        RECT 123.760 37.440 126.620 37.670 ;
        RECT 123.760 36.530 124.000 37.440 ;
        RECT 125.410 37.390 126.620 37.440 ;
        RECT 123.760 36.500 124.010 36.530 ;
        RECT 125.410 36.500 126.660 37.390 ;
        RECT 126.810 37.370 127.920 37.740 ;
        RECT 128.070 37.720 128.300 38.580 ;
        RECT 135.400 38.530 135.630 39.380 ;
        RECT 135.770 39.350 136.810 39.740 ;
        RECT 136.950 39.710 137.180 40.570 ;
        RECT 140.540 40.470 140.770 40.930 ;
        RECT 140.950 40.860 142.040 41.340 ;
        RECT 142.180 41.260 142.410 41.720 ;
        RECT 142.200 40.930 142.390 41.260 ;
        RECT 140.560 40.140 140.750 40.470 ;
        RECT 136.990 39.380 137.130 39.710 ;
        RECT 140.540 39.680 140.770 40.140 ;
        RECT 140.940 40.080 142.030 40.560 ;
        RECT 142.180 40.470 142.410 40.930 ;
        RECT 142.200 40.140 142.390 40.470 ;
        RECT 136.950 38.530 137.180 39.380 ;
        RECT 140.560 39.350 140.750 39.680 ;
        RECT 140.540 38.890 140.770 39.350 ;
        RECT 140.930 39.280 142.020 39.760 ;
        RECT 142.180 39.680 142.410 40.140 ;
        RECT 142.200 39.350 142.390 39.680 ;
        RECT 140.560 38.560 140.750 38.890 ;
        RECT 135.400 38.240 137.180 38.530 ;
        RECT 135.400 37.420 135.630 38.240 ;
        RECT 128.070 36.500 128.300 37.390 ;
        RECT 135.420 37.090 135.590 37.420 ;
        RECT 135.780 37.090 136.790 37.450 ;
        RECT 136.950 37.420 137.180 38.240 ;
        RECT 140.540 38.100 140.770 38.560 ;
        RECT 140.940 38.500 142.030 38.980 ;
        RECT 142.180 38.890 142.410 39.350 ;
        RECT 142.200 38.560 142.390 38.890 ;
        RECT 140.560 37.770 140.750 38.100 ;
        RECT 136.990 37.090 137.130 37.420 ;
        RECT 140.540 37.310 140.770 37.770 ;
        RECT 140.940 37.700 142.030 38.180 ;
        RECT 142.180 38.100 142.410 38.560 ;
        RECT 142.200 37.770 142.390 38.100 ;
        RECT 123.760 36.320 128.300 36.500 ;
        RECT 123.760 36.230 124.010 36.320 ;
        RECT 123.760 35.520 124.000 36.230 ;
        RECT 79.970 35.010 80.160 35.340 ;
        RECT 73.170 34.155 74.950 34.340 ;
        RECT 78.330 34.220 78.520 34.550 ;
        RECT 65.030 30.900 65.630 33.410 ;
        RECT 68.025 34.050 74.950 34.155 ;
        RECT 68.025 33.240 73.400 34.050 ;
        RECT 74.720 33.240 74.950 34.050 ;
        RECT 78.310 33.760 78.540 34.220 ;
        RECT 78.710 34.140 79.800 34.620 ;
        RECT 79.950 34.550 80.180 35.010 ;
        RECT 79.970 34.220 80.160 34.550 ;
        RECT 79.950 33.760 80.180 34.220 ;
        RECT 78.330 33.720 78.520 33.760 ;
        RECT 78.710 33.320 79.770 33.760 ;
        RECT 79.970 33.750 80.160 33.760 ;
        RECT 68.025 33.180 73.360 33.240 ;
        RECT 54.870 28.585 56.020 30.450 ;
        RECT 62.570 29.370 63.070 30.750 ;
        RECT 64.500 30.140 65.000 30.750 ;
        RECT 66.615 30.140 67.210 30.260 ;
        RECT 64.500 29.730 67.210 30.140 ;
        RECT 66.615 29.605 67.210 29.730 ;
        RECT 62.570 28.790 64.810 29.370 ;
        RECT 68.025 28.585 69.000 33.180 ;
        RECT 73.190 32.910 73.360 33.180 ;
        RECT 73.540 32.950 74.580 33.210 ;
        RECT 74.760 32.910 74.900 33.240 ;
        RECT 73.170 32.100 73.400 32.910 ;
        RECT 74.720 32.100 74.950 32.910 ;
        RECT 73.170 31.810 74.950 32.100 ;
        RECT 73.170 30.950 73.400 31.810 ;
        RECT 73.190 30.620 73.360 30.950 ;
        RECT 73.170 29.760 73.400 30.620 ;
        RECT 73.540 30.580 74.580 30.970 ;
        RECT 74.720 30.950 74.950 31.810 ;
        RECT 74.760 30.620 74.900 30.950 ;
        RECT 74.720 29.760 74.950 30.620 ;
        RECT 73.170 29.470 74.950 29.760 ;
        RECT 73.170 28.660 73.400 29.470 ;
        RECT 74.720 28.660 74.950 29.470 ;
        RECT 54.870 27.730 69.000 28.585 ;
        RECT 73.190 28.330 73.360 28.660 ;
        RECT 73.540 28.360 74.580 28.630 ;
        RECT 74.760 28.330 74.900 28.660 ;
        RECT 54.880 27.725 69.000 27.730 ;
        RECT 54.880 27.720 68.570 27.725 ;
        RECT 56.260 27.030 57.010 27.720 ;
        RECT 73.170 27.490 73.400 28.330 ;
        RECT 74.720 27.490 74.950 28.330 ;
        RECT 73.170 27.200 74.950 27.490 ;
        RECT 56.260 26.860 63.990 27.030 ;
        RECT 55.850 26.660 64.680 26.860 ;
        RECT 55.850 26.630 57.810 26.660 ;
        RECT 58.140 26.630 60.100 26.660 ;
        RECT 60.430 26.630 62.390 26.660 ;
        RECT 62.720 26.630 64.680 26.660 ;
        RECT 55.490 25.470 55.850 26.470 ;
        RECT 56.630 25.310 57.010 26.630 ;
        RECT 57.790 25.470 58.170 26.470 ;
        RECT 58.940 25.310 59.320 26.630 ;
        RECT 60.070 25.470 60.450 26.470 ;
        RECT 61.180 25.310 61.560 26.630 ;
        RECT 62.360 25.470 62.740 26.470 ;
        RECT 63.520 25.310 63.900 26.630 ;
        RECT 64.660 25.470 65.040 26.470 ;
        RECT 73.170 26.370 73.400 27.200 ;
        RECT 73.540 26.060 74.580 26.400 ;
        RECT 74.720 26.370 74.950 27.200 ;
        RECT 74.760 26.330 74.900 26.370 ;
        RECT 73.560 25.660 74.560 26.060 ;
        RECT 55.850 25.080 57.810 25.310 ;
        RECT 58.140 25.080 60.100 25.310 ;
        RECT 60.430 25.080 62.390 25.310 ;
        RECT 62.720 25.080 64.680 25.310 ;
        RECT 65.530 24.480 84.840 25.660 ;
        RECT 54.840 10.670 84.840 24.480 ;
        RECT 94.300 10.990 106.280 35.440 ;
        RECT 123.760 34.620 124.010 35.520 ;
        RECT 124.250 35.440 125.160 35.450 ;
        RECT 124.210 35.380 125.220 35.440 ;
        RECT 124.205 35.150 125.220 35.380 ;
        RECT 124.210 35.140 125.220 35.150 ;
        RECT 125.410 35.430 126.660 36.320 ;
        RECT 125.410 35.240 126.620 35.430 ;
        RECT 126.870 35.380 127.870 35.440 ;
        RECT 128.070 35.430 128.300 36.320 ;
        RECT 135.400 36.260 135.630 37.090 ;
        RECT 136.950 36.260 137.180 37.090 ;
        RECT 140.560 36.980 140.750 37.310 ;
        RECT 140.540 36.520 140.770 36.980 ;
        RECT 140.940 36.910 142.030 37.390 ;
        RECT 142.180 37.310 142.410 37.770 ;
        RECT 142.200 36.980 142.390 37.310 ;
        RECT 135.400 35.970 137.180 36.260 ;
        RECT 140.560 36.190 140.750 36.520 ;
        RECT 124.250 35.100 125.160 35.140 ;
        RECT 125.410 34.620 125.660 35.240 ;
        RECT 126.865 35.150 127.870 35.380 ;
        RECT 126.870 35.090 127.870 35.150 ;
        RECT 135.400 35.130 135.630 35.970 ;
        RECT 126.900 35.070 127.830 35.090 ;
        RECT 135.420 34.810 135.580 35.130 ;
        RECT 135.420 34.800 135.620 34.810 ;
        RECT 123.760 34.280 125.930 34.620 ;
        RECT 126.940 34.290 128.070 34.710 ;
        RECT 124.800 33.170 125.300 33.460 ;
        RECT 124.170 30.510 124.770 33.020 ;
        RECT 124.910 30.350 125.190 33.170 ;
        RECT 125.540 33.020 125.930 34.280 ;
        RECT 126.730 33.150 127.240 33.450 ;
        RECT 125.330 30.510 125.930 33.020 ;
        RECT 126.100 32.630 126.700 33.010 ;
        RECT 126.070 30.640 126.700 32.630 ;
        RECT 126.100 30.510 126.700 30.640 ;
        RECT 126.840 30.350 127.120 33.150 ;
        RECT 127.480 33.010 127.860 34.290 ;
        RECT 135.400 33.940 135.630 34.800 ;
        RECT 135.770 34.710 136.810 35.220 ;
        RECT 136.950 35.130 137.180 35.970 ;
        RECT 140.540 35.730 140.770 36.190 ;
        RECT 140.950 36.120 142.040 36.600 ;
        RECT 142.180 36.520 142.410 36.980 ;
        RECT 142.200 36.190 142.390 36.520 ;
        RECT 140.560 35.400 140.750 35.730 ;
        RECT 136.990 34.800 137.130 35.130 ;
        RECT 140.540 34.940 140.770 35.400 ;
        RECT 140.940 35.330 142.030 35.810 ;
        RECT 142.180 35.730 142.410 36.190 ;
        RECT 142.200 35.400 142.390 35.730 ;
        RECT 136.950 33.940 137.180 34.800 ;
        RECT 140.560 34.610 140.750 34.940 ;
        RECT 140.540 34.150 140.770 34.610 ;
        RECT 140.950 34.550 142.040 35.030 ;
        RECT 142.180 34.940 142.410 35.400 ;
        RECT 142.200 34.610 142.390 34.940 ;
        RECT 135.400 33.755 137.180 33.940 ;
        RECT 140.560 33.820 140.750 34.150 ;
        RECT 127.260 30.500 127.860 33.010 ;
        RECT 130.255 33.650 137.180 33.755 ;
        RECT 130.255 32.840 135.630 33.650 ;
        RECT 136.950 32.840 137.180 33.650 ;
        RECT 140.540 33.360 140.770 33.820 ;
        RECT 140.940 33.740 142.030 34.220 ;
        RECT 142.180 34.150 142.410 34.610 ;
        RECT 142.200 33.820 142.390 34.150 ;
        RECT 142.180 33.360 142.410 33.820 ;
        RECT 140.560 33.320 140.750 33.360 ;
        RECT 140.940 32.920 142.000 33.360 ;
        RECT 142.200 33.350 142.390 33.360 ;
        RECT 130.255 32.780 135.590 32.840 ;
        RECT 117.100 28.185 118.250 30.050 ;
        RECT 124.800 28.970 125.300 30.350 ;
        RECT 126.730 29.740 127.230 30.350 ;
        RECT 128.845 29.740 129.440 29.860 ;
        RECT 126.730 29.330 129.440 29.740 ;
        RECT 128.845 29.205 129.440 29.330 ;
        RECT 124.800 28.390 127.040 28.970 ;
        RECT 130.255 28.185 131.230 32.780 ;
        RECT 135.420 32.510 135.590 32.780 ;
        RECT 135.770 32.550 136.810 32.810 ;
        RECT 136.990 32.510 137.130 32.840 ;
        RECT 135.400 31.700 135.630 32.510 ;
        RECT 136.950 31.700 137.180 32.510 ;
        RECT 135.400 31.410 137.180 31.700 ;
        RECT 135.400 30.550 135.630 31.410 ;
        RECT 135.420 30.220 135.590 30.550 ;
        RECT 135.400 29.360 135.630 30.220 ;
        RECT 135.770 30.180 136.810 30.570 ;
        RECT 136.950 30.550 137.180 31.410 ;
        RECT 136.990 30.220 137.130 30.550 ;
        RECT 136.950 29.360 137.180 30.220 ;
        RECT 135.400 29.070 137.180 29.360 ;
        RECT 135.400 28.260 135.630 29.070 ;
        RECT 136.950 28.260 137.180 29.070 ;
        RECT 117.100 27.330 131.230 28.185 ;
        RECT 135.420 27.930 135.590 28.260 ;
        RECT 135.770 27.960 136.810 28.230 ;
        RECT 136.990 27.930 137.130 28.260 ;
        RECT 117.110 27.325 131.230 27.330 ;
        RECT 117.110 27.320 130.800 27.325 ;
        RECT 118.490 26.630 119.240 27.320 ;
        RECT 135.400 27.090 135.630 27.930 ;
        RECT 136.950 27.090 137.180 27.930 ;
        RECT 135.400 26.800 137.180 27.090 ;
        RECT 118.490 26.460 126.220 26.630 ;
        RECT 118.080 26.260 126.910 26.460 ;
        RECT 118.080 26.230 120.040 26.260 ;
        RECT 120.370 26.230 122.330 26.260 ;
        RECT 122.660 26.230 124.620 26.260 ;
        RECT 124.950 26.230 126.910 26.260 ;
        RECT 117.720 25.070 118.080 26.070 ;
        RECT 118.860 24.910 119.240 26.230 ;
        RECT 120.020 25.070 120.400 26.070 ;
        RECT 121.170 24.910 121.550 26.230 ;
        RECT 122.300 25.070 122.680 26.070 ;
        RECT 123.410 24.910 123.790 26.230 ;
        RECT 124.590 25.070 124.970 26.070 ;
        RECT 125.750 24.910 126.130 26.230 ;
        RECT 126.890 25.070 127.270 26.070 ;
        RECT 135.400 25.970 135.630 26.800 ;
        RECT 135.770 25.660 136.810 26.000 ;
        RECT 136.950 25.970 137.180 26.800 ;
        RECT 136.990 25.930 137.130 25.970 ;
        RECT 135.790 25.260 136.790 25.660 ;
        RECT 118.080 24.680 120.040 24.910 ;
        RECT 120.370 24.680 122.330 24.910 ;
        RECT 122.660 24.680 124.620 24.910 ;
        RECT 124.950 24.680 126.910 24.910 ;
        RECT 127.760 24.080 147.070 25.260 ;
        RECT 117.070 23.460 147.070 24.080 ;
        RECT 117.070 22.030 147.050 23.460 ;
        RECT 117.100 12.950 146.870 22.030 ;
        RECT 117.100 12.940 127.920 12.950 ;
      LAYER via ;
        RECT 55.340 55.020 76.610 59.300 ;
        RECT 95.400 55.090 105.220 59.770 ;
        RECT 62.000 49.290 62.940 49.650 ;
        RECT 64.680 49.300 65.590 49.700 ;
        RECT 78.760 49.160 79.750 49.640 ;
        RECT 78.760 48.380 79.750 48.860 ;
        RECT 78.750 47.580 79.740 48.060 ;
        RECT 64.630 46.910 65.640 47.280 ;
        RECT 77.540 46.870 78.230 47.310 ;
        RECT 78.750 46.800 79.740 47.280 ;
        RECT 81.010 47.560 82.950 51.910 ;
        RECT 117.310 54.830 134.530 58.370 ;
        RECT 62.000 44.650 62.940 45.010 ;
        RECT 64.680 44.630 65.590 45.030 ;
        RECT 78.740 46.010 79.730 46.490 ;
        RECT 78.750 45.210 79.740 45.690 ;
        RECT 78.770 44.420 79.760 44.900 ;
        RECT 64.630 42.350 65.640 42.720 ;
        RECT 78.760 43.640 79.750 44.120 ;
        RECT 78.770 42.840 79.760 43.320 ;
        RECT 62.010 40.080 62.950 40.440 ;
        RECT 64.670 40.060 65.580 40.460 ;
        RECT 73.610 42.040 74.520 42.400 ;
        RECT 78.760 42.060 79.750 42.540 ;
        RECT 78.770 41.260 79.760 41.740 ;
        RECT 106.985 41.740 108.715 43.470 ;
        RECT 73.590 39.820 74.540 40.100 ;
        RECT 64.630 37.770 65.640 38.140 ;
        RECT 78.760 40.480 79.750 40.960 ;
        RECT 78.750 39.680 79.740 40.160 ;
        RECT 73.600 37.490 74.510 37.850 ;
        RECT 78.760 38.900 79.750 39.380 ;
        RECT 78.760 38.100 79.750 38.580 ;
        RECT 62.030 35.540 62.940 35.840 ;
        RECT 64.690 35.490 65.590 35.840 ;
        RECT 78.760 37.310 79.750 37.790 ;
        RECT 95.110 38.110 96.110 39.110 ;
        RECT 97.400 38.090 98.400 39.090 ;
        RECT 99.690 38.070 100.690 39.070 ;
        RECT 101.950 38.090 102.950 39.090 ;
        RECT 104.240 38.090 105.240 39.090 ;
        RECT 64.760 34.690 65.790 35.110 ;
        RECT 61.960 31.020 62.410 33.080 ;
        RECT 63.890 31.040 64.310 33.030 ;
        RECT 73.580 35.110 74.540 35.620 ;
        RECT 78.770 36.520 79.760 37.000 ;
        RECT 78.760 35.730 79.750 36.210 ;
        RECT 124.230 48.890 125.170 49.250 ;
        RECT 126.910 48.900 127.820 49.300 ;
        RECT 140.990 48.760 141.980 49.240 ;
        RECT 140.990 47.980 141.980 48.460 ;
        RECT 140.980 47.180 141.970 47.660 ;
        RECT 126.860 46.510 127.870 46.880 ;
        RECT 139.770 46.470 140.460 46.910 ;
        RECT 140.980 46.400 141.970 46.880 ;
        RECT 143.240 47.160 145.180 51.510 ;
        RECT 124.230 44.250 125.170 44.610 ;
        RECT 126.910 44.230 127.820 44.630 ;
        RECT 140.970 45.610 141.960 46.090 ;
        RECT 140.980 44.810 141.970 45.290 ;
        RECT 141.000 44.020 141.990 44.500 ;
        RECT 126.860 41.950 127.870 42.320 ;
        RECT 140.990 43.240 141.980 43.720 ;
        RECT 141.000 42.440 141.990 42.920 ;
        RECT 124.240 39.680 125.180 40.040 ;
        RECT 126.900 39.660 127.810 40.060 ;
        RECT 135.840 41.640 136.750 42.000 ;
        RECT 140.990 41.660 141.980 42.140 ;
        RECT 141.000 40.860 141.990 41.340 ;
        RECT 135.820 39.420 136.770 39.700 ;
        RECT 95.580 36.400 104.840 36.500 ;
        RECT 78.770 34.950 79.760 35.430 ;
        RECT 95.500 35.670 104.860 36.400 ;
        RECT 126.860 37.370 127.870 37.740 ;
        RECT 140.990 40.080 141.980 40.560 ;
        RECT 140.980 39.280 141.970 39.760 ;
        RECT 135.830 37.090 136.740 37.450 ;
        RECT 140.990 38.500 141.980 38.980 ;
        RECT 140.990 37.700 141.980 38.180 ;
        RECT 78.760 34.140 79.750 34.620 ;
        RECT 78.760 33.320 79.720 33.760 ;
        RECT 54.960 28.560 55.960 30.370 ;
        RECT 66.615 29.635 67.210 30.230 ;
        RECT 64.290 28.820 64.810 29.340 ;
        RECT 73.570 32.950 74.550 33.210 ;
        RECT 73.580 30.620 74.540 30.940 ;
        RECT 73.570 28.360 74.540 28.630 ;
        RECT 55.540 25.470 55.800 26.470 ;
        RECT 57.840 25.470 58.120 26.470 ;
        RECT 60.120 25.470 60.400 26.470 ;
        RECT 62.410 25.470 62.690 26.470 ;
        RECT 64.710 25.470 64.990 26.470 ;
        RECT 73.590 26.100 74.540 26.360 ;
        RECT 55.560 23.840 64.950 24.420 ;
        RECT 55.390 11.400 64.190 18.240 ;
        RECT 74.330 11.280 83.680 18.120 ;
        RECT 124.260 35.140 125.170 35.440 ;
        RECT 126.920 35.090 127.820 35.440 ;
        RECT 140.990 36.910 141.980 37.390 ;
        RECT 126.990 34.290 128.020 34.710 ;
        RECT 124.190 30.620 124.640 32.680 ;
        RECT 126.120 30.640 126.540 32.630 ;
        RECT 135.810 34.710 136.770 35.220 ;
        RECT 141.000 36.120 141.990 36.600 ;
        RECT 140.990 35.330 141.980 35.810 ;
        RECT 141.000 34.550 141.990 35.030 ;
        RECT 140.990 33.740 141.980 34.220 ;
        RECT 140.990 32.920 141.950 33.360 ;
        RECT 117.190 28.160 118.190 29.970 ;
        RECT 128.845 29.235 129.440 29.830 ;
        RECT 126.520 28.420 127.040 28.940 ;
        RECT 135.800 32.550 136.780 32.810 ;
        RECT 135.810 30.220 136.770 30.540 ;
        RECT 135.800 27.960 136.770 28.230 ;
        RECT 117.770 25.070 118.030 26.070 ;
        RECT 120.070 25.070 120.350 26.070 ;
        RECT 122.350 25.070 122.630 26.070 ;
        RECT 124.640 25.070 124.920 26.070 ;
        RECT 126.940 25.070 127.220 26.070 ;
        RECT 135.820 25.700 136.770 25.960 ;
        RECT 117.790 23.440 127.180 24.020 ;
        RECT 94.640 11.670 105.730 18.200 ;
        RECT 117.320 13.120 127.600 18.610 ;
        RECT 135.980 13.520 146.160 18.400 ;
      LAYER met2 ;
        RECT 54.930 54.700 77.070 59.620 ;
        RECT 62.000 49.240 62.940 49.700 ;
        RECT 64.680 49.250 65.590 49.750 ;
        RECT 78.760 49.110 79.750 49.690 ;
        RECT 81.010 48.920 82.950 51.960 ;
        RECT 95.020 50.660 105.690 60.270 ;
        RECT 117.160 54.670 134.820 58.500 ;
        RECT 78.760 48.340 82.950 48.920 ;
        RECT 124.230 48.840 125.170 49.300 ;
        RECT 126.910 48.850 127.820 49.350 ;
        RECT 140.990 48.710 141.980 49.290 ;
        RECT 143.240 48.520 145.180 51.560 ;
        RECT 78.760 48.330 79.750 48.340 ;
        RECT 78.750 47.530 79.740 48.110 ;
        RECT 81.010 47.510 82.950 48.340 ;
        RECT 140.990 47.940 145.180 48.520 ;
        RECT 140.990 47.930 141.980 47.940 ;
        RECT 64.630 47.305 65.640 47.330 ;
        RECT 77.540 47.305 78.230 47.360 ;
        RECT 81.030 47.330 82.050 47.510 ;
        RECT 64.630 46.875 78.505 47.305 ;
        RECT 64.630 46.860 65.640 46.875 ;
        RECT 62.000 44.600 62.940 45.060 ;
        RECT 64.680 44.580 65.590 45.080 ;
        RECT 64.630 42.735 65.640 42.770 ;
        RECT 66.425 42.735 66.855 46.875 ;
        RECT 77.540 46.820 78.230 46.875 ;
        RECT 78.750 46.750 82.050 47.330 ;
        RECT 140.980 47.130 141.970 47.710 ;
        RECT 143.240 47.110 145.180 47.940 ;
        RECT 78.740 45.960 79.730 46.540 ;
        RECT 81.030 45.740 82.050 46.750 ;
        RECT 126.860 46.905 127.870 46.930 ;
        RECT 139.770 46.905 140.460 46.960 ;
        RECT 143.260 46.930 144.280 47.110 ;
        RECT 126.860 46.475 140.735 46.905 ;
        RECT 126.860 46.460 127.870 46.475 ;
        RECT 78.750 45.160 82.050 45.740 ;
        RECT 78.770 44.370 79.760 44.950 ;
        RECT 81.030 44.170 82.050 45.160 ;
        RECT 124.230 44.200 125.170 44.660 ;
        RECT 126.910 44.180 127.820 44.680 ;
        RECT 78.760 43.590 82.050 44.170 ;
        RECT 78.770 42.790 79.760 43.370 ;
        RECT 64.630 42.305 66.855 42.735 ;
        RECT 81.030 42.590 82.050 43.590 ;
        RECT 75.030 42.570 75.890 42.580 ;
        RECT 73.620 42.450 75.890 42.570 ;
        RECT 64.630 42.300 65.640 42.305 ;
        RECT 62.010 40.030 62.950 40.490 ;
        RECT 64.670 40.010 65.580 40.510 ;
        RECT 64.630 38.145 65.640 38.190 ;
        RECT 66.425 38.145 66.855 42.305 ;
        RECT 73.610 41.990 75.890 42.450 ;
        RECT 78.760 42.030 82.050 42.590 ;
        RECT 78.760 42.010 79.750 42.030 ;
        RECT 73.620 41.840 75.890 41.990 ;
        RECT 73.590 39.770 74.540 40.150 ;
        RECT 64.615 37.715 66.855 38.145 ;
        RECT 75.030 38.020 75.890 41.840 ;
        RECT 78.770 41.210 79.760 41.790 ;
        RECT 78.760 40.995 79.750 41.010 ;
        RECT 81.030 40.995 82.050 42.030 ;
        RECT 106.955 41.740 108.745 43.470 ;
        RECT 126.860 42.335 127.870 42.370 ;
        RECT 128.655 42.335 129.085 46.475 ;
        RECT 139.770 46.420 140.460 46.475 ;
        RECT 140.980 46.350 144.280 46.930 ;
        RECT 140.970 45.560 141.960 46.140 ;
        RECT 143.260 45.340 144.280 46.350 ;
        RECT 140.980 44.760 144.280 45.340 ;
        RECT 141.000 43.970 141.990 44.550 ;
        RECT 143.260 43.770 144.280 44.760 ;
        RECT 140.990 43.190 144.280 43.770 ;
        RECT 141.000 42.390 141.990 42.970 ;
        RECT 126.860 41.905 129.085 42.335 ;
        RECT 143.260 42.190 144.280 43.190 ;
        RECT 137.260 42.170 138.120 42.180 ;
        RECT 135.850 42.050 138.120 42.170 ;
        RECT 126.860 41.900 127.870 41.905 ;
        RECT 78.760 40.435 82.050 40.995 ;
        RECT 78.760 40.430 79.750 40.435 ;
        RECT 78.750 39.630 79.740 40.210 ;
        RECT 78.760 39.425 79.750 39.430 ;
        RECT 81.030 39.425 82.050 40.435 ;
        RECT 78.760 38.870 82.050 39.425 ;
        RECT 78.760 38.850 79.750 38.870 ;
        RECT 78.760 38.050 79.750 38.630 ;
        RECT 62.030 35.490 62.940 35.890 ;
        RECT 64.690 35.440 65.590 35.890 ;
        RECT 64.760 35.110 65.790 35.160 ;
        RECT 66.425 35.110 66.855 37.715 ;
        RECT 73.600 37.290 75.890 38.020 ;
        RECT 64.750 34.680 66.855 35.110 ;
        RECT 73.580 35.060 74.540 35.670 ;
        RECT 64.760 34.640 65.790 34.680 ;
        RECT 75.030 33.490 75.890 37.290 ;
        RECT 78.760 37.825 79.750 37.840 ;
        RECT 81.030 37.825 82.050 38.870 ;
        RECT 95.110 38.060 96.110 39.160 ;
        RECT 78.760 37.270 82.050 37.825 ;
        RECT 78.760 37.260 79.750 37.270 ;
        RECT 78.770 36.470 79.760 37.050 ;
        RECT 81.030 36.260 82.050 37.270 ;
        RECT 95.360 36.700 95.900 38.060 ;
        RECT 97.400 38.040 98.400 39.140 ;
        RECT 99.690 38.020 100.690 39.120 ;
        RECT 101.950 38.040 102.950 39.140 ;
        RECT 104.240 38.040 105.240 39.140 ;
        RECT 99.920 36.700 100.460 38.020 ;
        RECT 104.470 36.700 105.010 38.040 ;
        RECT 78.760 35.680 82.050 36.260 ;
        RECT 78.770 34.900 79.760 35.480 ;
        RECT 81.030 34.670 82.050 35.680 ;
        RECT 95.330 35.460 105.150 36.700 ;
        RECT 78.760 34.110 82.050 34.670 ;
        RECT 78.760 34.090 81.690 34.110 ;
        RECT 78.760 33.810 79.700 33.850 ;
        RECT 78.760 33.770 79.720 33.810 ;
        RECT 59.530 30.960 64.390 33.110 ;
        RECT 73.530 32.760 75.890 33.490 ;
        RECT 78.730 33.250 79.750 33.770 ;
        RECT 75.030 31.850 75.890 32.760 ;
        RECT 78.750 31.850 79.750 33.250 ;
        RECT 75.030 31.550 84.770 31.850 ;
        RECT 54.960 30.310 55.960 30.420 ;
        RECT 51.990 29.440 55.960 30.310 ;
        RECT 51.990 21.815 52.860 29.440 ;
        RECT 54.960 28.510 55.960 29.440 ;
        RECT 59.530 28.760 60.875 30.960 ;
        RECT 63.420 30.950 64.390 30.960 ;
        RECT 73.580 30.520 74.540 31.040 ;
        RECT 75.030 30.950 90.920 31.550 ;
        RECT 75.030 30.590 84.770 30.950 ;
        RECT 66.585 30.215 67.240 30.230 ;
        RECT 66.585 29.645 69.925 30.215 ;
        RECT 66.585 29.635 67.240 29.645 ;
        RECT 64.260 29.300 65.290 29.340 ;
        RECT 66.200 29.300 67.280 29.340 ;
        RECT 64.260 28.820 67.280 29.300 ;
        RECT 59.530 28.590 60.870 28.760 ;
        RECT 57.840 27.790 62.690 28.590 ;
        RECT 66.760 27.870 67.280 28.820 ;
        RECT 69.355 28.090 69.925 29.645 ;
        RECT 75.030 28.850 75.890 30.590 ;
        RECT 73.560 28.120 75.890 28.850 ;
        RECT 55.540 25.000 55.800 26.520 ;
        RECT 57.840 25.420 58.120 27.790 ;
        RECT 60.120 25.420 60.400 26.520 ;
        RECT 62.410 25.420 62.690 27.790 ;
        RECT 64.710 25.420 64.990 26.520 ;
        RECT 60.130 25.000 60.390 25.420 ;
        RECT 64.720 25.000 64.980 25.420 ;
        RECT 55.540 23.840 64.980 25.000 ;
        RECT 55.560 23.790 64.950 23.840 ;
        RECT 66.520 22.580 67.520 27.870 ;
        RECT 69.140 23.520 70.140 28.090 ;
        RECT 73.590 26.000 74.540 26.440 ;
        RECT 90.320 23.705 90.920 30.950 ;
        RECT 106.985 29.840 108.715 41.740 ;
        RECT 124.240 39.630 125.180 40.090 ;
        RECT 126.900 39.610 127.810 40.110 ;
        RECT 126.860 37.745 127.870 37.790 ;
        RECT 128.655 37.745 129.085 41.905 ;
        RECT 135.840 41.590 138.120 42.050 ;
        RECT 140.990 41.630 144.280 42.190 ;
        RECT 140.990 41.610 141.980 41.630 ;
        RECT 135.850 41.440 138.120 41.590 ;
        RECT 135.820 39.370 136.770 39.750 ;
        RECT 126.845 37.315 129.085 37.745 ;
        RECT 137.260 37.620 138.120 41.440 ;
        RECT 141.000 40.810 141.990 41.390 ;
        RECT 140.990 40.595 141.980 40.610 ;
        RECT 143.260 40.595 144.280 41.630 ;
        RECT 140.990 40.035 144.280 40.595 ;
        RECT 140.990 40.030 141.980 40.035 ;
        RECT 140.980 39.230 141.970 39.810 ;
        RECT 140.990 39.025 141.980 39.030 ;
        RECT 143.260 39.025 144.280 40.035 ;
        RECT 140.990 38.470 144.280 39.025 ;
        RECT 140.990 38.450 141.980 38.470 ;
        RECT 140.990 37.650 141.980 38.230 ;
        RECT 124.260 35.090 125.170 35.490 ;
        RECT 126.920 35.040 127.820 35.490 ;
        RECT 126.990 34.710 128.020 34.760 ;
        RECT 128.655 34.710 129.085 37.315 ;
        RECT 135.830 36.890 138.120 37.620 ;
        RECT 126.980 34.280 129.085 34.710 ;
        RECT 135.810 34.660 136.770 35.270 ;
        RECT 126.990 34.240 128.020 34.280 ;
        RECT 137.260 33.090 138.120 36.890 ;
        RECT 140.990 37.425 141.980 37.440 ;
        RECT 143.260 37.425 144.280 38.470 ;
        RECT 140.990 36.870 144.280 37.425 ;
        RECT 140.990 36.860 141.980 36.870 ;
        RECT 141.000 36.070 141.990 36.650 ;
        RECT 143.260 35.860 144.280 36.870 ;
        RECT 140.990 35.280 144.280 35.860 ;
        RECT 141.000 34.500 141.990 35.080 ;
        RECT 143.260 34.270 144.280 35.280 ;
        RECT 140.990 33.710 144.280 34.270 ;
        RECT 140.990 33.690 143.920 33.710 ;
        RECT 140.990 33.410 141.930 33.450 ;
        RECT 140.990 33.370 141.950 33.410 ;
        RECT 121.760 30.560 126.620 32.710 ;
        RECT 135.760 32.360 138.120 33.090 ;
        RECT 140.960 32.850 141.980 33.370 ;
        RECT 137.260 31.450 138.120 32.360 ;
        RECT 140.980 31.450 141.980 32.850 ;
        RECT 137.260 31.150 147.000 31.450 ;
        RECT 106.985 29.830 113.910 29.840 ;
        RECT 117.190 29.830 118.190 30.020 ;
        RECT 106.985 29.070 118.190 29.830 ;
        RECT 106.985 29.050 111.750 29.070 ;
        RECT 107.225 26.410 108.095 29.050 ;
        RECT 117.190 28.110 118.190 29.070 ;
        RECT 121.760 28.360 123.105 30.560 ;
        RECT 125.650 30.550 126.620 30.560 ;
        RECT 135.810 30.120 136.770 30.640 ;
        RECT 137.260 30.550 151.130 31.150 ;
        RECT 137.260 30.190 147.000 30.550 ;
        RECT 128.815 29.815 129.470 29.830 ;
        RECT 128.815 29.245 132.155 29.815 ;
        RECT 128.815 29.235 129.470 29.245 ;
        RECT 126.490 28.900 127.520 28.940 ;
        RECT 128.430 28.900 129.510 28.940 ;
        RECT 126.490 28.420 129.510 28.900 ;
        RECT 121.760 28.190 123.100 28.360 ;
        RECT 120.070 27.390 124.920 28.190 ;
        RECT 128.990 27.470 129.510 28.420 ;
        RECT 131.585 27.690 132.155 29.245 ;
        RECT 137.260 28.450 138.120 30.190 ;
        RECT 135.790 27.720 138.120 28.450 ;
        RECT 107.205 25.590 108.115 26.410 ;
        RECT 107.225 25.565 108.095 25.590 ;
        RECT 117.770 24.600 118.030 26.120 ;
        RECT 120.070 25.020 120.350 27.390 ;
        RECT 122.350 25.020 122.630 26.120 ;
        RECT 124.640 25.020 124.920 27.390 ;
        RECT 126.940 25.020 127.220 26.120 ;
        RECT 122.360 24.600 122.620 25.020 ;
        RECT 126.950 24.600 127.210 25.020 ;
        RECT 69.130 23.320 70.140 23.520 ;
        RECT 69.030 22.720 70.140 23.320 ;
        RECT 90.300 23.155 90.940 23.705 ;
        RECT 117.770 23.440 127.210 24.600 ;
        RECT 117.790 23.390 127.180 23.440 ;
        RECT 90.320 23.130 90.920 23.155 ;
        RECT 51.990 20.945 60.930 21.815 ;
        RECT 55.150 10.850 64.860 18.920 ;
        RECT 66.730 9.340 67.330 22.580 ;
        RECT 69.130 22.520 70.140 22.720 ;
        RECT 61.300 8.740 67.330 9.340 ;
        RECT 56.435 5.380 56.985 5.400 ;
        RECT 61.300 5.380 61.900 8.740 ;
        RECT 69.450 7.975 70.050 22.520 ;
        RECT 128.750 22.180 129.750 27.470 ;
        RECT 131.370 23.120 132.370 27.690 ;
        RECT 135.820 25.600 136.770 26.040 ;
        RECT 73.660 10.790 84.410 18.850 ;
        RECT 94.350 11.450 105.980 18.660 ;
        RECT 117.190 13.030 127.820 18.860 ;
        RECT 69.430 7.425 70.070 7.975 ;
        RECT 69.450 7.400 70.050 7.425 ;
        RECT 128.970 7.165 129.570 22.180 ;
        RECT 131.360 22.120 132.370 23.120 ;
        RECT 131.570 20.610 132.170 22.120 ;
        RECT 150.530 20.735 151.130 30.550 ;
        RECT 134.505 20.610 135.055 20.630 ;
        RECT 131.570 20.010 135.080 20.610 ;
        RECT 150.510 20.185 151.150 20.735 ;
        RECT 150.530 20.160 151.130 20.185 ;
        RECT 134.505 19.990 135.055 20.010 ;
        RECT 135.840 13.390 146.360 18.670 ;
        RECT 128.950 6.615 129.590 7.165 ;
        RECT 128.970 6.590 129.570 6.615 ;
        RECT 56.410 4.780 61.900 5.380 ;
        RECT 56.435 4.760 56.985 4.780 ;
      LAYER via2 ;
        RECT 55.340 55.020 76.610 59.300 ;
        RECT 95.400 55.090 105.220 59.770 ;
        RECT 62.000 49.290 62.940 49.650 ;
        RECT 64.680 49.300 65.590 49.700 ;
        RECT 78.760 49.160 79.750 49.640 ;
        RECT 117.310 54.830 134.530 58.370 ;
        RECT 124.230 48.890 125.170 49.250 ;
        RECT 126.910 48.900 127.820 49.300 ;
        RECT 140.990 48.760 141.980 49.240 ;
        RECT 78.750 47.580 79.740 48.060 ;
        RECT 62.000 44.650 62.940 45.010 ;
        RECT 64.680 44.630 65.590 45.030 ;
        RECT 140.980 47.180 141.970 47.660 ;
        RECT 78.740 46.010 79.730 46.490 ;
        RECT 78.770 44.420 79.760 44.900 ;
        RECT 124.230 44.250 125.170 44.610 ;
        RECT 126.910 44.230 127.820 44.630 ;
        RECT 78.770 42.840 79.760 43.320 ;
        RECT 62.010 40.080 62.950 40.440 ;
        RECT 64.670 40.060 65.580 40.460 ;
        RECT 73.590 39.820 74.540 40.100 ;
        RECT 78.770 41.260 79.760 41.740 ;
        RECT 140.970 45.610 141.960 46.090 ;
        RECT 141.000 44.020 141.990 44.500 ;
        RECT 141.000 42.440 141.990 42.920 ;
        RECT 78.750 39.680 79.740 40.160 ;
        RECT 78.760 38.100 79.750 38.580 ;
        RECT 62.030 35.540 62.940 35.840 ;
        RECT 64.690 35.490 65.590 35.840 ;
        RECT 73.580 35.110 74.540 35.620 ;
        RECT 78.770 36.520 79.760 37.000 ;
        RECT 78.770 34.950 79.760 35.430 ;
        RECT 78.760 33.230 79.700 33.800 ;
        RECT 73.580 30.570 74.540 30.990 ;
        RECT 73.590 26.050 74.540 26.390 ;
        RECT 124.240 39.680 125.180 40.040 ;
        RECT 126.900 39.660 127.810 40.060 ;
        RECT 135.820 39.420 136.770 39.700 ;
        RECT 141.000 40.860 141.990 41.340 ;
        RECT 140.980 39.280 141.970 39.760 ;
        RECT 140.990 37.700 141.980 38.180 ;
        RECT 124.260 35.140 125.170 35.440 ;
        RECT 126.920 35.090 127.820 35.440 ;
        RECT 135.810 34.710 136.770 35.220 ;
        RECT 141.000 36.120 141.990 36.600 ;
        RECT 141.000 34.550 141.990 35.030 ;
        RECT 140.990 32.830 141.930 33.400 ;
        RECT 135.810 30.170 136.770 30.590 ;
        RECT 107.250 25.590 108.070 26.410 ;
        RECT 90.345 23.155 90.895 23.705 ;
        RECT 60.015 20.945 60.885 21.815 ;
        RECT 55.390 11.400 64.190 18.240 ;
        RECT 135.820 25.650 136.770 25.990 ;
        RECT 74.330 11.280 83.680 18.120 ;
        RECT 94.640 11.670 105.730 18.200 ;
        RECT 117.320 13.120 127.600 18.610 ;
        RECT 69.475 7.425 70.025 7.975 ;
        RECT 134.505 20.035 135.055 20.585 ;
        RECT 150.555 20.185 151.105 20.735 ;
        RECT 135.980 13.520 146.160 18.400 ;
        RECT 128.995 6.615 129.545 7.165 ;
        RECT 56.435 4.805 56.985 5.355 ;
      LAYER met3 ;
        RECT 54.930 54.700 77.070 59.620 ;
        RECT 95.020 50.660 105.690 60.270 ;
        RECT 117.160 54.670 134.820 58.500 ;
        RECT 62.020 49.675 62.960 49.850 ;
        RECT 64.680 49.725 65.580 50.260 ;
        RECT 61.950 49.265 62.990 49.675 ;
        RECT 64.630 49.275 65.640 49.725 ;
        RECT 78.760 49.665 79.770 49.670 ;
        RECT 62.020 45.035 62.960 49.265 ;
        RECT 64.680 45.055 65.580 49.275 ;
        RECT 78.710 49.135 79.800 49.665 ;
        RECT 124.250 49.275 125.190 49.450 ;
        RECT 126.910 49.325 127.810 49.860 ;
        RECT 78.760 48.085 79.770 49.135 ;
        RECT 124.180 48.865 125.220 49.275 ;
        RECT 126.860 48.875 127.870 49.325 ;
        RECT 140.990 49.265 142.000 49.270 ;
        RECT 78.700 47.555 79.790 48.085 ;
        RECT 78.760 46.515 79.770 47.555 ;
        RECT 78.690 45.985 79.780 46.515 ;
        RECT 61.950 44.625 62.990 45.035 ;
        RECT 62.020 40.465 62.960 44.625 ;
        RECT 64.630 44.605 65.640 45.055 ;
        RECT 78.760 44.925 79.770 45.985 ;
        RECT 64.680 40.485 65.580 44.605 ;
        RECT 78.720 44.395 79.810 44.925 ;
        RECT 124.250 44.635 125.190 48.865 ;
        RECT 126.910 44.655 127.810 48.875 ;
        RECT 140.940 48.735 142.030 49.265 ;
        RECT 140.990 47.685 142.000 48.735 ;
        RECT 140.930 47.155 142.020 47.685 ;
        RECT 140.990 46.115 142.000 47.155 ;
        RECT 140.920 45.585 142.010 46.115 ;
        RECT 78.760 43.345 79.770 44.395 ;
        RECT 124.180 44.225 125.220 44.635 ;
        RECT 78.720 42.815 79.810 43.345 ;
        RECT 78.760 41.765 79.770 42.815 ;
        RECT 78.720 41.235 79.810 41.765 ;
        RECT 61.960 40.055 63.000 40.465 ;
        RECT 62.020 35.865 62.960 40.055 ;
        RECT 64.620 40.035 65.630 40.485 ;
        RECT 64.680 35.865 65.580 40.035 ;
        RECT 61.980 35.515 62.990 35.865 ;
        RECT 64.640 35.465 65.640 35.865 ;
        RECT 64.680 35.440 65.580 35.465 ;
        RECT 73.500 25.770 74.620 40.290 ;
        RECT 78.760 40.185 79.770 41.235 ;
        RECT 78.700 39.655 79.790 40.185 ;
        RECT 124.250 40.065 125.190 44.225 ;
        RECT 126.860 44.205 127.870 44.655 ;
        RECT 140.990 44.525 142.000 45.585 ;
        RECT 126.910 40.085 127.810 44.205 ;
        RECT 140.950 43.995 142.040 44.525 ;
        RECT 140.990 42.945 142.000 43.995 ;
        RECT 140.950 42.415 142.040 42.945 ;
        RECT 140.990 41.365 142.000 42.415 ;
        RECT 140.950 40.835 142.040 41.365 ;
        RECT 124.190 39.655 125.230 40.065 ;
        RECT 78.760 38.605 79.770 39.655 ;
        RECT 78.710 38.075 79.800 38.605 ;
        RECT 78.760 37.025 79.770 38.075 ;
        RECT 78.720 36.495 79.810 37.025 ;
        RECT 78.760 35.455 79.770 36.495 ;
        RECT 124.250 35.465 125.190 39.655 ;
        RECT 126.850 39.635 127.860 40.085 ;
        RECT 126.910 35.465 127.810 39.635 ;
        RECT 78.720 34.925 79.810 35.455 ;
        RECT 124.210 35.115 125.220 35.465 ;
        RECT 126.870 35.065 127.870 35.465 ;
        RECT 126.910 35.040 127.810 35.065 ;
        RECT 78.760 33.825 79.770 34.925 ;
        RECT 78.710 33.320 79.770 33.825 ;
        RECT 78.710 33.205 79.750 33.320 ;
        RECT 87.245 25.565 108.095 26.435 ;
        RECT 59.990 21.815 60.910 21.840 ;
        RECT 87.245 21.815 88.115 25.565 ;
        RECT 135.730 25.370 136.850 39.890 ;
        RECT 140.990 39.785 142.000 40.835 ;
        RECT 140.930 39.255 142.020 39.785 ;
        RECT 140.990 38.205 142.000 39.255 ;
        RECT 140.940 37.675 142.030 38.205 ;
        RECT 140.990 36.625 142.000 37.675 ;
        RECT 140.950 36.095 142.040 36.625 ;
        RECT 140.990 35.055 142.000 36.095 ;
        RECT 140.950 34.525 142.040 35.055 ;
        RECT 140.990 33.425 142.000 34.525 ;
        RECT 140.940 32.920 142.000 33.425 ;
        RECT 140.940 32.805 141.980 32.920 ;
        RECT 59.990 20.945 88.115 21.815 ;
        RECT 59.990 20.920 60.910 20.945 ;
        RECT 55.150 10.850 64.860 18.920 ;
        RECT 73.660 10.790 84.410 18.850 ;
        RECT 68.240 7.400 70.050 8.000 ;
        RECT 46.165 5.380 46.755 5.405 ;
        RECT 46.160 4.780 57.010 5.380 ;
        RECT 46.165 4.755 46.755 4.780 ;
        RECT 68.240 2.835 68.840 7.400 ;
        RECT 90.320 2.925 90.920 23.730 ;
        RECT 94.350 11.450 105.980 18.660 ;
        RECT 117.190 13.030 127.820 18.860 ;
        RECT 112.400 6.590 129.570 7.190 ;
        RECT 112.400 3.135 113.000 6.590 ;
        RECT 134.480 3.365 135.080 20.610 ;
        RECT 135.840 13.390 146.360 18.670 ;
        RECT 150.530 4.705 151.130 20.760 ;
        RECT 150.505 4.115 151.155 4.705 ;
        RECT 150.530 4.110 151.130 4.115 ;
        RECT 68.215 2.245 68.865 2.835 ;
        RECT 90.295 2.335 90.945 2.925 ;
        RECT 112.375 2.545 113.025 3.135 ;
        RECT 134.455 2.775 135.105 3.365 ;
        RECT 150.530 3.065 151.130 3.100 ;
        RECT 134.480 2.770 135.080 2.775 ;
        RECT 112.400 2.540 113.000 2.545 ;
        RECT 150.505 2.475 151.155 3.065 ;
        RECT 150.530 2.440 151.130 2.475 ;
        RECT 90.320 2.330 90.920 2.335 ;
        RECT 68.240 2.240 68.840 2.245 ;
      LAYER via3 ;
        RECT 55.340 55.020 76.610 59.300 ;
        RECT 95.400 55.090 105.220 59.770 ;
        RECT 117.310 54.830 134.530 58.370 ;
        RECT 55.390 11.400 64.190 18.240 ;
        RECT 74.330 11.280 83.680 18.120 ;
        RECT 46.165 4.785 46.755 5.375 ;
        RECT 94.640 11.670 105.730 18.200 ;
        RECT 117.320 13.120 127.600 18.610 ;
        RECT 135.980 13.520 146.160 18.400 ;
        RECT 150.535 4.115 151.125 4.705 ;
        RECT 68.245 2.245 68.835 2.835 ;
        RECT 90.325 2.335 90.915 2.925 ;
        RECT 112.405 2.545 112.995 3.135 ;
        RECT 134.485 2.775 135.075 3.365 ;
        RECT 150.530 2.470 151.130 3.070 ;
      LAYER met4 ;
        RECT 3.990 223.170 4.290 224.760 ;
        RECT 7.670 223.170 7.970 224.760 ;
        RECT 11.350 223.170 11.650 224.760 ;
        RECT 15.030 223.170 15.330 224.760 ;
        RECT 18.710 223.170 19.010 224.760 ;
        RECT 22.390 223.170 22.690 224.760 ;
        RECT 26.070 223.170 26.370 224.760 ;
        RECT 29.750 223.170 30.050 224.760 ;
        RECT 33.430 223.170 33.730 224.760 ;
        RECT 37.110 223.170 37.410 224.760 ;
        RECT 40.790 223.170 41.090 224.760 ;
        RECT 44.470 223.170 44.770 224.760 ;
        RECT 48.150 223.170 48.450 224.760 ;
        RECT 51.830 223.170 52.130 224.760 ;
        RECT 55.510 223.170 55.810 224.760 ;
        RECT 59.190 223.170 59.490 224.760 ;
        RECT 62.870 223.170 63.170 224.760 ;
        RECT 66.550 223.170 66.850 224.760 ;
        RECT 70.230 223.170 70.530 224.760 ;
        RECT 73.910 223.170 74.210 224.760 ;
        RECT 77.590 223.170 77.890 224.760 ;
        RECT 81.270 223.170 81.570 224.760 ;
        RECT 84.950 223.170 85.250 224.760 ;
        RECT 88.630 223.170 88.930 224.760 ;
        RECT 3.990 222.870 156.790 223.170 ;
        RECT 18.710 222.860 19.010 222.870 ;
        RECT 156.490 220.680 156.790 222.870 ;
        RECT 2.500 54.710 152.680 63.120 ;
        RECT 2.500 54.590 93.820 54.710 ;
        RECT 107.870 54.590 152.680 54.710 ;
        RECT 99.610 19.000 100.800 19.040 ;
        RECT 51.320 10.470 155.860 19.000 ;
        RECT 46.160 1.000 46.760 5.380 ;
        RECT 68.240 1.000 68.840 2.840 ;
        RECT 90.320 1.000 90.920 2.930 ;
        RECT 112.400 1.000 113.000 3.140 ;
        RECT 134.480 1.000 135.080 3.370 ;
        RECT 150.530 3.075 151.130 4.710 ;
        RECT 150.525 3.070 151.135 3.075 ;
        RECT 150.525 2.470 157.160 3.070 ;
        RECT 150.525 2.465 151.135 2.470 ;
        RECT 156.560 1.000 157.160 2.470 ;
  END
END tt_um_argunda_tiny_opamp
END LIBRARY

