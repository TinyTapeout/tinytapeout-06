module tt_um_MichaelBell_tinyQV (VGND,
    VPWR,
    clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input VGND;
 input VPWR;
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire _2933_;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire _2945_;
 wire _2946_;
 wire _2947_;
 wire _2948_;
 wire _2949_;
 wire _2950_;
 wire _2951_;
 wire _2952_;
 wire _2953_;
 wire _2954_;
 wire _2955_;
 wire _2956_;
 wire _2957_;
 wire _2958_;
 wire _2959_;
 wire _2960_;
 wire _2961_;
 wire _2962_;
 wire _2963_;
 wire _2964_;
 wire _2965_;
 wire _2966_;
 wire _2967_;
 wire _2968_;
 wire _2969_;
 wire _2970_;
 wire _2971_;
 wire _2972_;
 wire _2973_;
 wire _2974_;
 wire _2975_;
 wire _2976_;
 wire _2977_;
 wire _2978_;
 wire _2979_;
 wire _2980_;
 wire _2981_;
 wire _2982_;
 wire _2983_;
 wire _2984_;
 wire _2985_;
 wire _2986_;
 wire _2987_;
 wire _2988_;
 wire _2989_;
 wire _2990_;
 wire _2991_;
 wire _2992_;
 wire _2993_;
 wire _2994_;
 wire _2995_;
 wire _2996_;
 wire _2997_;
 wire _2998_;
 wire _2999_;
 wire _3000_;
 wire _3001_;
 wire _3002_;
 wire _3003_;
 wire _3004_;
 wire _3005_;
 wire _3006_;
 wire _3007_;
 wire _3008_;
 wire _3009_;
 wire _3010_;
 wire _3011_;
 wire _3012_;
 wire _3013_;
 wire _3014_;
 wire _3015_;
 wire _3016_;
 wire _3017_;
 wire _3018_;
 wire _3019_;
 wire _3020_;
 wire _3021_;
 wire _3022_;
 wire _3023_;
 wire _3024_;
 wire _3025_;
 wire _3026_;
 wire _3027_;
 wire _3028_;
 wire _3029_;
 wire _3030_;
 wire _3031_;
 wire _3032_;
 wire _3033_;
 wire _3034_;
 wire _3035_;
 wire _3036_;
 wire _3037_;
 wire _3038_;
 wire _3039_;
 wire _3040_;
 wire _3041_;
 wire _3042_;
 wire _3043_;
 wire _3044_;
 wire _3045_;
 wire _3046_;
 wire _3047_;
 wire _3048_;
 wire _3049_;
 wire _3050_;
 wire _3051_;
 wire _3052_;
 wire _3053_;
 wire _3054_;
 wire _3055_;
 wire _3056_;
 wire _3057_;
 wire _3058_;
 wire _3059_;
 wire _3060_;
 wire _3061_;
 wire _3062_;
 wire _3063_;
 wire _3064_;
 wire _3065_;
 wire _3066_;
 wire _3067_;
 wire _3068_;
 wire _3069_;
 wire _3070_;
 wire _3071_;
 wire _3072_;
 wire _3073_;
 wire _3074_;
 wire _3075_;
 wire _3076_;
 wire _3077_;
 wire _3078_;
 wire _3079_;
 wire _3080_;
 wire _3081_;
 wire _3082_;
 wire _3083_;
 wire _3084_;
 wire _3085_;
 wire _3086_;
 wire _3087_;
 wire _3088_;
 wire _3089_;
 wire _3090_;
 wire _3091_;
 wire _3092_;
 wire _3093_;
 wire _3094_;
 wire _3095_;
 wire _3096_;
 wire _3097_;
 wire _3098_;
 wire _3099_;
 wire _3100_;
 wire _3101_;
 wire _3102_;
 wire _3103_;
 wire _3104_;
 wire _3105_;
 wire _3106_;
 wire _3107_;
 wire _3108_;
 wire _3109_;
 wire _3110_;
 wire _3111_;
 wire _3112_;
 wire _3113_;
 wire _3114_;
 wire _3115_;
 wire _3116_;
 wire _3117_;
 wire _3118_;
 wire _3119_;
 wire _3120_;
 wire _3121_;
 wire _3122_;
 wire _3123_;
 wire _3124_;
 wire _3125_;
 wire _3126_;
 wire _3127_;
 wire _3128_;
 wire _3129_;
 wire _3130_;
 wire _3131_;
 wire _3132_;
 wire _3133_;
 wire _3134_;
 wire _3135_;
 wire _3136_;
 wire _3137_;
 wire _3138_;
 wire _3139_;
 wire _3140_;
 wire _3141_;
 wire _3142_;
 wire _3143_;
 wire _3144_;
 wire _3145_;
 wire _3146_;
 wire _3147_;
 wire _3148_;
 wire _3149_;
 wire _3150_;
 wire _3151_;
 wire _3152_;
 wire _3153_;
 wire _3154_;
 wire _3155_;
 wire _3156_;
 wire _3157_;
 wire _3158_;
 wire _3159_;
 wire _3160_;
 wire _3161_;
 wire _3162_;
 wire _3163_;
 wire _3164_;
 wire _3165_;
 wire _3166_;
 wire _3167_;
 wire _3168_;
 wire _3169_;
 wire _3170_;
 wire _3171_;
 wire _3172_;
 wire _3173_;
 wire _3174_;
 wire _3175_;
 wire _3176_;
 wire _3177_;
 wire _3178_;
 wire _3179_;
 wire _3180_;
 wire _3181_;
 wire _3182_;
 wire _3183_;
 wire _3184_;
 wire _3185_;
 wire _3186_;
 wire _3187_;
 wire _3188_;
 wire _3189_;
 wire _3190_;
 wire _3191_;
 wire _3192_;
 wire _3193_;
 wire _3194_;
 wire _3195_;
 wire _3196_;
 wire _3197_;
 wire _3198_;
 wire _3199_;
 wire _3200_;
 wire _3201_;
 wire _3202_;
 wire _3203_;
 wire _3204_;
 wire _3205_;
 wire _3206_;
 wire _3207_;
 wire _3208_;
 wire _3209_;
 wire _3210_;
 wire _3211_;
 wire _3212_;
 wire _3213_;
 wire _3214_;
 wire _3215_;
 wire _3216_;
 wire _3217_;
 wire _3218_;
 wire _3219_;
 wire _3220_;
 wire _3221_;
 wire _3222_;
 wire _3223_;
 wire _3224_;
 wire _3225_;
 wire _3226_;
 wire _3227_;
 wire _3228_;
 wire _3229_;
 wire _3230_;
 wire _3231_;
 wire _3232_;
 wire _3233_;
 wire _3234_;
 wire _3235_;
 wire _3236_;
 wire _3237_;
 wire _3238_;
 wire _3239_;
 wire _3240_;
 wire _3241_;
 wire _3242_;
 wire _3243_;
 wire _3244_;
 wire _3245_;
 wire _3246_;
 wire _3247_;
 wire _3248_;
 wire _3249_;
 wire _3250_;
 wire _3251_;
 wire _3252_;
 wire _3253_;
 wire _3254_;
 wire _3255_;
 wire _3256_;
 wire _3257_;
 wire _3258_;
 wire _3259_;
 wire _3260_;
 wire _3261_;
 wire _3262_;
 wire _3263_;
 wire _3264_;
 wire _3265_;
 wire _3266_;
 wire _3267_;
 wire _3268_;
 wire _3269_;
 wire _3270_;
 wire _3271_;
 wire _3272_;
 wire _3273_;
 wire _3274_;
 wire _3275_;
 wire _3276_;
 wire _3277_;
 wire _3278_;
 wire _3279_;
 wire _3280_;
 wire _3281_;
 wire _3282_;
 wire _3283_;
 wire _3284_;
 wire _3285_;
 wire _3286_;
 wire _3287_;
 wire _3288_;
 wire _3289_;
 wire _3290_;
 wire _3291_;
 wire _3292_;
 wire _3293_;
 wire _3294_;
 wire _3295_;
 wire _3296_;
 wire _3297_;
 wire _3298_;
 wire _3299_;
 wire _3300_;
 wire _3301_;
 wire _3302_;
 wire _3303_;
 wire _3304_;
 wire _3305_;
 wire _3306_;
 wire _3307_;
 wire _3308_;
 wire _3309_;
 wire _3310_;
 wire _3311_;
 wire _3312_;
 wire _3313_;
 wire _3314_;
 wire _3315_;
 wire _3316_;
 wire _3317_;
 wire _3318_;
 wire _3319_;
 wire _3320_;
 wire _3321_;
 wire _3322_;
 wire _3323_;
 wire _3324_;
 wire _3325_;
 wire _3326_;
 wire _3327_;
 wire _3328_;
 wire _3329_;
 wire _3330_;
 wire _3331_;
 wire _3332_;
 wire _3333_;
 wire _3334_;
 wire _3335_;
 wire _3336_;
 wire _3337_;
 wire _3338_;
 wire _3339_;
 wire _3340_;
 wire _3341_;
 wire _3342_;
 wire _3343_;
 wire _3344_;
 wire _3345_;
 wire _3346_;
 wire _3347_;
 wire _3348_;
 wire _3349_;
 wire _3350_;
 wire _3351_;
 wire _3352_;
 wire _3353_;
 wire _3354_;
 wire _3355_;
 wire _3356_;
 wire _3357_;
 wire _3358_;
 wire _3359_;
 wire _3360_;
 wire _3361_;
 wire _3362_;
 wire _3363_;
 wire _3364_;
 wire _3365_;
 wire _3366_;
 wire _3367_;
 wire _3368_;
 wire _3369_;
 wire _3370_;
 wire _3371_;
 wire _3372_;
 wire _3373_;
 wire _3374_;
 wire _3375_;
 wire _3376_;
 wire _3377_;
 wire _3378_;
 wire _3379_;
 wire _3380_;
 wire _3381_;
 wire _3382_;
 wire _3383_;
 wire _3384_;
 wire _3385_;
 wire _3386_;
 wire _3387_;
 wire _3388_;
 wire _3389_;
 wire _3390_;
 wire _3391_;
 wire _3392_;
 wire _3393_;
 wire _3394_;
 wire _3395_;
 wire _3396_;
 wire _3397_;
 wire _3398_;
 wire _3399_;
 wire _3400_;
 wire _3401_;
 wire _3402_;
 wire _3403_;
 wire _3404_;
 wire _3405_;
 wire _3406_;
 wire _3407_;
 wire _3408_;
 wire _3409_;
 wire _3410_;
 wire _3411_;
 wire _3412_;
 wire _3413_;
 wire _3414_;
 wire _3415_;
 wire _3416_;
 wire _3417_;
 wire _3418_;
 wire _3419_;
 wire _3420_;
 wire _3421_;
 wire _3422_;
 wire _3423_;
 wire _3424_;
 wire _3425_;
 wire _3426_;
 wire _3427_;
 wire _3428_;
 wire _3429_;
 wire _3430_;
 wire _3431_;
 wire _3432_;
 wire _3433_;
 wire _3434_;
 wire _3435_;
 wire _3436_;
 wire _3437_;
 wire _3438_;
 wire _3439_;
 wire _3440_;
 wire _3441_;
 wire _3442_;
 wire _3443_;
 wire _3444_;
 wire _3445_;
 wire _3446_;
 wire _3447_;
 wire _3448_;
 wire _3449_;
 wire _3450_;
 wire _3451_;
 wire _3452_;
 wire _3453_;
 wire _3454_;
 wire _3455_;
 wire _3456_;
 wire _3457_;
 wire _3458_;
 wire _3459_;
 wire _3460_;
 wire _3461_;
 wire _3462_;
 wire _3463_;
 wire _3464_;
 wire _3465_;
 wire _3466_;
 wire _3467_;
 wire _3468_;
 wire _3469_;
 wire _3470_;
 wire _3471_;
 wire _3472_;
 wire _3473_;
 wire _3474_;
 wire _3475_;
 wire _3476_;
 wire _3477_;
 wire _3478_;
 wire _3479_;
 wire _3480_;
 wire _3481_;
 wire _3482_;
 wire _3483_;
 wire _3484_;
 wire _3485_;
 wire _3486_;
 wire _3487_;
 wire _3488_;
 wire _3489_;
 wire _3490_;
 wire _3491_;
 wire _3492_;
 wire _3493_;
 wire _3494_;
 wire _3495_;
 wire _3496_;
 wire _3497_;
 wire _3498_;
 wire _3499_;
 wire _3500_;
 wire _3501_;
 wire _3502_;
 wire _3503_;
 wire _3504_;
 wire _3505_;
 wire _3506_;
 wire _3507_;
 wire _3508_;
 wire _3509_;
 wire _3510_;
 wire _3511_;
 wire _3512_;
 wire _3513_;
 wire _3514_;
 wire _3515_;
 wire _3516_;
 wire _3517_;
 wire _3518_;
 wire _3519_;
 wire _3520_;
 wire _3521_;
 wire _3522_;
 wire _3523_;
 wire _3524_;
 wire _3525_;
 wire _3526_;
 wire _3527_;
 wire _3528_;
 wire _3529_;
 wire _3530_;
 wire _3531_;
 wire _3532_;
 wire _3533_;
 wire _3534_;
 wire _3535_;
 wire _3536_;
 wire _3537_;
 wire _3538_;
 wire _3539_;
 wire _3540_;
 wire _3541_;
 wire _3542_;
 wire _3543_;
 wire _3544_;
 wire _3545_;
 wire _3546_;
 wire _3547_;
 wire _3548_;
 wire _3549_;
 wire _3550_;
 wire _3551_;
 wire _3552_;
 wire _3553_;
 wire _3554_;
 wire _3555_;
 wire _3556_;
 wire _3557_;
 wire _3558_;
 wire _3559_;
 wire _3560_;
 wire _3561_;
 wire _3562_;
 wire _3563_;
 wire _3564_;
 wire _3565_;
 wire _3566_;
 wire _3567_;
 wire _3568_;
 wire _3569_;
 wire _3570_;
 wire _3571_;
 wire _3572_;
 wire _3573_;
 wire _3574_;
 wire _3575_;
 wire _3576_;
 wire _3577_;
 wire _3578_;
 wire _3579_;
 wire _3580_;
 wire _3581_;
 wire _3582_;
 wire _3583_;
 wire _3584_;
 wire _3585_;
 wire _3586_;
 wire _3587_;
 wire _3588_;
 wire _3589_;
 wire _3590_;
 wire _3591_;
 wire _3592_;
 wire _3593_;
 wire _3594_;
 wire _3595_;
 wire _3596_;
 wire _3597_;
 wire _3598_;
 wire _3599_;
 wire _3600_;
 wire _3601_;
 wire _3602_;
 wire _3603_;
 wire _3604_;
 wire _3605_;
 wire _3606_;
 wire _3607_;
 wire _3608_;
 wire _3609_;
 wire _3610_;
 wire _3611_;
 wire _3612_;
 wire _3613_;
 wire _3614_;
 wire _3615_;
 wire _3616_;
 wire _3617_;
 wire _3618_;
 wire _3619_;
 wire _3620_;
 wire _3621_;
 wire _3622_;
 wire _3623_;
 wire _3624_;
 wire _3625_;
 wire _3626_;
 wire _3627_;
 wire _3628_;
 wire _3629_;
 wire _3630_;
 wire _3631_;
 wire _3632_;
 wire _3633_;
 wire _3634_;
 wire _3635_;
 wire _3636_;
 wire _3637_;
 wire _3638_;
 wire _3639_;
 wire _3640_;
 wire _3641_;
 wire _3642_;
 wire _3643_;
 wire _3644_;
 wire _3645_;
 wire _3646_;
 wire _3647_;
 wire _3648_;
 wire _3649_;
 wire _3650_;
 wire _3651_;
 wire _3652_;
 wire _3653_;
 wire _3654_;
 wire _3655_;
 wire _3656_;
 wire _3657_;
 wire _3658_;
 wire _3659_;
 wire _3660_;
 wire _3661_;
 wire _3662_;
 wire _3663_;
 wire _3664_;
 wire _3665_;
 wire _3666_;
 wire _3667_;
 wire _3668_;
 wire _3669_;
 wire _3670_;
 wire _3671_;
 wire _3672_;
 wire _3673_;
 wire _3674_;
 wire _3675_;
 wire _3676_;
 wire _3677_;
 wire _3678_;
 wire _3679_;
 wire _3680_;
 wire _3681_;
 wire _3682_;
 wire _3683_;
 wire _3684_;
 wire _3685_;
 wire _3686_;
 wire _3687_;
 wire _3688_;
 wire _3689_;
 wire _3690_;
 wire _3691_;
 wire _3692_;
 wire _3693_;
 wire _3694_;
 wire _3695_;
 wire _3696_;
 wire _3697_;
 wire _3698_;
 wire _3699_;
 wire _3700_;
 wire _3701_;
 wire _3702_;
 wire _3703_;
 wire _3704_;
 wire _3705_;
 wire _3706_;
 wire _3707_;
 wire _3708_;
 wire _3709_;
 wire _3710_;
 wire _3711_;
 wire _3712_;
 wire _3713_;
 wire _3714_;
 wire _3715_;
 wire _3716_;
 wire _3717_;
 wire _3718_;
 wire _3719_;
 wire _3720_;
 wire _3721_;
 wire _3722_;
 wire _3723_;
 wire _3724_;
 wire _3725_;
 wire _3726_;
 wire _3727_;
 wire _3728_;
 wire _3729_;
 wire _3730_;
 wire _3731_;
 wire _3732_;
 wire _3733_;
 wire _3734_;
 wire _3735_;
 wire _3736_;
 wire _3737_;
 wire _3738_;
 wire _3739_;
 wire _3740_;
 wire _3741_;
 wire _3742_;
 wire _3743_;
 wire _3744_;
 wire _3745_;
 wire _3746_;
 wire _3747_;
 wire _3748_;
 wire _3749_;
 wire _3750_;
 wire _3751_;
 wire _3752_;
 wire _3753_;
 wire _3754_;
 wire clknet_0_clk;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire clknet_leaf_0_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_52_clk;
 wire clknet_leaf_53_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_55_clk;
 wire clknet_leaf_56_clk;
 wire clknet_leaf_57_clk;
 wire clknet_leaf_58_clk;
 wire clknet_leaf_59_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire \debug_rd_r[0] ;
 wire \debug_rd_r[1] ;
 wire \debug_rd_r[2] ;
 wire \debug_rd_r[3] ;
 wire debug_register_data;
 wire \gpio_out[0] ;
 wire \gpio_out[1] ;
 wire \gpio_out[2] ;
 wire \gpio_out[3] ;
 wire \gpio_out[4] ;
 wire \gpio_out[5] ;
 wire \gpio_out[6] ;
 wire \gpio_out[7] ;
 wire \gpio_out_sel[0] ;
 wire \gpio_out_sel[1] ;
 wire \gpio_out_sel[2] ;
 wire \gpio_out_sel[3] ;
 wire \gpio_out_sel[4] ;
 wire \gpio_out_sel[5] ;
 wire \gpio_out_sel[6] ;
 wire \gpio_out_sel[7] ;
 wire \i_debug_uart_tx.cycle_counter[0] ;
 wire \i_debug_uart_tx.cycle_counter[1] ;
 wire \i_debug_uart_tx.cycle_counter[2] ;
 wire \i_debug_uart_tx.cycle_counter[3] ;
 wire \i_debug_uart_tx.cycle_counter[4] ;
 wire \i_debug_uart_tx.data_to_send[0] ;
 wire \i_debug_uart_tx.data_to_send[1] ;
 wire \i_debug_uart_tx.data_to_send[2] ;
 wire \i_debug_uart_tx.data_to_send[3] ;
 wire \i_debug_uart_tx.data_to_send[4] ;
 wire \i_debug_uart_tx.data_to_send[5] ;
 wire \i_debug_uart_tx.data_to_send[6] ;
 wire \i_debug_uart_tx.data_to_send[7] ;
 wire \i_debug_uart_tx.fsm_state[0] ;
 wire \i_debug_uart_tx.fsm_state[1] ;
 wire \i_debug_uart_tx.fsm_state[2] ;
 wire \i_debug_uart_tx.fsm_state[3] ;
 wire \i_debug_uart_tx.resetn ;
 wire \i_debug_uart_tx.txd_reg ;
 wire \i_debug_uart_tx.uart_tx_data[0] ;
 wire \i_debug_uart_tx.uart_tx_data[1] ;
 wire \i_debug_uart_tx.uart_tx_data[2] ;
 wire \i_debug_uart_tx.uart_tx_data[3] ;
 wire \i_debug_uart_tx.uart_tx_data[4] ;
 wire \i_debug_uart_tx.uart_tx_data[5] ;
 wire \i_debug_uart_tx.uart_tx_data[6] ;
 wire \i_debug_uart_tx.uart_tx_data[7] ;
 wire \i_spi.bits_remaining[0] ;
 wire \i_spi.bits_remaining[1] ;
 wire \i_spi.bits_remaining[2] ;
 wire \i_spi.bits_remaining[3] ;
 wire \i_spi.busy ;
 wire \i_spi.clock_count[0] ;
 wire \i_spi.clock_count[1] ;
 wire \i_spi.clock_divider[0] ;
 wire \i_spi.clock_divider[1] ;
 wire \i_spi.data[0] ;
 wire \i_spi.data[1] ;
 wire \i_spi.data[2] ;
 wire \i_spi.data[3] ;
 wire \i_spi.data[4] ;
 wire \i_spi.data[5] ;
 wire \i_spi.data[6] ;
 wire \i_spi.data[7] ;
 wire \i_spi.dc_in ;
 wire \i_spi.end_txn ;
 wire \i_spi.end_txn_reg ;
 wire \i_spi.read_latency ;
 wire \i_spi.spi_clk_out ;
 wire \i_spi.spi_dc ;
 wire \i_spi.spi_select ;
 wire \i_tinyqv.cpu.additional_mem_ops[0] ;
 wire \i_tinyqv.cpu.additional_mem_ops[1] ;
 wire \i_tinyqv.cpu.additional_mem_ops[2] ;
 wire \i_tinyqv.cpu.alu_op[0] ;
 wire \i_tinyqv.cpu.alu_op[1] ;
 wire \i_tinyqv.cpu.alu_op[2] ;
 wire \i_tinyqv.cpu.alu_op[3] ;
 wire \i_tinyqv.cpu.counter[2] ;
 wire \i_tinyqv.cpu.counter[3] ;
 wire \i_tinyqv.cpu.counter[4] ;
 wire \i_tinyqv.cpu.data_addr[0] ;
 wire \i_tinyqv.cpu.data_addr[10] ;
 wire \i_tinyqv.cpu.data_addr[11] ;
 wire \i_tinyqv.cpu.data_addr[12] ;
 wire \i_tinyqv.cpu.data_addr[13] ;
 wire \i_tinyqv.cpu.data_addr[14] ;
 wire \i_tinyqv.cpu.data_addr[15] ;
 wire \i_tinyqv.cpu.data_addr[16] ;
 wire \i_tinyqv.cpu.data_addr[17] ;
 wire \i_tinyqv.cpu.data_addr[18] ;
 wire \i_tinyqv.cpu.data_addr[19] ;
 wire \i_tinyqv.cpu.data_addr[1] ;
 wire \i_tinyqv.cpu.data_addr[20] ;
 wire \i_tinyqv.cpu.data_addr[21] ;
 wire \i_tinyqv.cpu.data_addr[22] ;
 wire \i_tinyqv.cpu.data_addr[23] ;
 wire \i_tinyqv.cpu.data_addr[24] ;
 wire \i_tinyqv.cpu.data_addr[25] ;
 wire \i_tinyqv.cpu.data_addr[26] ;
 wire \i_tinyqv.cpu.data_addr[27] ;
 wire \i_tinyqv.cpu.data_addr[2] ;
 wire \i_tinyqv.cpu.data_addr[3] ;
 wire \i_tinyqv.cpu.data_addr[4] ;
 wire \i_tinyqv.cpu.data_addr[5] ;
 wire \i_tinyqv.cpu.data_addr[6] ;
 wire \i_tinyqv.cpu.data_addr[7] ;
 wire \i_tinyqv.cpu.data_addr[8] ;
 wire \i_tinyqv.cpu.data_addr[9] ;
 wire \i_tinyqv.cpu.data_continue ;
 wire \i_tinyqv.cpu.data_out[10] ;
 wire \i_tinyqv.cpu.data_out[11] ;
 wire \i_tinyqv.cpu.data_out[12] ;
 wire \i_tinyqv.cpu.data_out[13] ;
 wire \i_tinyqv.cpu.data_out[14] ;
 wire \i_tinyqv.cpu.data_out[15] ;
 wire \i_tinyqv.cpu.data_out[16] ;
 wire \i_tinyqv.cpu.data_out[17] ;
 wire \i_tinyqv.cpu.data_out[18] ;
 wire \i_tinyqv.cpu.data_out[19] ;
 wire \i_tinyqv.cpu.data_out[20] ;
 wire \i_tinyqv.cpu.data_out[21] ;
 wire \i_tinyqv.cpu.data_out[22] ;
 wire \i_tinyqv.cpu.data_out[23] ;
 wire \i_tinyqv.cpu.data_out[24] ;
 wire \i_tinyqv.cpu.data_out[25] ;
 wire \i_tinyqv.cpu.data_out[26] ;
 wire \i_tinyqv.cpu.data_out[27] ;
 wire \i_tinyqv.cpu.data_out[28] ;
 wire \i_tinyqv.cpu.data_out[29] ;
 wire \i_tinyqv.cpu.data_out[30] ;
 wire \i_tinyqv.cpu.data_out[31] ;
 wire \i_tinyqv.cpu.data_read_n[0] ;
 wire \i_tinyqv.cpu.data_read_n[1] ;
 wire \i_tinyqv.cpu.data_ready_core ;
 wire \i_tinyqv.cpu.data_ready_latch ;
 wire \i_tinyqv.cpu.data_write_n[0] ;
 wire \i_tinyqv.cpu.data_write_n[1] ;
 wire \i_tinyqv.cpu.debug_instr_valid ;
 wire \i_tinyqv.cpu.debug_rd[0] ;
 wire \i_tinyqv.cpu.debug_rd[1] ;
 wire \i_tinyqv.cpu.debug_rd[2] ;
 wire \i_tinyqv.cpu.debug_rd[3] ;
 wire \i_tinyqv.cpu.i_core.cmp ;
 wire \i_tinyqv.cpu.i_core.cmp_out ;
 wire \i_tinyqv.cpu.i_core.cy ;
 wire \i_tinyqv.cpu.i_core.cy_out ;
 wire \i_tinyqv.cpu.i_core.cycle[0] ;
 wire \i_tinyqv.cpu.i_core.cycle[1] ;
 wire \i_tinyqv.cpu.i_core.cycle_count[0] ;
 wire \i_tinyqv.cpu.i_core.cycle_count[1] ;
 wire \i_tinyqv.cpu.i_core.cycle_count[2] ;
 wire \i_tinyqv.cpu.i_core.cycle_count[3] ;
 wire \i_tinyqv.cpu.i_core.cycle_count_wide[4] ;
 wire \i_tinyqv.cpu.i_core.cycle_count_wide[5] ;
 wire \i_tinyqv.cpu.i_core.cycle_count_wide[6] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.cy ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[10] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[11] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[12] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[13] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[14] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[15] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[16] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[17] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[18] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[19] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[20] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[21] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[22] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[23] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[24] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[25] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[26] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[27] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[28] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[29] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[30] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[31] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[4] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[5] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[6] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[7] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[8] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[9] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.register[0] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.register[11] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.register[12] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.register[13] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.register[14] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.register[15] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.register[16] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.register[17] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.register[18] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.register[19] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.register[1] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.register[20] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.register[21] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.register[22] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.register[23] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.register[24] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.register[25] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.register[26] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.register[27] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.register[28] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.register[29] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.register[2] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.register[30] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.register[31] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.register[3] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.rstn ;
 wire \i_tinyqv.cpu.i_core.i_instrret.add ;
 wire \i_tinyqv.cpu.i_core.i_instrret.cy ;
 wire \i_tinyqv.cpu.i_core.i_instrret.data[0] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.data[1] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.data[2] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.data[3] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[10] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[11] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[12] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[13] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[14] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[15] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[16] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[17] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[18] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[19] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[20] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[21] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[22] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[23] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[24] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[25] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[26] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[27] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[28] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[29] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[30] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[31] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[4] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[5] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[6] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[7] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[8] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[9] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.register[0] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.register[10] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.register[11] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.register[12] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.register[13] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.register[14] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.register[15] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.register[16] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.register[17] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.register[18] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.register[19] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.register[1] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.register[20] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.register[21] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.register[22] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.register[23] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.register[24] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.register[25] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.register[26] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.register[27] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.register[28] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.register[29] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.register[2] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.register[30] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.register[31] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.register[3] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.register[8] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.register[9] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.reg_buf[10] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.reg_buf[11] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.reg_buf[12] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.reg_buf[13] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.reg_buf[14] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.reg_buf[15] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.reg_buf[16] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.reg_buf[17] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.reg_buf[18] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.reg_buf[19] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.reg_buf[20] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.reg_buf[21] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.reg_buf[22] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.reg_buf[23] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.reg_buf[24] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.reg_buf[25] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.reg_buf[26] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.reg_buf[27] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.reg_buf[28] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.reg_buf[29] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.reg_buf[30] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.reg_buf[31] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.reg_buf[4] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.reg_buf[5] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.reg_buf[6] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.reg_buf[7] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.reg_buf[8] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.reg_buf[9] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.reg_buf[10] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.reg_buf[11] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.reg_buf[12] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.reg_buf[13] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.reg_buf[14] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.reg_buf[15] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.reg_buf[16] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.reg_buf[17] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.reg_buf[18] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.reg_buf[19] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.reg_buf[20] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.reg_buf[21] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.reg_buf[22] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.reg_buf[23] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.reg_buf[24] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.reg_buf[25] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.reg_buf[26] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.reg_buf[27] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.reg_buf[28] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.reg_buf[29] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.reg_buf[30] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.reg_buf[31] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.reg_buf[4] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.reg_buf[5] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.reg_buf[6] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.reg_buf[7] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.reg_buf[8] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.reg_buf[9] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.reg_buf[10] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.reg_buf[11] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.reg_buf[12] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.reg_buf[13] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.reg_buf[14] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.reg_buf[15] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.reg_buf[16] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.reg_buf[17] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.reg_buf[18] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.reg_buf[19] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.reg_buf[20] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.reg_buf[21] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.reg_buf[22] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.reg_buf[23] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.reg_buf[24] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.reg_buf[25] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.reg_buf[26] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.reg_buf[27] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.reg_buf[28] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.reg_buf[29] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.reg_buf[30] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.reg_buf[31] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.reg_buf[4] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.reg_buf[5] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.reg_buf[6] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.reg_buf[7] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.reg_buf[8] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.reg_buf[9] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.reg_buf[10] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.reg_buf[11] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.reg_buf[12] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.reg_buf[13] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.reg_buf[14] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.reg_buf[15] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.reg_buf[16] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.reg_buf[17] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.reg_buf[18] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.reg_buf[19] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.reg_buf[20] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.reg_buf[21] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.reg_buf[22] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.reg_buf[23] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.reg_buf[24] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.reg_buf[25] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.reg_buf[26] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.reg_buf[27] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.reg_buf[28] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.reg_buf[29] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.reg_buf[30] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.reg_buf[31] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.reg_buf[4] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.reg_buf[5] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.reg_buf[6] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.reg_buf[7] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.reg_buf[8] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.reg_buf[9] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.reg_buf[10] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.reg_buf[11] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.reg_buf[12] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.reg_buf[13] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.reg_buf[14] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.reg_buf[15] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.reg_buf[16] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.reg_buf[17] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.reg_buf[18] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.reg_buf[19] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.reg_buf[20] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.reg_buf[21] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.reg_buf[22] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.reg_buf[23] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.reg_buf[24] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.reg_buf[25] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.reg_buf[26] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.reg_buf[27] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.reg_buf[28] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.reg_buf[29] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.reg_buf[30] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.reg_buf[31] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.reg_buf[4] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.reg_buf[5] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.reg_buf[6] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.reg_buf[7] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.reg_buf[8] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.reg_buf[9] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.reg_buf[10] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.reg_buf[11] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.reg_buf[12] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.reg_buf[13] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.reg_buf[14] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.reg_buf[15] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.reg_buf[16] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.reg_buf[17] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.reg_buf[18] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.reg_buf[19] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.reg_buf[20] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.reg_buf[21] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.reg_buf[22] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.reg_buf[23] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.reg_buf[24] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.reg_buf[25] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.reg_buf[26] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.reg_buf[27] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.reg_buf[28] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.reg_buf[29] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.reg_buf[30] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.reg_buf[31] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.reg_buf[4] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.reg_buf[5] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.reg_buf[6] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.reg_buf[7] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.reg_buf[8] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.reg_buf[9] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.reg_buf[10] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.reg_buf[11] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.reg_buf[12] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.reg_buf[13] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.reg_buf[14] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.reg_buf[15] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.reg_buf[16] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.reg_buf[17] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.reg_buf[18] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.reg_buf[19] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.reg_buf[20] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.reg_buf[21] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.reg_buf[22] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.reg_buf[23] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.reg_buf[24] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.reg_buf[25] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.reg_buf[26] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.reg_buf[27] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.reg_buf[28] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.reg_buf[29] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.reg_buf[30] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.reg_buf[31] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.reg_buf[4] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.reg_buf[5] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.reg_buf[6] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.reg_buf[7] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.reg_buf[8] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.reg_buf[9] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.reg_buf[10] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.reg_buf[11] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.reg_buf[12] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.reg_buf[13] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.reg_buf[14] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.reg_buf[15] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.reg_buf[16] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.reg_buf[17] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.reg_buf[18] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.reg_buf[19] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.reg_buf[20] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.reg_buf[21] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.reg_buf[22] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.reg_buf[23] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.reg_buf[24] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.reg_buf[25] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.reg_buf[26] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.reg_buf[27] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.reg_buf[28] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.reg_buf[29] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.reg_buf[30] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.reg_buf[31] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.reg_buf[4] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.reg_buf[5] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.reg_buf[6] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.reg_buf[7] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.reg_buf[8] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.reg_buf[9] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.reg_buf[10] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.reg_buf[11] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.reg_buf[12] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.reg_buf[13] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.reg_buf[14] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.reg_buf[15] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.reg_buf[16] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.reg_buf[17] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.reg_buf[18] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.reg_buf[19] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.reg_buf[20] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.reg_buf[21] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.reg_buf[22] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.reg_buf[23] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.reg_buf[24] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.reg_buf[25] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.reg_buf[26] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.reg_buf[27] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.reg_buf[28] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.reg_buf[29] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.reg_buf[30] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.reg_buf[31] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.reg_buf[4] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.reg_buf[5] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.reg_buf[6] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.reg_buf[7] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.reg_buf[8] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.reg_buf[9] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.reg_buf[10] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.reg_buf[11] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.reg_buf[12] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.reg_buf[13] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.reg_buf[14] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.reg_buf[15] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.reg_buf[16] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.reg_buf[17] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.reg_buf[18] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.reg_buf[19] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.reg_buf[20] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.reg_buf[21] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.reg_buf[22] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.reg_buf[23] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.reg_buf[24] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.reg_buf[25] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.reg_buf[26] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.reg_buf[27] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.reg_buf[28] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.reg_buf[29] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.reg_buf[30] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.reg_buf[31] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.reg_buf[4] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.reg_buf[5] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.reg_buf[6] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.reg_buf[7] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.reg_buf[8] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.reg_buf[9] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.reg_buf[10] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.reg_buf[11] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.reg_buf[12] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.reg_buf[13] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.reg_buf[14] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.reg_buf[15] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.reg_buf[16] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.reg_buf[17] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.reg_buf[18] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.reg_buf[19] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.reg_buf[20] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.reg_buf[21] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.reg_buf[22] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.reg_buf[23] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.reg_buf[24] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.reg_buf[25] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.reg_buf[26] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.reg_buf[27] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.reg_buf[28] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.reg_buf[29] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.reg_buf[30] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.reg_buf[31] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.reg_buf[4] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.reg_buf[5] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.reg_buf[6] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.reg_buf[7] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.reg_buf[8] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.reg_buf[9] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.reg_buf[10] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.reg_buf[11] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.reg_buf[12] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.reg_buf[13] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.reg_buf[14] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.reg_buf[15] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.reg_buf[16] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.reg_buf[17] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.reg_buf[18] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.reg_buf[19] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.reg_buf[20] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.reg_buf[21] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.reg_buf[22] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.reg_buf[23] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.reg_buf[24] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.reg_buf[25] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.reg_buf[26] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.reg_buf[27] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.reg_buf[28] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.reg_buf[29] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.reg_buf[30] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.reg_buf[31] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.reg_buf[4] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.reg_buf[5] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.reg_buf[6] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.reg_buf[7] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.reg_buf[8] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.reg_buf[9] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.reg_buf[10] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.reg_buf[11] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.reg_buf[12] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.reg_buf[13] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.reg_buf[14] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.reg_buf[15] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.reg_buf[16] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.reg_buf[17] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.reg_buf[18] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.reg_buf[19] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.reg_buf[20] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.reg_buf[21] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.reg_buf[22] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.reg_buf[23] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.reg_buf[24] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.reg_buf[25] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.reg_buf[26] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.reg_buf[27] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.reg_buf[28] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.reg_buf[29] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.reg_buf[30] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.reg_buf[31] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.reg_buf[4] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.reg_buf[5] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.reg_buf[6] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.reg_buf[7] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.reg_buf[8] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.reg_buf[9] ;
 wire \i_tinyqv.cpu.i_core.i_registers.rd[0] ;
 wire \i_tinyqv.cpu.i_core.i_registers.rd[1] ;
 wire \i_tinyqv.cpu.i_core.i_registers.rd[2] ;
 wire \i_tinyqv.cpu.i_core.i_registers.rd[3] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[10][0] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[10][1] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[10][2] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[10][3] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[11][0] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[11][1] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[11][2] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[11][3] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[12][0] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[12][1] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[12][2] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[12][3] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[13][0] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[13][1] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[13][2] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[13][3] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[14][0] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[14][1] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[14][2] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[14][3] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[15][0] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[15][1] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[15][2] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[15][3] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[1][0] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[1][1] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[1][2] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[1][3] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[2][0] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[2][1] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[2][2] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[2][3] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[5][0] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[5][1] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[5][2] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[5][3] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[6][0] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[6][1] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[6][2] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[6][3] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[7][0] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[7][1] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[7][2] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[7][3] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[8][0] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[8][1] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[8][2] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[8][3] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[9][0] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[9][1] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[9][2] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[9][3] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[10][0] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[10][10] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[10][11] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[10][12] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[10][13] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[10][14] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[10][15] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[10][16] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[10][17] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[10][18] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[10][19] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[10][1] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[10][20] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[10][21] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[10][22] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[10][23] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[10][24] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[10][25] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[10][26] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[10][27] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[10][28] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[10][29] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[10][2] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[10][30] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[10][31] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[10][3] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[10][8] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[10][9] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[11][0] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[11][10] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[11][11] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[11][12] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[11][13] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[11][14] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[11][15] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[11][16] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[11][17] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[11][18] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[11][19] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[11][1] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[11][20] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[11][21] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[11][22] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[11][23] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[11][24] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[11][25] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[11][26] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[11][27] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[11][28] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[11][29] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[11][2] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[11][30] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[11][31] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[11][3] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[11][8] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[11][9] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[12][0] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[12][10] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[12][11] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[12][12] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[12][13] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[12][14] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[12][15] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[12][16] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[12][17] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[12][18] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[12][19] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[12][1] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[12][20] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[12][21] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[12][22] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[12][23] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[12][24] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[12][25] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[12][26] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[12][27] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[12][28] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[12][29] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[12][2] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[12][30] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[12][31] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[12][3] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[12][8] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[12][9] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[13][0] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[13][10] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[13][11] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[13][12] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[13][13] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[13][14] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[13][15] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[13][16] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[13][17] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[13][18] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[13][19] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[13][1] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[13][20] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[13][21] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[13][22] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[13][23] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[13][24] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[13][25] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[13][26] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[13][27] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[13][28] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[13][29] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[13][2] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[13][30] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[13][31] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[13][3] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[13][8] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[13][9] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[14][0] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[14][10] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[14][11] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[14][12] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[14][13] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[14][14] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[14][15] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[14][16] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[14][17] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[14][18] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[14][19] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[14][1] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[14][20] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[14][21] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[14][22] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[14][23] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[14][24] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[14][25] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[14][26] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[14][27] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[14][28] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[14][29] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[14][2] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[14][30] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[14][31] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[14][3] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[14][8] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[14][9] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[15][0] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[15][10] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[15][11] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[15][12] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[15][13] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[15][14] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[15][15] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[15][16] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[15][17] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[15][18] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[15][19] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[15][1] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[15][20] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[15][21] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[15][22] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[15][23] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[15][24] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[15][25] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[15][26] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[15][27] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[15][28] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[15][29] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[15][2] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[15][30] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[15][31] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[15][3] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[15][8] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[15][9] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[1][0] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[1][10] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[1][11] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[1][12] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[1][13] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[1][14] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[1][15] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[1][16] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[1][17] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[1][18] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[1][19] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[1][1] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[1][20] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[1][21] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[1][22] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[1][23] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[1][24] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[1][25] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[1][26] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[1][27] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[1][28] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[1][29] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[1][2] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[1][30] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[1][31] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[1][3] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[1][8] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[1][9] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[2][0] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[2][10] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[2][11] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[2][12] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[2][13] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[2][14] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[2][15] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[2][16] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[2][17] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[2][18] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[2][19] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[2][1] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[2][20] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[2][21] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[2][22] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[2][23] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[2][24] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[2][25] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[2][26] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[2][27] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[2][28] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[2][29] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[2][2] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[2][30] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[2][31] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[2][3] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[2][8] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[2][9] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[5][0] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[5][10] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[5][11] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[5][12] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[5][13] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[5][14] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[5][15] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[5][16] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[5][17] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[5][18] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[5][19] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[5][1] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[5][20] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[5][21] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[5][22] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[5][23] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[5][24] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[5][25] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[5][26] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[5][27] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[5][28] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[5][29] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[5][2] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[5][30] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[5][31] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[5][3] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[5][8] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[5][9] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[6][0] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[6][10] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[6][11] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[6][12] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[6][13] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[6][14] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[6][15] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[6][16] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[6][17] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[6][18] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[6][19] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[6][1] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[6][20] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[6][21] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[6][22] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[6][23] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[6][24] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[6][25] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[6][26] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[6][27] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[6][28] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[6][29] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[6][2] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[6][30] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[6][31] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[6][3] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[6][8] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[6][9] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[7][0] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[7][10] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[7][11] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[7][12] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[7][13] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[7][14] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[7][15] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[7][16] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[7][17] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[7][18] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[7][19] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[7][1] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[7][20] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[7][21] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[7][22] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[7][23] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[7][24] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[7][25] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[7][26] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[7][27] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[7][28] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[7][29] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[7][2] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[7][30] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[7][31] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[7][3] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[7][8] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[7][9] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[8][0] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[8][10] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[8][11] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[8][12] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[8][13] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[8][14] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[8][15] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[8][16] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[8][17] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[8][18] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[8][19] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[8][1] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[8][20] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[8][21] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[8][22] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[8][23] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[8][24] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[8][25] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[8][26] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[8][27] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[8][28] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[8][29] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[8][2] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[8][30] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[8][31] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[8][3] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[8][8] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[8][9] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[9][0] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[9][10] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[9][11] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[9][12] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[9][13] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[9][14] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[9][15] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[9][16] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[9][17] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[9][18] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[9][19] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[9][1] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[9][20] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[9][21] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[9][22] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[9][23] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[9][24] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[9][25] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[9][26] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[9][27] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[9][28] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[9][29] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[9][2] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[9][30] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[9][31] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[9][3] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[9][8] ;
 wire \i_tinyqv.cpu.i_core.i_registers.registers[9][9] ;
 wire \i_tinyqv.cpu.i_core.i_registers.rs1[0] ;
 wire \i_tinyqv.cpu.i_core.i_registers.rs1[1] ;
 wire \i_tinyqv.cpu.i_core.i_registers.rs1[2] ;
 wire \i_tinyqv.cpu.i_core.i_registers.rs1[3] ;
 wire \i_tinyqv.cpu.i_core.i_registers.rs2[0] ;
 wire \i_tinyqv.cpu.i_core.i_registers.rs2[1] ;
 wire \i_tinyqv.cpu.i_core.i_registers.rs2[2] ;
 wire \i_tinyqv.cpu.i_core.i_registers.rs2[3] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[0] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[10] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[11] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[12] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[13] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[14] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[15] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[16] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[17] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[18] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[19] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[1] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[20] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[21] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[22] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[23] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[24] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[25] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[26] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[27] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[28] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[29] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[2] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[30] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[31] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[3] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[4] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[5] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[6] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[7] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[8] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[9] ;
 wire \i_tinyqv.cpu.i_core.i_shift.adjusted_shift_amt[0] ;
 wire \i_tinyqv.cpu.i_core.i_shift.adjusted_shift_amt[1] ;
 wire \i_tinyqv.cpu.i_core.i_shift.b[2] ;
 wire \i_tinyqv.cpu.i_core.i_shift.b[3] ;
 wire \i_tinyqv.cpu.i_core.i_shift.b[4] ;
 wire \i_tinyqv.cpu.i_core.imm_lo[0] ;
 wire \i_tinyqv.cpu.i_core.imm_lo[10] ;
 wire \i_tinyqv.cpu.i_core.imm_lo[11] ;
 wire \i_tinyqv.cpu.i_core.imm_lo[1] ;
 wire \i_tinyqv.cpu.i_core.imm_lo[2] ;
 wire \i_tinyqv.cpu.i_core.imm_lo[3] ;
 wire \i_tinyqv.cpu.i_core.imm_lo[4] ;
 wire \i_tinyqv.cpu.i_core.imm_lo[5] ;
 wire \i_tinyqv.cpu.i_core.imm_lo[6] ;
 wire \i_tinyqv.cpu.i_core.imm_lo[7] ;
 wire \i_tinyqv.cpu.i_core.imm_lo[8] ;
 wire \i_tinyqv.cpu.i_core.imm_lo[9] ;
 wire \i_tinyqv.cpu.i_core.interrupt_req[0] ;
 wire \i_tinyqv.cpu.i_core.interrupt_req[1] ;
 wire \i_tinyqv.cpu.i_core.is_double_fault_r ;
 wire \i_tinyqv.cpu.i_core.is_interrupt ;
 wire \i_tinyqv.cpu.i_core.last_interrupt_req[0] ;
 wire \i_tinyqv.cpu.i_core.last_interrupt_req[1] ;
 wire \i_tinyqv.cpu.i_core.load_done ;
 wire \i_tinyqv.cpu.i_core.load_top_bit ;
 wire \i_tinyqv.cpu.i_core.mcause[0] ;
 wire \i_tinyqv.cpu.i_core.mcause[1] ;
 wire \i_tinyqv.cpu.i_core.mcause[3] ;
 wire \i_tinyqv.cpu.i_core.mcause[4] ;
 wire \i_tinyqv.cpu.i_core.mem_op[0] ;
 wire \i_tinyqv.cpu.i_core.mem_op[1] ;
 wire \i_tinyqv.cpu.i_core.mem_op[2] ;
 wire \i_tinyqv.cpu.i_core.mepc[0] ;
 wire \i_tinyqv.cpu.i_core.mepc[10] ;
 wire \i_tinyqv.cpu.i_core.mepc[11] ;
 wire \i_tinyqv.cpu.i_core.mepc[12] ;
 wire \i_tinyqv.cpu.i_core.mepc[13] ;
 wire \i_tinyqv.cpu.i_core.mepc[14] ;
 wire \i_tinyqv.cpu.i_core.mepc[15] ;
 wire \i_tinyqv.cpu.i_core.mepc[16] ;
 wire \i_tinyqv.cpu.i_core.mepc[17] ;
 wire \i_tinyqv.cpu.i_core.mepc[18] ;
 wire \i_tinyqv.cpu.i_core.mepc[19] ;
 wire \i_tinyqv.cpu.i_core.mepc[1] ;
 wire \i_tinyqv.cpu.i_core.mepc[20] ;
 wire \i_tinyqv.cpu.i_core.mepc[21] ;
 wire \i_tinyqv.cpu.i_core.mepc[22] ;
 wire \i_tinyqv.cpu.i_core.mepc[23] ;
 wire \i_tinyqv.cpu.i_core.mepc[2] ;
 wire \i_tinyqv.cpu.i_core.mepc[3] ;
 wire \i_tinyqv.cpu.i_core.mepc[4] ;
 wire \i_tinyqv.cpu.i_core.mepc[5] ;
 wire \i_tinyqv.cpu.i_core.mepc[6] ;
 wire \i_tinyqv.cpu.i_core.mepc[7] ;
 wire \i_tinyqv.cpu.i_core.mepc[8] ;
 wire \i_tinyqv.cpu.i_core.mepc[9] ;
 wire \i_tinyqv.cpu.i_core.mie[16] ;
 wire \i_tinyqv.cpu.i_core.mie[17] ;
 wire \i_tinyqv.cpu.i_core.mie[18] ;
 wire \i_tinyqv.cpu.i_core.mie[19] ;
 wire \i_tinyqv.cpu.i_core.mip[16] ;
 wire \i_tinyqv.cpu.i_core.mip[17] ;
 wire \i_tinyqv.cpu.i_core.mstatus_mie ;
 wire \i_tinyqv.cpu.i_core.mstatus_mpie ;
 wire \i_tinyqv.cpu.i_core.mstatus_mte ;
 wire \i_tinyqv.cpu.i_core.multiplier.accum[0] ;
 wire \i_tinyqv.cpu.i_core.multiplier.accum[10] ;
 wire \i_tinyqv.cpu.i_core.multiplier.accum[11] ;
 wire \i_tinyqv.cpu.i_core.multiplier.accum[12] ;
 wire \i_tinyqv.cpu.i_core.multiplier.accum[13] ;
 wire \i_tinyqv.cpu.i_core.multiplier.accum[14] ;
 wire \i_tinyqv.cpu.i_core.multiplier.accum[15] ;
 wire \i_tinyqv.cpu.i_core.multiplier.accum[1] ;
 wire \i_tinyqv.cpu.i_core.multiplier.accum[2] ;
 wire \i_tinyqv.cpu.i_core.multiplier.accum[3] ;
 wire \i_tinyqv.cpu.i_core.multiplier.accum[4] ;
 wire \i_tinyqv.cpu.i_core.multiplier.accum[5] ;
 wire \i_tinyqv.cpu.i_core.multiplier.accum[6] ;
 wire \i_tinyqv.cpu.i_core.multiplier.accum[7] ;
 wire \i_tinyqv.cpu.i_core.multiplier.accum[8] ;
 wire \i_tinyqv.cpu.i_core.multiplier.accum[9] ;
 wire \i_tinyqv.cpu.i_core.time_hi[0] ;
 wire \i_tinyqv.cpu.i_core.time_hi[1] ;
 wire \i_tinyqv.cpu.i_core.time_hi[2] ;
 wire \i_tinyqv.cpu.imm[12] ;
 wire \i_tinyqv.cpu.imm[13] ;
 wire \i_tinyqv.cpu.imm[14] ;
 wire \i_tinyqv.cpu.imm[15] ;
 wire \i_tinyqv.cpu.imm[16] ;
 wire \i_tinyqv.cpu.imm[17] ;
 wire \i_tinyqv.cpu.imm[18] ;
 wire \i_tinyqv.cpu.imm[19] ;
 wire \i_tinyqv.cpu.imm[20] ;
 wire \i_tinyqv.cpu.imm[21] ;
 wire \i_tinyqv.cpu.imm[22] ;
 wire \i_tinyqv.cpu.imm[23] ;
 wire \i_tinyqv.cpu.imm[24] ;
 wire \i_tinyqv.cpu.imm[25] ;
 wire \i_tinyqv.cpu.imm[26] ;
 wire \i_tinyqv.cpu.imm[27] ;
 wire \i_tinyqv.cpu.imm[28] ;
 wire \i_tinyqv.cpu.imm[29] ;
 wire \i_tinyqv.cpu.imm[30] ;
 wire \i_tinyqv.cpu.imm[31] ;
 wire \i_tinyqv.cpu.instr_data[0][0] ;
 wire \i_tinyqv.cpu.instr_data[0][10] ;
 wire \i_tinyqv.cpu.instr_data[0][11] ;
 wire \i_tinyqv.cpu.instr_data[0][12] ;
 wire \i_tinyqv.cpu.instr_data[0][13] ;
 wire \i_tinyqv.cpu.instr_data[0][14] ;
 wire \i_tinyqv.cpu.instr_data[0][15] ;
 wire \i_tinyqv.cpu.instr_data[0][1] ;
 wire \i_tinyqv.cpu.instr_data[0][2] ;
 wire \i_tinyqv.cpu.instr_data[0][3] ;
 wire \i_tinyqv.cpu.instr_data[0][4] ;
 wire \i_tinyqv.cpu.instr_data[0][5] ;
 wire \i_tinyqv.cpu.instr_data[0][6] ;
 wire \i_tinyqv.cpu.instr_data[0][7] ;
 wire \i_tinyqv.cpu.instr_data[0][8] ;
 wire \i_tinyqv.cpu.instr_data[0][9] ;
 wire \i_tinyqv.cpu.instr_data[1][0] ;
 wire \i_tinyqv.cpu.instr_data[1][10] ;
 wire \i_tinyqv.cpu.instr_data[1][11] ;
 wire \i_tinyqv.cpu.instr_data[1][12] ;
 wire \i_tinyqv.cpu.instr_data[1][13] ;
 wire \i_tinyqv.cpu.instr_data[1][14] ;
 wire \i_tinyqv.cpu.instr_data[1][15] ;
 wire \i_tinyqv.cpu.instr_data[1][1] ;
 wire \i_tinyqv.cpu.instr_data[1][2] ;
 wire \i_tinyqv.cpu.instr_data[1][3] ;
 wire \i_tinyqv.cpu.instr_data[1][4] ;
 wire \i_tinyqv.cpu.instr_data[1][5] ;
 wire \i_tinyqv.cpu.instr_data[1][6] ;
 wire \i_tinyqv.cpu.instr_data[1][7] ;
 wire \i_tinyqv.cpu.instr_data[1][8] ;
 wire \i_tinyqv.cpu.instr_data[1][9] ;
 wire \i_tinyqv.cpu.instr_data[2][0] ;
 wire \i_tinyqv.cpu.instr_data[2][10] ;
 wire \i_tinyqv.cpu.instr_data[2][11] ;
 wire \i_tinyqv.cpu.instr_data[2][12] ;
 wire \i_tinyqv.cpu.instr_data[2][13] ;
 wire \i_tinyqv.cpu.instr_data[2][14] ;
 wire \i_tinyqv.cpu.instr_data[2][15] ;
 wire \i_tinyqv.cpu.instr_data[2][1] ;
 wire \i_tinyqv.cpu.instr_data[2][2] ;
 wire \i_tinyqv.cpu.instr_data[2][3] ;
 wire \i_tinyqv.cpu.instr_data[2][4] ;
 wire \i_tinyqv.cpu.instr_data[2][5] ;
 wire \i_tinyqv.cpu.instr_data[2][6] ;
 wire \i_tinyqv.cpu.instr_data[2][7] ;
 wire \i_tinyqv.cpu.instr_data[2][8] ;
 wire \i_tinyqv.cpu.instr_data[2][9] ;
 wire \i_tinyqv.cpu.instr_data[3][0] ;
 wire \i_tinyqv.cpu.instr_data[3][10] ;
 wire \i_tinyqv.cpu.instr_data[3][11] ;
 wire \i_tinyqv.cpu.instr_data[3][12] ;
 wire \i_tinyqv.cpu.instr_data[3][13] ;
 wire \i_tinyqv.cpu.instr_data[3][14] ;
 wire \i_tinyqv.cpu.instr_data[3][15] ;
 wire \i_tinyqv.cpu.instr_data[3][1] ;
 wire \i_tinyqv.cpu.instr_data[3][2] ;
 wire \i_tinyqv.cpu.instr_data[3][3] ;
 wire \i_tinyqv.cpu.instr_data[3][4] ;
 wire \i_tinyqv.cpu.instr_data[3][5] ;
 wire \i_tinyqv.cpu.instr_data[3][6] ;
 wire \i_tinyqv.cpu.instr_data[3][7] ;
 wire \i_tinyqv.cpu.instr_data[3][8] ;
 wire \i_tinyqv.cpu.instr_data[3][9] ;
 wire \i_tinyqv.cpu.instr_data_in[0] ;
 wire \i_tinyqv.cpu.instr_data_in[10] ;
 wire \i_tinyqv.cpu.instr_data_in[11] ;
 wire \i_tinyqv.cpu.instr_data_in[12] ;
 wire \i_tinyqv.cpu.instr_data_in[13] ;
 wire \i_tinyqv.cpu.instr_data_in[14] ;
 wire \i_tinyqv.cpu.instr_data_in[15] ;
 wire \i_tinyqv.cpu.instr_data_in[1] ;
 wire \i_tinyqv.cpu.instr_data_in[2] ;
 wire \i_tinyqv.cpu.instr_data_in[3] ;
 wire \i_tinyqv.cpu.instr_data_in[4] ;
 wire \i_tinyqv.cpu.instr_data_in[5] ;
 wire \i_tinyqv.cpu.instr_data_in[6] ;
 wire \i_tinyqv.cpu.instr_data_in[7] ;
 wire \i_tinyqv.cpu.instr_data_in[8] ;
 wire \i_tinyqv.cpu.instr_data_in[9] ;
 wire \i_tinyqv.cpu.instr_data_start[10] ;
 wire \i_tinyqv.cpu.instr_data_start[11] ;
 wire \i_tinyqv.cpu.instr_data_start[12] ;
 wire \i_tinyqv.cpu.instr_data_start[13] ;
 wire \i_tinyqv.cpu.instr_data_start[14] ;
 wire \i_tinyqv.cpu.instr_data_start[15] ;
 wire \i_tinyqv.cpu.instr_data_start[16] ;
 wire \i_tinyqv.cpu.instr_data_start[17] ;
 wire \i_tinyqv.cpu.instr_data_start[18] ;
 wire \i_tinyqv.cpu.instr_data_start[19] ;
 wire \i_tinyqv.cpu.instr_data_start[20] ;
 wire \i_tinyqv.cpu.instr_data_start[21] ;
 wire \i_tinyqv.cpu.instr_data_start[22] ;
 wire \i_tinyqv.cpu.instr_data_start[23] ;
 wire \i_tinyqv.cpu.instr_data_start[3] ;
 wire \i_tinyqv.cpu.instr_data_start[4] ;
 wire \i_tinyqv.cpu.instr_data_start[5] ;
 wire \i_tinyqv.cpu.instr_data_start[6] ;
 wire \i_tinyqv.cpu.instr_data_start[7] ;
 wire \i_tinyqv.cpu.instr_data_start[8] ;
 wire \i_tinyqv.cpu.instr_data_start[9] ;
 wire \i_tinyqv.cpu.instr_fetch_running ;
 wire \i_tinyqv.cpu.instr_fetch_started ;
 wire \i_tinyqv.cpu.instr_fetch_stopped ;
 wire \i_tinyqv.cpu.instr_len[1] ;
 wire \i_tinyqv.cpu.instr_len[2] ;
 wire \i_tinyqv.cpu.instr_write_offset[1] ;
 wire \i_tinyqv.cpu.instr_write_offset[2] ;
 wire \i_tinyqv.cpu.instr_write_offset[3] ;
 wire \i_tinyqv.cpu.is_alu_imm ;
 wire \i_tinyqv.cpu.is_alu_reg ;
 wire \i_tinyqv.cpu.is_auipc ;
 wire \i_tinyqv.cpu.is_branch ;
 wire \i_tinyqv.cpu.is_jal ;
 wire \i_tinyqv.cpu.is_jalr ;
 wire \i_tinyqv.cpu.is_load ;
 wire \i_tinyqv.cpu.is_lui ;
 wire \i_tinyqv.cpu.is_store ;
 wire \i_tinyqv.cpu.is_system ;
 wire \i_tinyqv.cpu.load_started ;
 wire \i_tinyqv.cpu.mem_op_increment_reg ;
 wire \i_tinyqv.cpu.no_write_in_progress ;
 wire \i_tinyqv.cpu.pc[1] ;
 wire \i_tinyqv.cpu.pc[2] ;
 wire \i_tinyqv.cpu.was_early_branch ;
 wire \i_tinyqv.mem.data_from_read[16] ;
 wire \i_tinyqv.mem.data_from_read[17] ;
 wire \i_tinyqv.mem.data_from_read[18] ;
 wire \i_tinyqv.mem.data_from_read[19] ;
 wire \i_tinyqv.mem.data_from_read[20] ;
 wire \i_tinyqv.mem.data_from_read[21] ;
 wire \i_tinyqv.mem.data_from_read[22] ;
 wire \i_tinyqv.mem.data_from_read[23] ;
 wire \i_tinyqv.mem.data_stall ;
 wire \i_tinyqv.mem.instr_active ;
 wire \i_tinyqv.mem.q_ctrl.addr[0] ;
 wire \i_tinyqv.mem.q_ctrl.addr[10] ;
 wire \i_tinyqv.mem.q_ctrl.addr[11] ;
 wire \i_tinyqv.mem.q_ctrl.addr[12] ;
 wire \i_tinyqv.mem.q_ctrl.addr[13] ;
 wire \i_tinyqv.mem.q_ctrl.addr[14] ;
 wire \i_tinyqv.mem.q_ctrl.addr[15] ;
 wire \i_tinyqv.mem.q_ctrl.addr[16] ;
 wire \i_tinyqv.mem.q_ctrl.addr[17] ;
 wire \i_tinyqv.mem.q_ctrl.addr[18] ;
 wire \i_tinyqv.mem.q_ctrl.addr[19] ;
 wire \i_tinyqv.mem.q_ctrl.addr[1] ;
 wire \i_tinyqv.mem.q_ctrl.addr[20] ;
 wire \i_tinyqv.mem.q_ctrl.addr[21] ;
 wire \i_tinyqv.mem.q_ctrl.addr[22] ;
 wire \i_tinyqv.mem.q_ctrl.addr[23] ;
 wire \i_tinyqv.mem.q_ctrl.addr[2] ;
 wire \i_tinyqv.mem.q_ctrl.addr[3] ;
 wire \i_tinyqv.mem.q_ctrl.addr[4] ;
 wire \i_tinyqv.mem.q_ctrl.addr[5] ;
 wire \i_tinyqv.mem.q_ctrl.addr[6] ;
 wire \i_tinyqv.mem.q_ctrl.addr[7] ;
 wire \i_tinyqv.mem.q_ctrl.addr[8] ;
 wire \i_tinyqv.mem.q_ctrl.addr[9] ;
 wire \i_tinyqv.mem.q_ctrl.data_ready ;
 wire \i_tinyqv.mem.q_ctrl.data_req ;
 wire \i_tinyqv.mem.q_ctrl.delay_cycles_cfg[0] ;
 wire \i_tinyqv.mem.q_ctrl.delay_cycles_cfg[1] ;
 wire \i_tinyqv.mem.q_ctrl.delay_cycles_cfg[2] ;
 wire \i_tinyqv.mem.q_ctrl.fsm_state[0] ;
 wire \i_tinyqv.mem.q_ctrl.fsm_state[1] ;
 wire \i_tinyqv.mem.q_ctrl.fsm_state[2] ;
 wire \i_tinyqv.mem.q_ctrl.is_writing ;
 wire \i_tinyqv.mem.q_ctrl.last_ram_a_sel ;
 wire \i_tinyqv.mem.q_ctrl.last_ram_b_sel ;
 wire \i_tinyqv.mem.q_ctrl.nibbles_remaining[0] ;
 wire \i_tinyqv.mem.q_ctrl.nibbles_remaining[1] ;
 wire \i_tinyqv.mem.q_ctrl.nibbles_remaining[2] ;
 wire \i_tinyqv.mem.q_ctrl.read_cycles_count[0] ;
 wire \i_tinyqv.mem.q_ctrl.read_cycles_count[1] ;
 wire \i_tinyqv.mem.q_ctrl.read_cycles_count[2] ;
 wire \i_tinyqv.mem.q_ctrl.spi_clk_out ;
 wire \i_tinyqv.mem.q_ctrl.spi_data_oe[0] ;
 wire \i_tinyqv.mem.q_ctrl.spi_flash_select ;
 wire \i_tinyqv.mem.q_ctrl.spi_in_buffer[0] ;
 wire \i_tinyqv.mem.q_ctrl.spi_in_buffer[1] ;
 wire \i_tinyqv.mem.q_ctrl.spi_in_buffer[2] ;
 wire \i_tinyqv.mem.q_ctrl.spi_in_buffer[3] ;
 wire \i_tinyqv.mem.q_ctrl.spi_in_buffer[4] ;
 wire \i_tinyqv.mem.q_ctrl.spi_in_buffer[5] ;
 wire \i_tinyqv.mem.q_ctrl.spi_in_buffer[6] ;
 wire \i_tinyqv.mem.q_ctrl.spi_in_buffer[7] ;
 wire \i_tinyqv.mem.q_ctrl.spi_ram_a_select ;
 wire \i_tinyqv.mem.q_ctrl.spi_ram_b_select ;
 wire \i_tinyqv.mem.q_ctrl.stop_txn_reg ;
 wire \i_tinyqv.mem.qspi_data_buf[10] ;
 wire \i_tinyqv.mem.qspi_data_buf[11] ;
 wire \i_tinyqv.mem.qspi_data_buf[12] ;
 wire \i_tinyqv.mem.qspi_data_buf[13] ;
 wire \i_tinyqv.mem.qspi_data_buf[14] ;
 wire \i_tinyqv.mem.qspi_data_buf[15] ;
 wire \i_tinyqv.mem.qspi_data_buf[24] ;
 wire \i_tinyqv.mem.qspi_data_buf[25] ;
 wire \i_tinyqv.mem.qspi_data_buf[26] ;
 wire \i_tinyqv.mem.qspi_data_buf[27] ;
 wire \i_tinyqv.mem.qspi_data_buf[28] ;
 wire \i_tinyqv.mem.qspi_data_buf[29] ;
 wire \i_tinyqv.mem.qspi_data_buf[30] ;
 wire \i_tinyqv.mem.qspi_data_buf[31] ;
 wire \i_tinyqv.mem.qspi_data_buf[8] ;
 wire \i_tinyqv.mem.qspi_data_buf[9] ;
 wire \i_tinyqv.mem.qspi_data_byte_idx[0] ;
 wire \i_tinyqv.mem.qspi_data_byte_idx[1] ;
 wire \i_tinyqv.mem.qspi_write_done ;
 wire \i_uart_rx.bit_sample ;
 wire \i_uart_rx.cycle_counter[0] ;
 wire \i_uart_rx.cycle_counter[10] ;
 wire \i_uart_rx.cycle_counter[1] ;
 wire \i_uart_rx.cycle_counter[2] ;
 wire \i_uart_rx.cycle_counter[3] ;
 wire \i_uart_rx.cycle_counter[4] ;
 wire \i_uart_rx.cycle_counter[5] ;
 wire \i_uart_rx.cycle_counter[6] ;
 wire \i_uart_rx.cycle_counter[7] ;
 wire \i_uart_rx.cycle_counter[8] ;
 wire \i_uart_rx.cycle_counter[9] ;
 wire \i_uart_rx.fsm_state[0] ;
 wire \i_uart_rx.fsm_state[1] ;
 wire \i_uart_rx.fsm_state[2] ;
 wire \i_uart_rx.fsm_state[3] ;
 wire \i_uart_rx.recieved_data[0] ;
 wire \i_uart_rx.recieved_data[1] ;
 wire \i_uart_rx.recieved_data[2] ;
 wire \i_uart_rx.recieved_data[3] ;
 wire \i_uart_rx.recieved_data[4] ;
 wire \i_uart_rx.recieved_data[5] ;
 wire \i_uart_rx.recieved_data[6] ;
 wire \i_uart_rx.recieved_data[7] ;
 wire \i_uart_rx.rxd_reg[0] ;
 wire \i_uart_rx.rxd_reg[1] ;
 wire \i_uart_rx.uart_rts ;
 wire \i_uart_tx.cycle_counter[0] ;
 wire \i_uart_tx.cycle_counter[10] ;
 wire \i_uart_tx.cycle_counter[1] ;
 wire \i_uart_tx.cycle_counter[2] ;
 wire \i_uart_tx.cycle_counter[3] ;
 wire \i_uart_tx.cycle_counter[4] ;
 wire \i_uart_tx.cycle_counter[5] ;
 wire \i_uart_tx.cycle_counter[6] ;
 wire \i_uart_tx.cycle_counter[7] ;
 wire \i_uart_tx.cycle_counter[8] ;
 wire \i_uart_tx.cycle_counter[9] ;
 wire \i_uart_tx.data_to_send[0] ;
 wire \i_uart_tx.data_to_send[1] ;
 wire \i_uart_tx.data_to_send[2] ;
 wire \i_uart_tx.data_to_send[3] ;
 wire \i_uart_tx.data_to_send[4] ;
 wire \i_uart_tx.data_to_send[5] ;
 wire \i_uart_tx.data_to_send[6] ;
 wire \i_uart_tx.data_to_send[7] ;
 wire \i_uart_tx.fsm_state[0] ;
 wire \i_uart_tx.fsm_state[1] ;
 wire \i_uart_tx.fsm_state[2] ;
 wire \i_uart_tx.fsm_state[3] ;
 wire \i_uart_tx.txd_reg ;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net29;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net3;
 wire net30;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net31;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net32;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net4;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net5;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net6;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;

 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(_0865_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(_3068_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(\i_tinyqv.cpu.data_addr[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(\i_tinyqv.cpu.i_core.imm_lo[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_13 (.DIODE(\i_tinyqv.cpu.i_core.imm_lo[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_14 (.DIODE(\i_tinyqv.cpu.i_core.mepc[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_15 (.DIODE(\i_tinyqv.cpu.imm[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_16 (.DIODE(\i_tinyqv.cpu.imm[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_17 (.DIODE(\i_tinyqv.cpu.imm[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_18 (.DIODE(\i_tinyqv.mem.q_ctrl.addr[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_19 (.DIODE(\i_tinyqv.mem.q_ctrl.addr[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(_0991_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_20 (.DIODE(\i_tinyqv.mem.q_ctrl.addr[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_21 (.DIODE(\i_tinyqv.mem.q_ctrl.addr[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_22 (.DIODE(\i_tinyqv.mem.q_ctrl.addr[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_23 (.DIODE(\i_tinyqv.mem.q_ctrl.addr[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_24 (.DIODE(\i_uart_rx.recieved_data[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_25 (.DIODE(net69),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_26 (.DIODE(_1302_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_27 (.DIODE(_3010_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_28 (.DIODE(\i_debug_uart_tx.uart_tx_data[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_29 (.DIODE(\i_tinyqv.cpu.i_core.i_registers.registers[6][3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(_1054_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_30 (.DIODE(\i_tinyqv.cpu.i_core.imm_lo[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_31 (.DIODE(\i_tinyqv.cpu.i_core.imm_lo[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_32 (.DIODE(\i_tinyqv.cpu.i_core.is_interrupt ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_33 (.DIODE(\i_tinyqv.cpu.i_core.mepc[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_34 (.DIODE(\i_tinyqv.cpu.i_core.imm_lo[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_35 (.DIODE(\i_tinyqv.cpu.i_core.imm_lo[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_36 (.DIODE(\i_tinyqv.cpu.i_core.imm_lo[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_37 (.DIODE(\i_tinyqv.cpu.i_core.imm_lo[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_38 (.DIODE(\i_tinyqv.cpu.i_core.imm_lo[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_39 (.DIODE(\i_tinyqv.cpu.i_core.imm_lo[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(_1185_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_40 (.DIODE(\i_tinyqv.cpu.i_core.imm_lo[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_41 (.DIODE(\i_tinyqv.cpu.i_core.imm_lo[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_42 (.DIODE(\i_tinyqv.cpu.i_core.imm_lo[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_43 (.DIODE(\i_tinyqv.cpu.i_core.imm_lo[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_44 (.DIODE(\i_tinyqv.cpu.i_core.imm_lo[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_45 (.DIODE(\i_tinyqv.cpu.i_core.imm_lo[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_46 (.DIODE(\i_tinyqv.cpu.i_core.imm_lo[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_47 (.DIODE(\i_tinyqv.cpu.i_core.imm_lo[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_48 (.DIODE(\i_tinyqv.cpu.i_core.imm_lo[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(_1729_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(_2507_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(_2734_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(_2930_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(_2938_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_129 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_15 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_0_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_0_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_177 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_0_186 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_0_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_0_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_0_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_0_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_0_331 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_335 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_337 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_0_365 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_369 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_0_386 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_401 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_41 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_421 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_473 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_501 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_0_521 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_529 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_533 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_545 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_557 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_561 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_573 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_585 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_589 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_601 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_613 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_617 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_629 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_641 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_645 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_657 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_669 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_673 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_685 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_69 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_697 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_701 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_0_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_103 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_10_112 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_10_193 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_10_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_201 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_234 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_10_246 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_10_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_10_273 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_10_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_10_301 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_309 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_10_321 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_33 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_10_345 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_10_368 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_10_395 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_403 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_10_413 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_419 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_10_421 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_10_464 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_475 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_50 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_10_525 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_531 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_10_533 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_10_554 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_10_561 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_10_580 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_586 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_10_589 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_10_603 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_10_618 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_10_625 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_643 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_645 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_10_660 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_664 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_10_676 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_687 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_10_693 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_10_710 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_10_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_10_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_11_106 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_11_121 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_11_135 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_11_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_11_209 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_215 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_229 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_271 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_11_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_285 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_11_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_11_326 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_11_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_11_370 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_11_382 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_11_441 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_447 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_11_449 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_11_468 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_11_482 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_11_498 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_11_505 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_11_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_11_543 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_11_550 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_559 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_564 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_11_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_576 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_11_592 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_11_605 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_11_613 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_11_627 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_638 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_11_653 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_11_662 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_11_670 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_11_673 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_677 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_11_68 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_682 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_696 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_12_136 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_12_157 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_12_193 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_209 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_226 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_12_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_12_296 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_12_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_313 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_12_344 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_12_413 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_419 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_421 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_430 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_456 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_474 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_477 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_12_518 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_12_533 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_541 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_12_556 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_12_581 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_587 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_602 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_12_614 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_632 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_643 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_650 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_656 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_12_664 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_670 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_12_690 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_698 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_701 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_12_78 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_12_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_13_107 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_13_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_117 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_13_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_151 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_13_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_13_183 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_13_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_201 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_13_210 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_214 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_13_241 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_245 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_13_254 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_13_275 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_13_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_13_305 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_13_325 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_13_353 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_13_367 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_371 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_13_380 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_13_393 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_13_415 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_13_442 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_13_46 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_13_465 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_13_476 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_13_490 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_13_505 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_13_543 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_13_553 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_559 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_13_561 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_13_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_570 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_13_582 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_590 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_13_605 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_61 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_615 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_13_627 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_13_635 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_13_645 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_13_658 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_664 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_13_670 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_13_676 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_13_683 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_13_691 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_13_70 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_13_710 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_13_95 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_14_101 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_14_121 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_14_136 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_14_160 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_14_171 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_14_191 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_213 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_14_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_230 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_14_247 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_14_269 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_273 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_14_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_14_297 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_14_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_14_317 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_14_359 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_363 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_14_417 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_14_437 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_475 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_14_525 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_531 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_14_533 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_537 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_545 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_14_561 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_569 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_573 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_587 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_14_589 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_597 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_14_601 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_605 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_14_625 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_14_633 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_14_639 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_643 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_14_645 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_651 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_655 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_14_667 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_673 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_681 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_14_689 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_14_697 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_14_711 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_14_80 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_102 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_15_12 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_130 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_147 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_164 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_18 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_185 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_15_202 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_27 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_326 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_335 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_15_337 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_15_364 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_376 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_15_388 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_15_425 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_429 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_438 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_15_449 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_455 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_15_48 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_15_480 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_15_499 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_503 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_15_505 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_15_520 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_15_536 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_15_546 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_15_556 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_15_564 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_15_572 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_15_587 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_15_595 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_608 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_624 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_15_643 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_65 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_671 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_15_691 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_101 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_16_118 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_126 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_16_136 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_178 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_206 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_224 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_16_242 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_16_261 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_16_272 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_285 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_16_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_316 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_16_360 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_16_365 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_369 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_16_37 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_16_386 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_394 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_419 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_429 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_16_471 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_475 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_16_501 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_505 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_16_528 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_539 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_16_551 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_555 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_575 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_16_58 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_587 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_16_614 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_618 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_625 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_16_633 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_637 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_64 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_16_641 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_648 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_665 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_16_686 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_699 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_16_707 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_16_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_17_107 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_148 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_17_165 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_187 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_191 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_218 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_17_259 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_265 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_272 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_17_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_17_294 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_17_313 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_17_332 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_351 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_17_369 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_393 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_17_403 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_43 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_17_438 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_446 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_457 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_17_498 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_17_519 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_527 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_17_536 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_17_551 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_559 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_17_568 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_17_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_17_576 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_591 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_17_609 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_615 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_17_633 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_641 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_658 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_670 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_17_690 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_17_708 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_712 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_79 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_17_96 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_18_160 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_188 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_18_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_239 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_18_273 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_277 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_18_288 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_18_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_294 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_18_298 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_306 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_18_318 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_329 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_354 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_18_389 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_397 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_18_414 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_18_429 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_18_472 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_493 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_519 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_554 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_18_578 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_18_599 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_603 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_642 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_18_656 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_18_689 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_693 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_711 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_19_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_19_121 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_19_186 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_190 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_215 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_19_277 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_19_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_19_298 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_19_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_304 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_327 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_335 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_19_337 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_19_357 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_19_364 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_19_404 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_19_434 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_19_457 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_19_466 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_470 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_19_474 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_19_49 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_19_500 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_549 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_19_561 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_572 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_19_586 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_19_601 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_19_613 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_19_617 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_19_640 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_19_648 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_19_659 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_19_667 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_673 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_19_679 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_687 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_19_691 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_19_703 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_19_711 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_19_89 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_1_121 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_142 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_151 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_1_177 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_1_198 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_1_220 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_1_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_1_245 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_297 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_1_322 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_1_361 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_1_373 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_39 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_1_441 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_447 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_1_481 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_487 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_529 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_541 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_1_553 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_559 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_561 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_1_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_573 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_585 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_597 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_1_609 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_615 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_617 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_629 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_641 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_653 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_1_665 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_671 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_673 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_685 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_697 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_1_709 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_1_71 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_87 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_20_157 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_161 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_164 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_20_177 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_269 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_292 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_328 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_20_345 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_20_365 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_377 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_418 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_20_421 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_20_437 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_441 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_474 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_20_485 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_493 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_20_523 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_531 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_20_560 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_20_579 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_587 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_589 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_594 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_606 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_611 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_626 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_20_639 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_643 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_20_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_663 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_20_684 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_20_692 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_20_709 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_20_79 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_20_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_89 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_21_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_21_161 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_21_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_21_179 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_21_189 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_21_207 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_21_277 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_286 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_21_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_21_304 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_310 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_21_321 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_325 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_21_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_371 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_21_384 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_21_401 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_444 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_21_449 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_453 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_21_500 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_21_534 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_538 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_21_555 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_21_577 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_21_604 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_615 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_21_643 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_651 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_21_659 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_667 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_671 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_21_680 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_21_711 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_21_90 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_22_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_22_152 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_188 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_213 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_22_231 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_248 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_269 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_280 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_22_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_22_299 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_22_343 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_347 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_22_365 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_373 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_22_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_22_415 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_419 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_22_421 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_427 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_47 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_480 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_22_529 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_22_533 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_541 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_22_561 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_22_585 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_616 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_624 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_642 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_22_645 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_657 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_22_675 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_695 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_22_710 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_22_72 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_23_108 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_23_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_23_159 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_23_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_175 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_19 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_23_219 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_23_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_23_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_23_277 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_23_31 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_23_316 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_320 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_325 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_346 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_23_387 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_391 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_393 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_23_442 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_23_468 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_23_49 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_23_495 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_23_508 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_23_536 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_23_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_23_588 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_23_596 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_63 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_643 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_23_670 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_694 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_712 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_23_96 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_24_101 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_24_122 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_126 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_136 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_24_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_24_159 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_24_189 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_24_210 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_24_246 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_24_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_272 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_24_294 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_24_302 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_24_312 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_24_330 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_24_365 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_369 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_24_37 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_24_390 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_394 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_24_411 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_419 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_24_421 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_24_432 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_438 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_24_509 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_517 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_24_522 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_24_530 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_545 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_553 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_24_560 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_24_573 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_24_586 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_24_614 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_24_66 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_24_710 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_72 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_24_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_25_108 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_25_129 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_25_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_25_220 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_25_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_25_257 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_25_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_326 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_353 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_365 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_409 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_426 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_25_443 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_447 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_449 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_25_459 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_25_485 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_530 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_545 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_25_557 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_25_600 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_25_612 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_617 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_671 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_25_691 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_711 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_98 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_26_101 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_26_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_26_157 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_163 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_219 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_230 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_276 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_26_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_26_312 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_318 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_33 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_345 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_362 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_380 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_418 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_26_42 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_26_424 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_26_448 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_474 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_26_50 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_26_509 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_517 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_26_522 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_530 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_26_540 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_554 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_578 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_26_589 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_639 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_65 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_657 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_26_695 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_699 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_26_710 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_26_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_27_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_27_12 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_129 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_27_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_27_149 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_27_178 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_18 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_27_196 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_27_206 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_27_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_273 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_27_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_313 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_27_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_27_365 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_27_396 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_404 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_422 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_447 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_27_468 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_27_484 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_27_498 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_27_529 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_27_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_27_542 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_550 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_27_570 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_574 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_27_587 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_27_599 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_603 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_27_613 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_27_617 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_671 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_27_673 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_712 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_73 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_27_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_130 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_28_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_28_175 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_179 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_28_216 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_28_234 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_28_25 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_28_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_28_313 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_319 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_28_343 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_28_397 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_28_405 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_28_412 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_416 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_28_421 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_28_429 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_28_445 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_28_45 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_28_452 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_458 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_28_490 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_498 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_28_515 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_28_520 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_28_538 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_572 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_28_607 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_699 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_71 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_28_710 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_28_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_89 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_29_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_178 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_29_190 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_29_204 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_29_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_29_228 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_232 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_252 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_29_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_29_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_29_300 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_319 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_337 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_29_357 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_391 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_409 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_29_414 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_29_441 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_447 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_29_464 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_485 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_29_499 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_503 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_29_505 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_509 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_29_517 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_525 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_533 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_29_545 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_559 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_29_567 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_29_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_586 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_596 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_29_608 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_29_614 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_617 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_624 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_29_629 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_29_641 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_29_656 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_29_668 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_29_673 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_29_91 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_2_101 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_123 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_2_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_2_160 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_164 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_2_189 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_2_233 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_2_261 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_2_293 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_299 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_2_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_2_344 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_2_381 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_403 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_2_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_2_421 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_443 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_2_452 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_456 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_47 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_2_473 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_2_525 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_531 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_533 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_545 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_557 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_2_56 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_569 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_2_581 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_587 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_589 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_601 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_613 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_625 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_2_637 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_64 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_643 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_645 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_657 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_669 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_681 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_2_693 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_699 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_701 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_2_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_30_101 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_30_120 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_126 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_30_135 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_30_188 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_30_226 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_245 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_256 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_266 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_30_283 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_30_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_303 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_337 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_341 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_30_349 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_369 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_30_390 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_418 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_30_421 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_30_432 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_440 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_449 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_465 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_474 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_483 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_30_499 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_503 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_520 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_531 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_30_541 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_545 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_557 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_30_563 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_30_584 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_30_589 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_30_60 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_611 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_30_640 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_699 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_30_710 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_30_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_103 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_129 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_31_146 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_31_177 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_31_202 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_207 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_31_218 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_31_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_31_268 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_31_357 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_362 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_38 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_31_389 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_31_445 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_449 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_31_465 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_471 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_31_496 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_503 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_505 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_31_512 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_524 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_31_534 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_31_556 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_561 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_606 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_31_617 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_635 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_31_646 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_31_668 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_31_691 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_74 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_31_99 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_32_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_32_13 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_32_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_32_149 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_32_168 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_172 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_32_189 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_32_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_32_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_32_229 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_32_248 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_32_270 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_32_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_325 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_32_349 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_32_362 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_32_395 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_32_403 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_412 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_32_418 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_32_42 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_32_431 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_32_436 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_32_448 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_456 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_32_460 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_32_468 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_32_474 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_482 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_32_496 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_50 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_32_520 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_531 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_32_539 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_553 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_573 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_32_580 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_584 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_32_589 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_32_636 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_32_67 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_699 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_32_710 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_32_78 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_101 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_33_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_33_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_117 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_33_158 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_33_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_33_174 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_33_200 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_33_206 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_33_218 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_33_260 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_284 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_293 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_33_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_308 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_318 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_33_337 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_33_357 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_33_364 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_33_426 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_442 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_33_454 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_33_471 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_475 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_33_502 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_33_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_33_542 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_551 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_559 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_33_567 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_33_582 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_33_601 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_33_612 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_617 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_33_627 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_33_640 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_671 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_33_682 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_686 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_33_696 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_702 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_33_709 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_33_73 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_33_95 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_34_120 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_34_132 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_34_144 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_151 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_34_160 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_178 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_34_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_34_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_34_205 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_34_217 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_221 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_34_231 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_275 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_34_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_322 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_34_336 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_342 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_360 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_34_365 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_34_373 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_383 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_34_393 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_34_402 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_406 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_34_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_34_428 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_34_438 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_34_446 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_34_454 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_475 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_34_477 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_49 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_34_530 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_34_542 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_546 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_34_563 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_34_572 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_34_58 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_34_583 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_587 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_595 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_34_626 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_632 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_34_642 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_34_66 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_34_663 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_683 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_34_710 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_34_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_35_100 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_35_121 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_132 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_156 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_35_163 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_35_175 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_179 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_185 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_35_192 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_198 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_35_206 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_35_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_243 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_278 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_305 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_318 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_358 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_371 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_35_445 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_35_458 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_35_491 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_503 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_35_52 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_35_547 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_559 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_35_561 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_35_576 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_35_583 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_35_603 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_615 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_617 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_35_640 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_673 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_35_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_36_14 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_36_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_36_149 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_36_154 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_36_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_36_227 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_36_239 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_36_248 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_36_25 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_36_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_36_265 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_36_288 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_36_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_36_306 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_346 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_360 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_372 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_36_38 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_36_416 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_42 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_36_421 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_427 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_36_464 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_36_485 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_36_507 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_36_530 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_36_539 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_547 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_36_560 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_566 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_36_589 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_601 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_36_605 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_36_616 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_643 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_36_645 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_36_657 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_36_698 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_36_710 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_37_107 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_37_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_37_12 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_135 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_37_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_180 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_37_203 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_37_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_231 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_37_240 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_254 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_272 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_278 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_37_287 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_37_299 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_37_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_37_313 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_324 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_34 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_359 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_363 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_381 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_37_393 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_37_405 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_37_414 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_418 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_37_437 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_37_445 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_37_464 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_468 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_474 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_489 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_37_500 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_505 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_37_524 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_559 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_561 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_582 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_37_586 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_651 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_37_665 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_671 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_37_673 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_677 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_38_106 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_118 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_38_135 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_161 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_168 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_178 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_183 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_191 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_38_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_218 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_38_247 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_38_25 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_38_261 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_38_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_38_299 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_344 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_363 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_38_378 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_382 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_38_394 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_418 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_38_421 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_425 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_38_442 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_460 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_470 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_38_505 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_518 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_530 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_38_566 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_578 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_60 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_38_686 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_38_694 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_38_710 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_79 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_96 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_39_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_39_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_39_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_39_157 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_39_183 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_39_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_39_202 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_39_219 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_39_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_39_231 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_39_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_39_259 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_39_28 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_39_287 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_39_325 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_39_337 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_39_370 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_39_378 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_39_384 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_39_401 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_39_430 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_39_465 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_39_482 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_39_494 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_39_50 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_39_503 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_39_533 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_39_558 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_39_588 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_39_597 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_39_617 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_39_625 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_39_63 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_39_670 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_39_689 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_39_693 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_3_107 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_3_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_3_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_3_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_3_213 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_3_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_257 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_3_274 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_3_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_285 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_337 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_347 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_3_365 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_3_385 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_391 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_3_425 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_431 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_3_45 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_3_481 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_487 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_505 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_539 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_3_551 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_559 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_561 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_573 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_585 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_597 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_3_609 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_615 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_624 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_636 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_648 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_660 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_673 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_685 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_697 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_3_709 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_3_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_89 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_40_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_40_119 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_40_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_40_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_40_189 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_40_202 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_40_215 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_40_237 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_40_246 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_40_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_40_261 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_40_272 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_40_306 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_40_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_40_313 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_40_32 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_40_344 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_40_362 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_40_365 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_40_38 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_40_386 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_40_396 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_40_411 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_40_421 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_40_429 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_40_447 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_40_462 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_40_474 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_40_486 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_40_525 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_40_531 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_40_533 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_40_539 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_40_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_40_583 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_40_587 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_40_605 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_40_643 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_40_679 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_40_689 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_40_699 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_40_710 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_40_80 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_40_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_40_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_41_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_41_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_41_159 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_41_190 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_41_20 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_41_218 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_41_255 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_41_264 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_41_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_41_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_41_310 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_41_337 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_41_400 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_41_406 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_41_424 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_41_430 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_41_438 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_41_446 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_41_457 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_41_46 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_41_474 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_41_485 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_41_501 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_41_519 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_41_526 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_41_544 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_41_557 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_41_570 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_41_581 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_41_591 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_41_607 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_41_615 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_41_617 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_41_621 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_41_652 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_41_670 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_41_76 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_42_107 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_42_115 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_42_136 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_42_149 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_42_159 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_42_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_42_177 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_42_183 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_42_190 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_42_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_42_20 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_42_202 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_42_206 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_42_214 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_42_218 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_42_24 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_42_241 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_42_256 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_42_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_42_323 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_42_337 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_42_362 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_42_365 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_42_375 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_42_388 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_42_404 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_42_416 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_42_421 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_42_441 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_42_470 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_42_493 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_42_502 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_42_506 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_42_514 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_42_530 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_42_533 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_42_563 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_42_587 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_42_589 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_42_609 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_42_61 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_42_624 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_42_642 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_42_654 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_42_665 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_42_679 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_42_710 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_42_80 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_43_102 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_43_118 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_43_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_43_145 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_43_152 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_43_163 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_43_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_43_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_43_180 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_43_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_43_207 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_43_217 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_43_222 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_43_235 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_43_248 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_43_252 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_43_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_43_287 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_43_291 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_43_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_43_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_43_344 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_43_349 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_43_355 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_43_369 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_43_375 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_43_409 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_43_429 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_43_434 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_43_441 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_43_449 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_43_477 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_43_494 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_43_502 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_43_512 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_43_521 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_43_527 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_43_536 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_43_558 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_43_570 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_43_574 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_43_578 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_43_595 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_43_614 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_43_664 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_43_682 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_43_711 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_43_76 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_44_122 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_44_126 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_44_134 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_44_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_44_174 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_44_186 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_44_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_44_190 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_44_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_44_201 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_44_207 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_44_234 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_44_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_44_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_44_298 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_44_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_44_317 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_44_332 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_44_358 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_44_392 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_44_406 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_44_418 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_44_421 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_44_449 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_44_453 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_44_515 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_44_549 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_44_568 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_44_587 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_44_600 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_44_61 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_44_632 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_44_642 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_44_648 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_44_689 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_44_79 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_44_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_44_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_45_101 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_45_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_45_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_45_117 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_45_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_45_154 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_45_165 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_45_175 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_45_180 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_45_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_45_221 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_45_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_45_232 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_45_255 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_45_268 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_45_278 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_45_28 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_45_294 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_45_324 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_45_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_45_34 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_45_343 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_45_393 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_45_408 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_45_443 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_45_447 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_45_455 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_45_462 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_45_474 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_45_488 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_45_500 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_45_513 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_45_52 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_45_528 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_45_532 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_45_561 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_45_570 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_45_604 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_45_612 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_45_617 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_45_654 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_45_66 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_45_671 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_45_673 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_45_693 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_45_80 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_46_121 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_46_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_46_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_46_147 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_46_158 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_46_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_46_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_46_234 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_46_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_46_258 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_46_264 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_46_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_46_288 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_46_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_46_306 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_46_32 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_46_372 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_46_388 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_46_401 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_46_406 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_46_416 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_46_430 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_46_449 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_46_462 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_46_470 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_46_474 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_46_477 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_46_503 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_46_521 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_46_533 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_46_552 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_46_564 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_46_587 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_46_592 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_46_602 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_46_614 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_46_631 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_46_654 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_46_672 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_46_676 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_46_698 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_46_710 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_46_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_46_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_47_103 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_47_119 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_47_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_47_146 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_47_163 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_47_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_47_177 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_47_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_47_192 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_47_210 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_47_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_47_236 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_47_25 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_47_261 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_47_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_47_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_47_305 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_47_325 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_47_353 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_47_365 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_47_385 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_47_389 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_47_409 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_47_42 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_47_436 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_47_447 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_47_453 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_47_491 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_47_503 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_47_529 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_47_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_47_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_47_584 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_47_601 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_47_612 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_47_617 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_47_643 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_47_676 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_47_701 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_47_74 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_47_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_48_104 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_48_118 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_48_144 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_48_155 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_48_182 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_48_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_48_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_48_224 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_48_249 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_48_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_48_257 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_48_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_48_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_48_296 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_48_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_48_330 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_48_363 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_48_368 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_48_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_48_392 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_48_397 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_48_415 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_48_433 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_48_464 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_48_472 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_48_481 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_48_498 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_48_516 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_48_524 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_48_541 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_48_553 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_48_587 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_48_603 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_48_613 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_48_617 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_48_627 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_48_63 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_48_639 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_48_643 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_48_653 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_48_663 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_48_689 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_48_695 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_48_699 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_48_701 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_48_75 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_48_94 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_49_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_49_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_49_159 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_49_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_49_185 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_49_192 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_49_209 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_49_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_49_240 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_49_257 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_49_275 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_49_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_49_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_49_285 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_49_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_49_302 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_49_306 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_49_329 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_49_359 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_49_37 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_49_377 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_49_391 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_49_405 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_49_441 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_49_446 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_49_449 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_49_480 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_49_493 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_49_501 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_49_511 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_49_528 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_49_532 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_49_552 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_49_569 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_49_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_49_577 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_49_583 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_49_597 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_49_605 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_49_611 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_49_615 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_49_623 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_49_629 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_49_635 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_49_647 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_49_651 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_49_660 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_49_673 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_49_683 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_49_687 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_49_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_49_95 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_4_108 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_4_136 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_4_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_4_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_157 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_4_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_4_249 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_288 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_4_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_298 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_4_325 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_33 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_4_357 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_363 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_381 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_4_415 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_419 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_437 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_4_471 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_475 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_4_485 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_50 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_4_529 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_549 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_561 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_4_573 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_605 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_4_626 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_4_634 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_642 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_4_645 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_4_655 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_663 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_673 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_685 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_4_697 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_701 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_4_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_50_101 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_50_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_50_121 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_50_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_50_156 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_50_168 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_50_172 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_50_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_50_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_50_220 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_50_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_50_257 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_50_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_50_298 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_50_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_50_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_50_336 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_50_354 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_50_373 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_50_377 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_50_381 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_50_396 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_50_403 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_50_437 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_50_446 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_50_456 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_50_472 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_50_506 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_50_510 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_50_518 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_50_528 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_50_533 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_50_587 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_50_589 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_50_611 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_50_62 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_50_627 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_50_653 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_50_668 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_50_695 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_50_704 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_50_712 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_50_76 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_50_80 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_50_94 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_51_122 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_51_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_51_162 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_51_191 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_51_206 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_51_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_51_231 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_51_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_51_254 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_51_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_51_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_51_300 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_51_350 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_51_368 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_51_38 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_51_387 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_51_414 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_51_422 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_51_449 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_51_471 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_51_483 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_51_489 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_51_505 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_51_509 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_51_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_51_529 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_51_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_51_556 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_51_567 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_51_578 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_51_586 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_51_596 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_51_605 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_51_613 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_51_617 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_51_629 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_51_634 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_51_642 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_51_649 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_51_673 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_51_685 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_51_711 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_51_76 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_52_112 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_52_131 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_52_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_52_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_52_200 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_52_231 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_52_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_52_288 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_52_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_52_312 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_52_379 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_52_390 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_52_394 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_52_398 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_52_419 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_52_430 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_52_440 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_52_444 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_52_464 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_52_475 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_52_493 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_52_499 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_52_508 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_52_512 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_52_540 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_52_548 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_52_558 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_52_586 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_52_589 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_52_600 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_52_609 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_52_618 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_52_628 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_52_655 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_52_689 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_52_697 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_52_710 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_52_74 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_52_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_52_94 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_53_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_53_121 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_53_186 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_53_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_53_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_53_236 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_53_244 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_53_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_53_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_53_351 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_53_358 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_53_384 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_53_388 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_53_399 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_53_416 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_53_434 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_53_447 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_53_476 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_53_482 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_53_500 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_53_521 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_53_531 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_53_545 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_53_559 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_53_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_53_586 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_53_611 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_53_615 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_53_617 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_53_625 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_53_637 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_53_648 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_53_669 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_53_711 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_53_78 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_53_84 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_53_94 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_54_121 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_54_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_54_148 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_54_168 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_54_190 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_54_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_54_214 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_54_241 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_54_269 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_54_282 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_54_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_54_381 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_54_418 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_54_469 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_54_477 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_54_492 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_54_533 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_54_551 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_54_559 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_54_569 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_54_581 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_54_587 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_54_589 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_54_593 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_54_605 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_54_629 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_54_635 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_54_642 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_54_651 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_54_665 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_54_669 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_54_686 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_54_690 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_54_698 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_54_704 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_54_712 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_54_78 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_55_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_55_159 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_55_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_55_202 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_55_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_55_234 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_55_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_55_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_55_322 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_55_340 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_55_367 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_55_371 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_55_379 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_55_402 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_55_406 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_55_439 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_55_447 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_55_461 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_55_469 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_55_475 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_55_491 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_55_499 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_55_514 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_55_527 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_55_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_55_558 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_55_561 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_55_593 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_55_597 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_55_610 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_55_620 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_55_631 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_55_639 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_55_643 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_55_651 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_55_658 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_55_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_55_75 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_55_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_56_157 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_56_177 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_56_190 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_56_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_56_217 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_56_269 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_56_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_56_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_56_345 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_56_362 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_56_38 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_56_382 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_56_386 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_56_397 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_56_416 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_56_421 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_56_427 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_56_444 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_56_496 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_56_507 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_56_525 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_56_544 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_56_551 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_56_571 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_56_579 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_56_583 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_56_587 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_56_611 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_56_653 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_56_712 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_56_94 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_57_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_57_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_57_130 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_57_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_57_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_57_221 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_57_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_57_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_57_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_57_304 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_57_311 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_57_324 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_57_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_57_337 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_57_34 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_57_347 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_57_359 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_57_402 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_57_417 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_57_421 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_57_426 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_57_438 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_57_446 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_57_461 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_57_467 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_57_492 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_57_513 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_57_519 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_57_523 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_57_533 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_57_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_57_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_57_584 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_57_594 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_57_605 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_57_613 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_57_62 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_57_631 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_57_640 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_57_647 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_57_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_57_92 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_58_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_58_114 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_58_118 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_58_172 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_58_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_58_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_58_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_58_216 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_58_232 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_58_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_58_256 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_58_274 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_58_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_58_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_58_318 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_58_356 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_58_379 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_58_38 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_58_385 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_58_396 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_58_421 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_58_425 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_58_441 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_58_445 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_58_474 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_58_484 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_58_494 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_58_502 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_58_510 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_58_530 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_58_533 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_58_537 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_58_546 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_58_572 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_58_583 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_58_587 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_58_604 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_58_612 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_58_637 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_58_643 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_58_645 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_58_664 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_58_710 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_58_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_58_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_59_149 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_59_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_59_186 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_59_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_59_270 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_59_287 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_59_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_59_337 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_59_348 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_59_355 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_59_366 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_59_393 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_59_403 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_59_424 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_59_428 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_59_446 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_59_449 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_59_469 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_59_482 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_59_512 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_59_541 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_59_561 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_59_565 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_59_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_59_575 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_59_590 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_59_600 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_59_614 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_59_661 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_59_689 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_59_70 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_59_712 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_59_94 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_103 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_5_121 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_5_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_5_191 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_5_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_236 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_5_249 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_5_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_5_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_5_330 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_337 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_354 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_376 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_5_388 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_5_393 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_401 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_5_419 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_5_445 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_5_449 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_5_460 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_464 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_5_481 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_487 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_5_513 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_5_52 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_533 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_559 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_5_561 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_573 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_585 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_598 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_5_610 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_625 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_635 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_659 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_681 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_693 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_5_705 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_5_99 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_60_114 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_60_150 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_60_184 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_60_221 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_60_24 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_60_268 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_60_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_60_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_60_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_60_359 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_60_365 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_60_382 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_60_394 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_60_399 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_60_409 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_60_419 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_60_427 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_60_436 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_60_449 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_60_458 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_60_47 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_60_474 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_60_480 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_60_501 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_60_510 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_60_518 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_60_522 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_60_538 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_60_566 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_60_580 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_60_615 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_60_623 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_60_639 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_60_661 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_60_699 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_60_712 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_60_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_60_94 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_61_100 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_61_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_61_117 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_61_130 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_61_152 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_61_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_61_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_61_192 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_61_210 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_61_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_61_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_61_235 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_61_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_61_293 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_61_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_61_312 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_61_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_61_345 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_61_356 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_61_362 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_61_372 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_61_400 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_61_418 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_61_440 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_61_472 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_61_481 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_61_503 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_61_540 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_61_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_61_559 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_61_561 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_61_599 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_61_640 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_61_655 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_61_673 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_61_677 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_61_686 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_61_712 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_62_115 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_62_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_62_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_62_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_62_152 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_62_20 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_62_217 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_62_226 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_62_230 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_62_24 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_62_241 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_62_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_62_270 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_62_317 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_62_321 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_62_363 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_62_414 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_62_425 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_62_449 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_62_45 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_62_455 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_62_469 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_62_475 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_62_485 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_62_505 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_62_514 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_62_520 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_62_542 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_62_557 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_62_589 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_62_63 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_62_712 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_62_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_62_89 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_62_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_63_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_63_154 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_63_164 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_63_201 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_63_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_63_28 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_63_284 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_63_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_63_351 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_63_40 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_63_417 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_63_431 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_63_445 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_63_484 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_63_503 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_63_505 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_63_522 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_63_543 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_63_557 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_63_561 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_63_565 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_63_569 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_63_585 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_63_60 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_63_604 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_63_614 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_63_617 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_63_658 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_63_708 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_63_712 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_63_98 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_64_144 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_64_189 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_64_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_64_224 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_64_245 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_64_266 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_64_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_64_306 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_64_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_64_356 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_64_363 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_64_389 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_64_399 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_64_470 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_64_477 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_64_488 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_64_494 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_64_52 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_64_530 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_64_541 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_64_587 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_64_589 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_64_62 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_64_637 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_64_709 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_64_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_64_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_65_119 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_65_158 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_65_179 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_65_206 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_65_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_65_234 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_65_277 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_65_292 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_65_298 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_65_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_65_33 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_65_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_65_337 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_65_351 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_65_449 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_65_466 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_65_503 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_65_505 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_65_545 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_65_590 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_65_617 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_65_653 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_65_681 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_65_693 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_65_710 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_65_73 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_66_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_66_128 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_66_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_66_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_66_217 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_66_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_66_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_66_283 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_66_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_66_302 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_66_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_66_313 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_66_338 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_66_363 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_66_38 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_66_454 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_66_475 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_66_477 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_66_504 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_66_512 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_66_517 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_66_529 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_66_613 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_66_64 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_66_642 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_66_654 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_66_674 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_66_709 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_66_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_67_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_67_155 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_67_212 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_67_327 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_67_34 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_67_363 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_67_391 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_67_447 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_67_452 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_67_465 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_67_482 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_67_514 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_67_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_67_544 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_67_552 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_67_569 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_67_590 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_67_607 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_67_634 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_67_638 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_67_66 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_67_670 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_67_692 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_67_709 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_68_101 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_68_122 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_68_128 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_68_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_68_156 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_68_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_68_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_68_235 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_68_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_68_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_68_296 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_68_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_68_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_68_365 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_68_377 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_68_381 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_68_453 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_68_463 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_68_475 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_68_477 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_68_558 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_68_587 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_68_609 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_68_617 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_68_635 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_68_64 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_68_683 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_68_70 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_68_74 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_68_78 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_68_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_68_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_68_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_69_108 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_69_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_69_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_69_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_69_222 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_69_230 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_69_235 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_69_243 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_69_255 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_69_262 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_69_267 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_69_286 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_69_362 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_69_381 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_69_447 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_69_449 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_69_46 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_69_488 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_69_501 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_69_514 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_69_534 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_69_570 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_69_584 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_69_634 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_6_112 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_6_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_148 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_6_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_6_175 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_6_191 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_213 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_6_230 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_6_266 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_6_285 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_6_304 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_6_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_313 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_354 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_6_365 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_6_387 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_395 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_453 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_6_470 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_6_493 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_512 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_6_529 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_533 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_6_584 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_589 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_6_608 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_616 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_624 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_629 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_6_641 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_6_645 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_6_659 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_668 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_6_677 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_685 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_699 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_6_704 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_6_71 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_712 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_75 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_6_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_70_132 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_70_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_70_182 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_70_208 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_70_212 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_70_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_70_257 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_70_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_70_291 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_70_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_70_325 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_70_360 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_70_402 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_70_419 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_70_421 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_70_489 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_70_514 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_70_533 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_70_544 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_70_560 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_70_581 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_70_589 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_70_612 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_70_618 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_70_63 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_70_645 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_70_674 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_70_72 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_70_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_70_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_71_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_71_120 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_71_132 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_71_136 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_71_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_71_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_71_205 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_71_236 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_71_246 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_71_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_71_285 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_71_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_71_306 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_71_331 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_71_335 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_71_354 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_71_391 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_71_401 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_71_410 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_71_432 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_71_440 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_71_512 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_71_528 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_71_532 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_71_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_71_557 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_71_583 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_71_607 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_71_625 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_71_630 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_71_653 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_71_657 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_71_671 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_71_673 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_71_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_71_98 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_72_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_72_16 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_72_160 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_72_201 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_72_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_72_231 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_72_249 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_72_271 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_72_290 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_72_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_72_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_72_329 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_72_359 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_72_363 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_72_381 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_72_392 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_72_411 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_72_429 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_72_433 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_72_44 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_72_456 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_72_493 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_72_527 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_72_533 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_72_543 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_72_561 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_72_589 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_72_602 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_72_608 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_72_628 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_72_635 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_72_643 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_72_661 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_72_682 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_72_690 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_72_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_72_712 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_72_74 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_72_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_72_95 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_73_104 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_73_108 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_73_146 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_73_156 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_73_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_73_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_73_206 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_73_212 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_73_218 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_73_222 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_73_244 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_73_262 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_73_266 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_73_269 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_73_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_73_28 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_73_316 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_73_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_73_34 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_73_380 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_73_390 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_73_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_73_417 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_73_447 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_73_456 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_73_476 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_73_491 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_73_520 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_73_535 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_73_559 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_73_584 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_73_594 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_73_599 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_73_633 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_73_64 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_73_641 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_73_712 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_73_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_74_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_117 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_74_120 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_172 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_74_179 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_74_200 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_224 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_74_230 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_74_243 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_74_25 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_74_285 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_74_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_74_304 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_34 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_74_342 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_346 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_358 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_74_373 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_74_399 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_74_418 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_74_425 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_443 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_452 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_74_466 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_493 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_74_510 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_74_520 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_74_529 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_74_551 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_56 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_603 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_74_645 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_651 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_74_67 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_681 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_74_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_75_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_122 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_75_135 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_75_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_150 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_158 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_75_178 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_75_206 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_212 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_75_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_75_252 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_263 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_75_290 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_335 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_75_342 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_75_37 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_391 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_75_398 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_447 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_75_456 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_75_485 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_491 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_75_500 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_75_505 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_75_52 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_75_522 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_537 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_75_600 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_624 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_75_640 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_644 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_680 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_75_72 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_75_92 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_76_100 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_76_136 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_76_157 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_76_191 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_76_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_76_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_76_230 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_76_236 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_76_278 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_76_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_76_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_76_305 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_76_373 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_76_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_76_436 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_76_44 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_76_462 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_76_469 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_76_48 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_76_483 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_76_493 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_76_498 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_76_506 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_76_530 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_76_587 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_76_589 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_76_604 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_76_613 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_76_635 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_76_645 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_76_75 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_76_92 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_77_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_77_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_77_14 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_77_151 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_77_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_77_201 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_77_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_77_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_77_24 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_77_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_77_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_77_345 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_77_391 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_77_402 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_77_449 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_77_45 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_77_466 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_77_485 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_77_503 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_77_505 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_77_523 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_77_527 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_77_544 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_77_556 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_77_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_77_596 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_77_614 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_77_620 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_77_628 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_77_633 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_77_650 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_77_94 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_77_99 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_78_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_78_157 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_78_176 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_78_222 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_78_226 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_78_245 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_78_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_78_306 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_78_32 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_78_320 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_78_338 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_78_350 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_78_356 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_78_363 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_78_370 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_78_398 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_78_442 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_78_454 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_78_469 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_78_475 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_78_490 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_78_499 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_78_507 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_78_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_78_530 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_78_533 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_78_559 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_78_570 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_78_586 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_78_609 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_78_617 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_78_623 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_78_640 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_78_72 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_79_12 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_79_129 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_79_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_79_151 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_79_193 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_79_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_79_259 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_79_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_79_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_79_300 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_79_310 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_79_314 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_79_325 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_79_352 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_79_370 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_79_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_79_396 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_79_421 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_79_43 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_79_471 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_79_480 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_79_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_79_545 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_79_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_79_587 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_79_605 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_79_613 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_79_671 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_79_75 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_79_98 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_7_121 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_129 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_7_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_7_162 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_7_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_7_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_222 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_7_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_7_261 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_7_276 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_7_297 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_30 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_7_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_337 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_7_355 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_363 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_7_393 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_7_405 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_409 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_7_434 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_438 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_447 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_449 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_7_458 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_462 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_503 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_7_545 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_7_556 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_565 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_569 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_7_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_7_583 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_602 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_7_607 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_7_621 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_7_669 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_673 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_679 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_79 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_80_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_80_157 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_80_175 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_80_192 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_80_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_80_220 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_80_241 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_80_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_80_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_80_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_80_325 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_80_358 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_80_365 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_80_369 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_80_386 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_80_393 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_80_410 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_80_415 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_80_419 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_80_449 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_80_474 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_80_477 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_80_487 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_80_491 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_80_502 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_80_530 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_80_533 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_80_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_80_551 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_80_559 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_80_561 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_80_567 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_80_587 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_80_589 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_80_611 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_80_615 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_80_617 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_80_623 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_80_66 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_80_670 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_80_699 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_80_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_80_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_80_89 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_103 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_8_112 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_8_134 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_8_149 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_206 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_8_240 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_8_278 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_8_305 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_317 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_8_326 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_338 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_365 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_8_395 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_8_414 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_8_421 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_8_440 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_444 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_8_45 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_8_469 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_475 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_8_477 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_8_528 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_8_541 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_558 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_8_576 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_580 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_8_585 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_8_589 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_593 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_8_598 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_606 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_8_628 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_8_641 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_8_645 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_653 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_659 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_8_687 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_691 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_701 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_8_75 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_9_107 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_9_129 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_135 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_9_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_183 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_9_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_9_211 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_9_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_229 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_262 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_9_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_335 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_337 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_346 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_355 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_367 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_9_376 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_9_417 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_425 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_43 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_435 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_9_445 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_9_481 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_9_492 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_9_513 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_521 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_9_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_538 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_9_548 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_9_566 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_9_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_9_574 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_584 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_9_589 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_598 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_9_607 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_615 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_617 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_9_629 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_63 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_633 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_9_642 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_650 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_660 (.VGND(VGND),
    .VPWR(VPWR),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_9_686 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_9_88 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_91 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_92 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_94 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_95 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_96 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_98 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_99 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_100 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_101 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_102 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_103 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_104 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_106 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_107 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_108 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_112 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_114 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_115 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_116 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_117 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_118 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_119 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Left_120 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Right_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_84 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Left_121 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Right_40 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Left_122 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Right_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Left_123 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Right_42 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Left_124 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Right_43 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Left_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Right_44 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Left_126 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Right_45 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Left_127 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Right_46 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Left_128 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Right_47 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Left_129 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Right_48 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Left_130 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Right_49 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Left_131 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Right_50 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Left_132 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Right_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Left_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Right_52 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Left_134 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Right_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Left_135 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Right_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Left_136 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Right_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Left_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Right_56 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Left_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Right_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Left_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Right_58 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Left_140 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Right_59 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_86 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Left_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Right_60 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Left_142 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Right_61 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Left_143 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Right_62 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Left_144 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Right_63 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Left_145 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Right_64 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Left_146 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Right_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Left_147 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Right_66 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Left_148 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Right_67 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Left_149 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Right_68 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Left_150 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Right_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_87 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Left_151 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Right_70 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Left_152 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Right_71 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Left_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Right_72 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Left_154 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Right_73 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Left_155 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Right_74 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Left_156 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Right_75 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Left_157 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Right_76 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Left_158 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Right_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Left_159 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Right_78 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Left_160 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Right_79 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_88 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Left_161 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Right_80 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_89 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_90 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_162 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_163 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_164 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_165 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_166 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_167 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_168 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_169 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_170 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_171 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_172 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_173 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_174 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_175 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_176 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_177 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_178 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_179 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_180 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_181 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_182 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_183 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_184 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_185 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_186 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_299 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_300 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_301 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_302 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_303 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_304 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_305 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_306 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_307 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_308 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_309 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_310 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_311 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_312 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_313 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_314 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_315 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_316 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_317 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_318 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_319 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_320 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_321 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_322 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_323 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_324 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_325 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_326 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_327 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_328 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_329 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_330 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_331 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_332 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_333 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_334 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_335 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_336 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_337 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_338 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_339 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_340 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_341 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_342 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_343 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_344 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_345 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_346 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_347 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_348 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_349 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_350 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_351 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_352 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_353 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_354 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_355 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_356 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_357 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_358 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_359 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_360 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_361 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_362 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_363 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_364 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_365 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_366 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_367 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_368 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_369 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_370 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_371 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_372 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_373 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_374 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_375 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_376 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_377 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_378 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_379 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_380 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_381 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_382 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_383 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_384 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_385 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_386 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_387 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_388 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_389 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_390 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_391 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_392 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_393 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_394 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_395 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_396 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_397 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_398 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_399 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_400 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_401 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_402 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_403 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_404 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_405 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_406 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_407 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_408 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_409 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_410 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_411 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_412 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_413 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_414 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_415 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_416 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_417 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_418 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_419 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_420 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_421 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_422 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_423 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_187 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_188 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_189 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_190 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_191 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_192 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_193 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_194 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_195 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_196 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_197 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_198 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_424 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_425 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_426 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_427 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_428 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_429 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_430 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_431 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_432 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_433 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_434 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_435 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_436 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_437 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_438 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_439 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_440 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_441 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_442 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_443 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_444 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_445 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_446 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_447 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_448 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_449 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_450 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_451 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_452 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_453 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_454 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_455 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_456 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_457 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_458 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_459 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_460 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_461 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_462 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_463 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_464 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_465 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_466 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_467 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_468 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_469 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_470 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_471 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_472 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_473 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_474 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_475 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_476 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_477 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_478 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_479 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_480 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_481 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_482 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_483 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_484 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_485 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_486 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_487 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_488 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_489 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_490 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_491 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_492 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_493 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_494 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_495 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_496 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_497 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_498 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_499 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_500 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_501 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_502 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_503 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_504 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_505 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_506 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_507 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_508 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_509 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_510 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_511 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_512 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_513 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_514 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_515 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_516 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_517 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_518 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_519 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_520 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_521 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_522 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_523 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_524 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_525 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_526 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_527 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_528 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_529 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_530 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_531 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_532 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_533 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_534 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_535 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_536 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_537 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_538 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_539 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_540 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_541 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_542 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_543 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_544 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_545 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_546 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_547 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_548 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_199 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_200 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_201 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_202 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_203 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_204 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_205 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_206 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_207 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_208 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_209 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_210 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_211 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_549 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_550 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_551 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_552 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_553 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_554 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_555 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_556 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_557 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_558 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_559 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_560 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_561 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_562 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_563 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_564 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_565 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_566 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_567 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_568 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_569 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_570 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_571 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_572 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_573 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_574 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_575 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_576 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_577 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_578 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_579 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_580 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_581 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_582 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_583 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_584 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_585 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_586 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_587 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_588 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_589 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_590 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_591 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_592 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_593 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_594 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_595 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_596 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_597 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_598 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_599 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_600 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_601 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_602 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_603 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_604 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_605 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_606 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_607 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_608 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_609 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_610 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_611 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_612 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_613 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_614 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_615 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_616 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_617 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_618 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_619 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_620 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_621 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_622 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_623 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_624 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_625 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_626 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_627 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_628 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_629 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_630 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_631 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_632 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_633 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_634 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_635 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_636 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_637 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_638 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_639 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_640 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_641 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_642 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_643 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_644 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_645 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_646 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_647 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_648 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_649 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_650 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_651 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_652 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_653 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_654 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_655 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_656 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_657 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_658 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_659 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_660 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_661 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_662 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_663 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_664 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_665 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_666 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_667 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_668 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_669 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_670 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_671 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_672 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_673 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_212 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_213 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_214 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_215 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_216 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_217 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_218 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_219 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_220 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_221 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_222 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_223 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_674 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_675 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_676 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_677 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_678 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_679 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_680 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_681 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_682 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_683 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_684 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_685 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_686 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_687 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_688 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_689 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_690 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_691 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_692 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_693 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_694 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_695 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_696 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_697 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_698 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_699 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_700 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_701 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_702 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_703 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_704 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_705 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_706 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_707 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_708 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_709 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_710 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_711 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_712 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_713 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_714 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_715 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_716 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_717 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_718 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_719 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_720 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_721 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_722 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_723 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_724 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_725 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_726 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_727 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_728 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_729 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_730 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_731 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_732 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_733 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_734 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_735 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_736 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_737 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_738 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_739 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_740 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_741 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_742 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_743 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_744 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_745 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_746 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_747 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_748 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_749 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_750 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_751 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_752 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_753 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_754 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_755 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_756 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_757 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_758 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_759 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_760 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_761 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_762 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_763 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_764 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_765 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_766 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_767 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_768 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_769 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_770 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_771 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_772 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_773 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_774 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_775 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_776 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_777 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_778 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_779 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_780 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_781 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_782 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_783 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_784 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_785 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_786 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_787 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_788 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_789 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_790 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_791 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_792 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_793 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_794 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_795 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_796 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_797 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_798 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_224 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_225 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_226 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_227 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_228 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_229 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_230 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_231 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_232 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_233 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_234 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_235 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_236 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_799 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_800 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_801 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_802 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_803 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_804 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_805 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_806 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_807 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_808 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_809 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_810 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_811 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_812 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_813 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_814 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_815 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_816 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_817 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_818 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_819 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_820 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_821 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_822 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_823 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_824 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_825 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_826 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_827 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_828 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_829 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_830 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_831 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_832 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_833 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_834 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_835 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_836 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_837 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_838 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_839 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_840 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_841 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_842 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_843 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_844 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_845 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_846 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_847 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_848 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_849 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_850 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_851 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_852 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_853 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_854 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_855 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_856 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_857 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_858 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_859 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_860 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_861 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_862 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_863 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_864 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_865 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_866 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_867 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_868 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_869 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_870 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_871 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_872 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_873 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_874 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_875 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_876 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_877 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_878 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_879 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_880 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_881 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_882 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_883 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_884 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_885 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_886 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_887 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_888 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_889 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_890 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_891 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_892 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_893 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_894 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_895 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_896 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_897 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_898 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_899 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_900 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_901 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_902 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_903 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_904 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_905 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_906 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_907 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_908 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_909 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_910 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_911 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_912 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_913 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_914 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_915 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_916 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_917 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_918 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_919 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_920 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_921 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_922 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_923 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_237 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_238 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_239 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_240 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_241 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_242 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_243 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_244 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_245 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_246 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_247 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_248 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_924 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_925 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_926 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_927 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_928 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_929 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_930 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_931 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_932 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_933 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_934 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_935 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_936 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_937 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_938 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_939 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_940 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_941 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_942 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_943 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_944 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_945 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_946 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_947 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_948 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_949 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_950 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_951 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_952 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_953 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_954 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_955 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_956 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_957 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_958 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_959 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_960 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_961 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_962 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_963 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_964 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_965 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_966 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_967 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_968 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_969 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_970 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_971 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_972 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_973 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_974 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_975 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_976 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_977 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_978 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_979 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_980 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_981 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_982 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_983 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_984 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_985 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_986 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_987 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_988 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_989 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_990 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_991 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_992 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_993 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_994 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_995 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_996 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_997 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_998 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1000 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1001 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1002 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1003 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1004 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1005 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1006 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1007 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1008 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1009 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1010 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1011 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_999 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1012 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1013 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1014 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1015 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1016 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1017 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1018 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1019 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1020 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1021 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1022 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1023 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1024 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1025 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1026 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1027 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1028 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1029 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1030 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1031 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1032 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1033 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1034 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1035 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1036 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1037 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1038 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1039 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1040 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1041 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1042 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1043 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1044 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1045 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1046 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1047 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1048 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_249 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_250 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_251 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_252 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_253 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_254 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_255 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_256 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_257 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_258 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_259 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_260 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_261 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1049 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1050 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1051 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1052 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1053 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1054 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1055 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1056 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1057 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1058 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1059 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1060 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1061 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1062 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1063 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1064 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1065 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1066 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1067 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1068 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1069 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1070 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1071 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1072 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1073 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1074 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1075 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1076 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1077 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1078 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1079 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1080 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1081 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1082 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1083 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1084 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1085 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1086 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1087 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1088 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1089 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1090 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1091 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1092 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1093 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1094 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1095 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1096 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1097 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1098 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1099 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1100 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1101 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1102 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1103 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1104 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1105 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1106 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1107 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1108 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1109 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1110 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1111 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1112 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1113 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1114 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1115 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1116 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1117 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1118 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1119 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1120 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1121 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1122 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1123 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1124 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1125 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1126 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1127 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1128 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1129 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1130 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1131 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1132 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1133 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1134 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1135 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1136 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1137 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1138 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1139 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1140 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1141 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1142 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1143 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1144 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1145 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1146 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1147 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1148 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1149 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1150 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1151 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1152 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1153 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1154 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1155 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1156 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1157 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1158 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1159 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1160 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1161 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1162 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1163 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1164 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1165 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1166 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1167 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1168 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1169 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1170 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1171 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1172 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1173 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_262 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_263 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_264 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_265 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_266 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_267 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_268 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_269 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_270 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_271 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_272 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_273 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1174 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1175 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1176 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1177 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1178 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1179 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1180 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1181 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1182 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1183 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1184 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1185 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1186 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1187 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1188 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1189 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1190 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1191 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1192 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1193 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1194 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1195 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1196 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1197 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1198 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_274 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_275 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_276 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_277 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_278 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_279 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_280 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_281 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_282 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_283 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_284 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_285 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_286 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_287 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_288 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_289 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_290 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_291 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_292 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_293 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_294 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_295 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_296 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_297 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_298 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_2 _3755_ (.A(\i_tinyqv.cpu.counter[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0607_));
 sky130_fd_sc_hd__clkbuf_4 _3756_ (.A(\i_tinyqv.cpu.counter[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0608_));
 sky130_fd_sc_hd__or2b_1 _3757_ (.A(\i_tinyqv.cpu.counter[3] ),
    .B_N(_0608_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0609_));
 sky130_fd_sc_hd__nor2_2 _3758_ (.A(_0607_),
    .B(_0609_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0610_));
 sky130_fd_sc_hd__clkbuf_4 _3759_ (.A(_0607_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0611_));
 sky130_fd_sc_hd__or2_4 _3760_ (.A(\i_tinyqv.cpu.counter[3] ),
    .B(_0608_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0612_));
 sky130_fd_sc_hd__nor2_2 _3761_ (.A(_0611_),
    .B(_0612_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0613_));
 sky130_fd_sc_hd__buf_4 _3762_ (.A(\i_tinyqv.cpu.counter[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0614_));
 sky130_fd_sc_hd__nor2_2 _3763_ (.A(_0614_),
    .B(_0608_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0615_));
 sky130_fd_sc_hd__and2_1 _3764_ (.A(\i_tinyqv.cpu.counter[3] ),
    .B(\i_tinyqv.cpu.counter[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0616_));
 sky130_fd_sc_hd__buf_2 _3765_ (.A(_0616_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0617_));
 sky130_fd_sc_hd__a22o_1 _3766_ (.A1(\i_tinyqv.cpu.instr_data_start[3] ),
    .A2(_0615_),
    .B1(_0617_),
    .B2(\i_tinyqv.cpu.instr_data_start[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0618_));
 sky130_fd_sc_hd__nor2b_4 _3767_ (.A(_0614_),
    .B_N(_0608_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0619_));
 sky130_fd_sc_hd__and2b_2 _3768_ (.A_N(\i_tinyqv.cpu.counter[2] ),
    .B(\i_tinyqv.cpu.counter[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0620_));
 sky130_fd_sc_hd__a22o_1 _3769_ (.A1(\i_tinyqv.cpu.instr_data_start[7] ),
    .A2(_0619_),
    .B1(_0620_),
    .B2(\i_tinyqv.cpu.instr_data_start[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0621_));
 sky130_fd_sc_hd__o21a_1 _3770_ (.A1(_0618_),
    .A2(_0621_),
    .B1(_0611_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0622_));
 sky130_fd_sc_hd__a221o_1 _3771_ (.A1(\i_tinyqv.cpu.instr_data_start[23] ),
    .A2(_0610_),
    .B1(_0613_),
    .B2(\i_tinyqv.cpu.instr_data_start[19] ),
    .C1(_0622_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0623_));
 sky130_fd_sc_hd__buf_4 _3772_ (.A(\i_tinyqv.cpu.i_core.i_registers.rs1[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0624_));
 sky130_fd_sc_hd__buf_6 _3773_ (.A(\i_tinyqv.cpu.i_core.i_registers.rs1[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0625_));
 sky130_fd_sc_hd__buf_6 _3774_ (.A(\i_tinyqv.cpu.i_core.i_registers.rs1[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0626_));
 sky130_fd_sc_hd__buf_4 _3775_ (.A(\i_tinyqv.cpu.i_core.i_registers.rs1[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0627_));
 sky130_fd_sc_hd__and4b_1 _3776_ (.A_N(_0624_),
    .B(_0625_),
    .C(net324),
    .D(_0627_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0628_));
 sky130_fd_sc_hd__or4b_1 _3777_ (.A(\i_tinyqv.cpu.i_core.i_registers.rs1[0] ),
    .B(net53),
    .C(net56),
    .D_N(net52),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0629_));
 sky130_fd_sc_hd__nand3b_2 _3778_ (.A_N(\i_tinyqv.cpu.counter[2] ),
    .B(_0614_),
    .C(\i_tinyqv.cpu.counter[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0630_));
 sky130_fd_sc_hd__and4bb_1 _3779_ (.A_N(\i_tinyqv.cpu.i_core.i_registers.rs1[0] ),
    .B_N(\i_tinyqv.cpu.i_core.i_registers.rs1[1] ),
    .C(\i_tinyqv.cpu.i_core.i_registers.rs1[2] ),
    .D(\i_tinyqv.cpu.i_core.i_registers.rs1[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0631_));
 sky130_fd_sc_hd__a2bb2o_1 _3780_ (.A1_N(_0629_),
    .A2_N(_0630_),
    .B1(_0631_),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[12][3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0632_));
 sky130_fd_sc_hd__and4_1 _3781_ (.A(_0627_),
    .B(net53),
    .C(net52),
    .D(net56),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0633_));
 sky130_fd_sc_hd__nor4b_1 _3782_ (.A(_0627_),
    .B(_0624_),
    .C(_0625_),
    .D_N(_0626_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0634_));
 sky130_fd_sc_hd__a22o_1 _3783_ (.A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[15][3] ),
    .A2(_0633_),
    .B1(net321),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[8][3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0635_));
 sky130_fd_sc_hd__a211o_4 _3784_ (.A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[13][3] ),
    .A2(net62),
    .B1(_0632_),
    .C1(_0635_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0636_));
 sky130_fd_sc_hd__and4b_2 _3785_ (.A_N(_0625_),
    .B(net324),
    .C(_0627_),
    .D(_0624_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0637_));
 sky130_fd_sc_hd__nor4b_2 _3786_ (.A(_0627_),
    .B(_0625_),
    .C(_0626_),
    .D_N(_0624_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0638_));
 sky130_fd_sc_hd__and4bb_2 _3787_ (.A_N(_0627_),
    .B_N(_0626_),
    .C(_0625_),
    .D(_0624_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0639_));
 sky130_fd_sc_hd__a22o_1 _3788_ (.A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[2][3] ),
    .A2(_0638_),
    .B1(_0639_),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[6][3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0640_));
 sky130_fd_sc_hd__a21o_1 _3789_ (.A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[11][3] ),
    .A2(_0637_),
    .B1(_0640_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0641_));
 sky130_fd_sc_hd__and4bb_2 _3790_ (.A_N(_0624_),
    .B_N(_0625_),
    .C(net324),
    .D(_0627_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0642_));
 sky130_fd_sc_hd__and4b_1 _3791_ (.A_N(\i_tinyqv.cpu.i_core.i_registers.rs1[0] ),
    .B(net70),
    .C(net51),
    .D(net30),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0643_));
 sky130_fd_sc_hd__and2_1 _3792_ (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[14][3] ),
    .B(_0643_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0644_));
 sky130_fd_sc_hd__and4bb_1 _3793_ (.A_N(\i_tinyqv.cpu.i_core.i_registers.rs1[1] ),
    .B_N(\i_tinyqv.cpu.i_core.i_registers.rs1[3] ),
    .C(\i_tinyqv.cpu.i_core.i_registers.rs1[2] ),
    .D(\i_tinyqv.cpu.i_core.i_registers.rs1[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0645_));
 sky130_fd_sc_hd__and4bb_1 _3794_ (.A_N(\i_tinyqv.cpu.i_core.i_registers.rs1[0] ),
    .B_N(\i_tinyqv.cpu.i_core.i_registers.rs1[2] ),
    .C(\i_tinyqv.cpu.i_core.i_registers.rs1[3] ),
    .D(\i_tinyqv.cpu.i_core.i_registers.rs1[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0646_));
 sky130_fd_sc_hd__a22o_1 _3795_ (.A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[5][3] ),
    .A2(_0645_),
    .B1(_0646_),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[10][3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0647_));
 sky130_fd_sc_hd__nor4b_4 _3796_ (.A(_0624_),
    .B(_0625_),
    .C(_0626_),
    .D_N(net87),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0648_));
 sky130_fd_sc_hd__and4b_1 _3797_ (.A_N(_0626_),
    .B(_0625_),
    .C(_0624_),
    .D(_0627_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0649_));
 sky130_fd_sc_hd__a22o_1 _3798_ (.A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[1][3] ),
    .A2(_0648_),
    .B1(_0649_),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[7][3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0650_));
 sky130_fd_sc_hd__a2111o_1 _3799_ (.A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[9][3] ),
    .A2(_0642_),
    .B1(_0644_),
    .C1(_0647_),
    .D1(_0650_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0651_));
 sky130_fd_sc_hd__or3_4 _3800_ (.A(_0636_),
    .B(_0641_),
    .C(_0651_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0652_));
 sky130_fd_sc_hd__buf_4 _3801_ (.A(\i_tinyqv.cpu.debug_instr_valid ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0653_));
 sky130_fd_sc_hd__o21ai_4 _3802_ (.A1(\i_tinyqv.cpu.is_jal ),
    .A2(\i_tinyqv.cpu.is_auipc ),
    .B1(_0653_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0654_));
 sky130_fd_sc_hd__mux2_4 _3803_ (.A0(_0623_),
    .A1(_0652_),
    .S(_0654_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0655_));
 sky130_fd_sc_hd__clkbuf_4 _3804_ (.A(\i_tinyqv.cpu.alu_op[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0656_));
 sky130_fd_sc_hd__or2_1 _3805_ (.A(_0656_),
    .B(\i_tinyqv.cpu.alu_op[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0657_));
 sky130_fd_sc_hd__clkbuf_2 _3806_ (.A(_0657_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0658_));
 sky130_fd_sc_hd__or4b_1 _3807_ (.A(net38),
    .B(net37),
    .C(\i_tinyqv.cpu.i_core.i_registers.rs2[3] ),
    .D_N(\i_tinyqv.cpu.i_core.i_registers.rs2[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0659_));
 sky130_fd_sc_hd__buf_2 _3808_ (.A(\i_tinyqv.cpu.i_core.i_registers.rs2[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0660_));
 sky130_fd_sc_hd__buf_2 _3809_ (.A(\i_tinyqv.cpu.i_core.i_registers.rs2[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0661_));
 sky130_fd_sc_hd__buf_2 _3810_ (.A(\i_tinyqv.cpu.i_core.i_registers.rs2[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0662_));
 sky130_fd_sc_hd__buf_6 _3811_ (.A(\i_tinyqv.cpu.i_core.i_registers.rs2[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0663_));
 sky130_fd_sc_hd__and4b_1 _3812_ (.A_N(_0660_),
    .B(_0661_),
    .C(_0662_),
    .D(_0663_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0664_));
 sky130_fd_sc_hd__a2bb2o_1 _3813_ (.A1_N(_0630_),
    .A2_N(_0659_),
    .B1(_0664_),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[11][3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0665_));
 sky130_fd_sc_hd__and2b_1 _3814_ (.A_N(_0660_),
    .B(_0661_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0666_));
 sky130_fd_sc_hd__nor2b_2 _3815_ (.A(net39),
    .B_N(_0663_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0667_));
 sky130_fd_sc_hd__and4b_2 _3816_ (.A_N(_0662_),
    .B(_0663_),
    .C(_0660_),
    .D(\i_tinyqv.cpu.i_core.i_registers.rs2[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0668_));
 sky130_fd_sc_hd__a32o_1 _3817_ (.A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[10][3] ),
    .A2(_0666_),
    .A3(_0667_),
    .B1(_0668_),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[14][3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0669_));
 sky130_fd_sc_hd__nor2_2 _3818_ (.A(_0660_),
    .B(_0661_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0670_));
 sky130_fd_sc_hd__nor4b_2 _3819_ (.A(_0662_),
    .B(_0663_),
    .C(_0660_),
    .D_N(_0661_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0671_));
 sky130_fd_sc_hd__a32o_1 _3820_ (.A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[2][3] ),
    .A2(_0667_),
    .A3(_0670_),
    .B1(net25),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[8][3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0672_));
 sky130_fd_sc_hd__or3_1 _3821_ (.A(_0665_),
    .B(_0669_),
    .C(_0672_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0673_));
 sky130_fd_sc_hd__and4bb_2 _3822_ (.A_N(net38),
    .B_N(net37),
    .C(\i_tinyqv.cpu.i_core.i_registers.rs2[2] ),
    .D(\i_tinyqv.cpu.i_core.i_registers.rs2[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0674_));
 sky130_fd_sc_hd__and4bb_2 _3823_ (.A_N(_0663_),
    .B_N(\i_tinyqv.cpu.i_core.i_registers.rs2[3] ),
    .C(\i_tinyqv.cpu.i_core.i_registers.rs2[2] ),
    .D(net38),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0675_));
 sky130_fd_sc_hd__a22o_1 _3824_ (.A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[12][3] ),
    .A2(_0674_),
    .B1(_0675_),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[5][3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0676_));
 sky130_fd_sc_hd__and4_2 _3825_ (.A(net38),
    .B(net37),
    .C(\i_tinyqv.cpu.i_core.i_registers.rs2[2] ),
    .D(\i_tinyqv.cpu.i_core.i_registers.rs2[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0677_));
 sky130_fd_sc_hd__and4b_2 _3826_ (.A_N(_0661_),
    .B(\i_tinyqv.cpu.i_core.i_registers.rs2[2] ),
    .C(net37),
    .D(net38),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0678_));
 sky130_fd_sc_hd__a22o_1 _3827_ (.A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[15][3] ),
    .A2(_0677_),
    .B1(_0678_),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[7][3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0679_));
 sky130_fd_sc_hd__and4bb_2 _3828_ (.A_N(net37),
    .B_N(\i_tinyqv.cpu.i_core.i_registers.rs2[2] ),
    .C(\i_tinyqv.cpu.i_core.i_registers.rs2[3] ),
    .D(net38),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0680_));
 sky130_fd_sc_hd__and4bb_2 _3829_ (.A_N(_0662_),
    .B_N(_0661_),
    .C(\i_tinyqv.cpu.i_core.i_registers.rs2[2] ),
    .D(net37),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0681_));
 sky130_fd_sc_hd__a22o_1 _3830_ (.A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[9][3] ),
    .A2(_0680_),
    .B1(_0681_),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[6][3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0682_));
 sky130_fd_sc_hd__nor4b_1 _3831_ (.A(_0663_),
    .B(_0660_),
    .C(_0661_),
    .D_N(_0662_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0683_));
 sky130_fd_sc_hd__and4b_2 _3832_ (.A_N(_0663_),
    .B(_0660_),
    .C(_0661_),
    .D(_0662_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0684_));
 sky130_fd_sc_hd__a22o_1 _3833_ (.A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[1][3] ),
    .A2(net24),
    .B1(_0684_),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[13][3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0685_));
 sky130_fd_sc_hd__or4_4 _3834_ (.A(_0676_),
    .B(_0679_),
    .C(_0682_),
    .D(_0685_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0686_));
 sky130_fd_sc_hd__nor2_2 _3835_ (.A(_0673_),
    .B(_0686_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0687_));
 sky130_fd_sc_hd__clkbuf_8 _3836_ (.A(\i_tinyqv.cpu.counter[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0688_));
 sky130_fd_sc_hd__buf_4 _3837_ (.A(_0615_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0689_));
 sky130_fd_sc_hd__clkbuf_4 _3838_ (.A(_0620_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0690_));
 sky130_fd_sc_hd__clkbuf_4 _3839_ (.A(_0690_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0691_));
 sky130_fd_sc_hd__a22o_1 _3840_ (.A1(\i_tinyqv.cpu.imm[15] ),
    .A2(_0617_),
    .B1(_0619_),
    .B2(\i_tinyqv.cpu.i_core.imm_lo[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0692_));
 sky130_fd_sc_hd__a221o_1 _3841_ (.A1(\i_tinyqv.cpu.i_core.imm_lo[3] ),
    .A2(_0689_),
    .B1(_0691_),
    .B2(\i_tinyqv.cpu.i_core.imm_lo[11] ),
    .C1(_0692_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0693_));
 sky130_fd_sc_hd__and3_1 _3842_ (.A(_0614_),
    .B(_0608_),
    .C(\i_tinyqv.cpu.imm[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0694_));
 sky130_fd_sc_hd__a221o_1 _3843_ (.A1(\i_tinyqv.cpu.imm[23] ),
    .A2(_0619_),
    .B1(_0690_),
    .B2(\i_tinyqv.cpu.imm[27] ),
    .C1(_0694_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0695_));
 sky130_fd_sc_hd__a211o_1 _3844_ (.A1(\i_tinyqv.cpu.imm[19] ),
    .A2(_0689_),
    .B1(_0695_),
    .C1(_0611_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0696_));
 sky130_fd_sc_hd__o21ai_2 _3845_ (.A1(_0688_),
    .A2(_0693_),
    .B1(_0696_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0697_));
 sky130_fd_sc_hd__o21ai_4 _3846_ (.A1(\i_tinyqv.cpu.is_branch ),
    .A2(\i_tinyqv.cpu.is_alu_reg ),
    .B1(\i_tinyqv.cpu.debug_instr_valid ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0698_));
 sky130_fd_sc_hd__mux2_4 _3847_ (.A0(_0687_),
    .A1(_0697_),
    .S(_0698_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0699_));
 sky130_fd_sc_hd__xnor2_1 _3848_ (.A(_0658_),
    .B(_0699_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0700_));
 sky130_fd_sc_hd__or2_1 _3849_ (.A(net80),
    .B(_0700_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0701_));
 sky130_fd_sc_hd__inv_2 _3850_ (.A(_0698_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0702_));
 sky130_fd_sc_hd__a22o_1 _3851_ (.A1(\i_tinyqv.cpu.imm[12] ),
    .A2(_0617_),
    .B1(_0619_),
    .B2(\i_tinyqv.cpu.i_core.imm_lo[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0703_));
 sky130_fd_sc_hd__a221o_1 _3852_ (.A1(\i_tinyqv.cpu.i_core.imm_lo[0] ),
    .A2(_0615_),
    .B1(_0620_),
    .B2(\i_tinyqv.cpu.i_core.imm_lo[8] ),
    .C1(\i_tinyqv.cpu.counter[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0704_));
 sky130_fd_sc_hd__mux4_1 _3853_ (.A0(\i_tinyqv.cpu.imm[16] ),
    .A1(\i_tinyqv.cpu.imm[20] ),
    .A2(\i_tinyqv.cpu.imm[24] ),
    .A3(\i_tinyqv.cpu.imm[28] ),
    .S0(_0608_),
    .S1(_0614_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0705_));
 sky130_fd_sc_hd__nor2_1 _3854_ (.A(_0611_),
    .B(_0705_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0706_));
 sky130_fd_sc_hd__o21bai_4 _3855_ (.A1(_0703_),
    .A2(_0704_),
    .B1_N(_0706_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0707_));
 sky130_fd_sc_hd__nor2_2 _3856_ (.A(_0702_),
    .B(_0707_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0708_));
 sky130_fd_sc_hd__a22o_1 _3857_ (.A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[15][0] ),
    .A2(_0677_),
    .B1(net24),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[1][0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0709_));
 sky130_fd_sc_hd__a32o_1 _3858_ (.A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[2][0] ),
    .A2(_0667_),
    .A3(_0670_),
    .B1(net25),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[8][0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0710_));
 sky130_fd_sc_hd__and2_1 _3859_ (.A(_0662_),
    .B(_0663_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0711_));
 sky130_fd_sc_hd__and4_1 _3860_ (.A(\i_tinyqv.cpu.counter[4] ),
    .B(_0620_),
    .C(_0711_),
    .D(_0670_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0712_));
 sky130_fd_sc_hd__a22o_1 _3861_ (.A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[11][0] ),
    .A2(_0664_),
    .B1(_0678_),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[7][0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0713_));
 sky130_fd_sc_hd__nor4_1 _3862_ (.A(_0709_),
    .B(_0710_),
    .C(_0712_),
    .D(_0713_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0714_));
 sky130_fd_sc_hd__and3_1 _3863_ (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[10][0] ),
    .B(_0666_),
    .C(_0667_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0715_));
 sky130_fd_sc_hd__a22o_1 _3864_ (.A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[14][0] ),
    .A2(_0668_),
    .B1(_0680_),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[9][0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0716_));
 sky130_fd_sc_hd__a22o_1 _3865_ (.A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[12][0] ),
    .A2(_0674_),
    .B1(_0684_),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[13][0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0717_));
 sky130_fd_sc_hd__a22o_1 _3866_ (.A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[5][0] ),
    .A2(_0675_),
    .B1(_0681_),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[6][0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0718_));
 sky130_fd_sc_hd__nor4_2 _3867_ (.A(_0715_),
    .B(_0716_),
    .C(_0717_),
    .D(_0718_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0719_));
 sky130_fd_sc_hd__a21oi_2 _3868_ (.A1(net23),
    .A2(net21),
    .B1(_0698_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0720_));
 sky130_fd_sc_hd__or3_4 _3869_ (.A(_0658_),
    .B(_0708_),
    .C(_0720_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0721_));
 sky130_fd_sc_hd__o21ai_1 _3870_ (.A1(_0708_),
    .A2(net77),
    .B1(_0658_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0722_));
 sky130_fd_sc_hd__and3_1 _3871_ (.A(\i_tinyqv.cpu.instr_data_start[8] ),
    .B(_0611_),
    .C(_0690_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0723_));
 sky130_fd_sc_hd__nand2_4 _3872_ (.A(_0614_),
    .B(_0608_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0724_));
 sky130_fd_sc_hd__nor2_1 _3873_ (.A(\i_tinyqv.cpu.counter[4] ),
    .B(_0724_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0725_));
 sky130_fd_sc_hd__clkbuf_4 _3874_ (.A(\i_tinyqv.cpu.instr_data_start[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0726_));
 sky130_fd_sc_hd__a22o_1 _3875_ (.A1(\i_tinyqv.cpu.instr_data_start[20] ),
    .A2(_0610_),
    .B1(_0725_),
    .B2(_0726_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0727_));
 sky130_fd_sc_hd__a32o_1 _3876_ (.A1(\i_tinyqv.cpu.instr_data_start[4] ),
    .A2(_0611_),
    .A3(_0619_),
    .B1(_0613_),
    .B2(\i_tinyqv.cpu.instr_data_start[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0728_));
 sky130_fd_sc_hd__or3_2 _3877_ (.A(_0723_),
    .B(_0727_),
    .C(_0728_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0729_));
 sky130_fd_sc_hd__a22o_1 _3878_ (.A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[12][0] ),
    .A2(net74),
    .B1(_0642_),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[9][0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0730_));
 sky130_fd_sc_hd__a22o_1 _3879_ (.A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[13][0] ),
    .A2(_0628_),
    .B1(_0646_),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[10][0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0731_));
 sky130_fd_sc_hd__and2_1 _3880_ (.A(_0627_),
    .B(_0624_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0732_));
 sky130_fd_sc_hd__nor2_1 _3881_ (.A(_0625_),
    .B(net324),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0733_));
 sky130_fd_sc_hd__and4_1 _3882_ (.A(\i_tinyqv.cpu.counter[4] ),
    .B(_0690_),
    .C(_0732_),
    .D(_0733_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0734_));
 sky130_fd_sc_hd__a22o_1 _3883_ (.A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[6][0] ),
    .A2(_0639_),
    .B1(net55),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[7][0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0735_));
 sky130_fd_sc_hd__nor4_2 _3884_ (.A(_0730_),
    .B(_0731_),
    .C(_0734_),
    .D(_0735_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0736_));
 sky130_fd_sc_hd__a22o_1 _3885_ (.A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[15][0] ),
    .A2(net84),
    .B1(net47),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[14][0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0737_));
 sky130_fd_sc_hd__a22o_1 _3886_ (.A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[5][0] ),
    .A2(net58),
    .B1(_0637_),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[11][0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0738_));
 sky130_fd_sc_hd__a22o_1 _3887_ (.A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[8][0] ),
    .A2(net321),
    .B1(_0638_),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[2][0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0739_));
 sky130_fd_sc_hd__a2111oi_4 _3888_ (.A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[1][0] ),
    .A2(_0648_),
    .B1(_0737_),
    .C1(_0738_),
    .D1(_0739_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0740_));
 sky130_fd_sc_hd__nand2_1 _3889_ (.A(net20),
    .B(_0740_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0741_));
 sky130_fd_sc_hd__mux2_4 _3890_ (.A0(_0729_),
    .A1(_0741_),
    .S(_0654_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0742_));
 sky130_fd_sc_hd__a21o_1 _3891_ (.A1(_0721_),
    .A2(_0722_),
    .B1(_0742_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0743_));
 sky130_fd_sc_hd__nor2_4 _3892_ (.A(_0688_),
    .B(_0612_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0744_));
 sky130_fd_sc_hd__mux2_1 _3893_ (.A0(\i_tinyqv.cpu.i_core.cy ),
    .A1(_0658_),
    .S(_0744_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0745_));
 sky130_fd_sc_hd__and3_1 _3894_ (.A(_0742_),
    .B(_0721_),
    .C(_0722_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0746_));
 sky130_fd_sc_hd__a21o_1 _3895_ (.A1(_0743_),
    .A2(_0745_),
    .B1(_0746_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0747_));
 sky130_fd_sc_hd__buf_4 _3896_ (.A(_0619_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0748_));
 sky130_fd_sc_hd__clkbuf_4 _3897_ (.A(\i_tinyqv.cpu.pc[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0749_));
 sky130_fd_sc_hd__a22o_1 _3898_ (.A1(_0749_),
    .A2(_0615_),
    .B1(_0617_),
    .B2(\i_tinyqv.cpu.instr_data_start[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0750_));
 sky130_fd_sc_hd__a221o_1 _3899_ (.A1(\i_tinyqv.cpu.instr_data_start[5] ),
    .A2(_0748_),
    .B1(_0690_),
    .B2(\i_tinyqv.cpu.instr_data_start[9] ),
    .C1(_0750_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0751_));
 sky130_fd_sc_hd__buf_4 _3900_ (.A(_0611_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0752_));
 sky130_fd_sc_hd__a22o_1 _3901_ (.A1(\i_tinyqv.cpu.instr_data_start[21] ),
    .A2(_0610_),
    .B1(_0751_),
    .B2(_0752_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0753_));
 sky130_fd_sc_hd__a21oi_1 _3902_ (.A1(\i_tinyqv.cpu.instr_data_start[17] ),
    .A2(_0613_),
    .B1(_0753_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0754_));
 sky130_fd_sc_hd__a22o_1 _3903_ (.A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[12][1] ),
    .A2(net75),
    .B1(net46),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[14][1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0755_));
 sky130_fd_sc_hd__a221o_1 _3904_ (.A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[2][1] ),
    .A2(net26),
    .B1(_0646_),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[10][1] ),
    .C1(_0755_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0756_));
 sky130_fd_sc_hd__a221o_1 _3905_ (.A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[8][1] ),
    .A2(net27),
    .B1(_0648_),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[1][1] ),
    .C1(_0756_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0757_));
 sky130_fd_sc_hd__a22o_1 _3906_ (.A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[5][1] ),
    .A2(net57),
    .B1(_0639_),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[6][1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0758_));
 sky130_fd_sc_hd__a22o_1 _3907_ (.A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[7][1] ),
    .A2(net88),
    .B1(_0637_),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[11][1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0759_));
 sky130_fd_sc_hd__a221o_1 _3908_ (.A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[15][1] ),
    .A2(net83),
    .B1(net54),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[9][1] ),
    .C1(_0759_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0760_));
 sky130_fd_sc_hd__a211o_1 _3909_ (.A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[13][1] ),
    .A2(net63),
    .B1(_0758_),
    .C1(_0760_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0761_));
 sky130_fd_sc_hd__nor2_2 _3910_ (.A(_0757_),
    .B(_0761_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0762_));
 sky130_fd_sc_hd__mux2_2 _3911_ (.A0(_0754_),
    .A1(_0762_),
    .S(_0654_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0763_));
 sky130_fd_sc_hd__a22o_1 _3912_ (.A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[8][1] ),
    .A2(_0671_),
    .B1(_0674_),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[12][1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0764_));
 sky130_fd_sc_hd__a22o_1 _3913_ (.A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[15][1] ),
    .A2(_0677_),
    .B1(_0680_),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[9][1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0765_));
 sky130_fd_sc_hd__a211o_1 _3914_ (.A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[14][1] ),
    .A2(net61),
    .B1(_0764_),
    .C1(_0765_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0766_));
 sky130_fd_sc_hd__and3_1 _3915_ (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[2][1] ),
    .B(_0667_),
    .C(_0670_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0767_));
 sky130_fd_sc_hd__a221o_1 _3916_ (.A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[11][1] ),
    .A2(_0664_),
    .B1(_0681_),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[6][1] ),
    .C1(_0767_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0768_));
 sky130_fd_sc_hd__a22o_1 _3917_ (.A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[7][1] ),
    .A2(_0678_),
    .B1(net320),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[1][1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0769_));
 sky130_fd_sc_hd__a22o_1 _3918_ (.A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[5][1] ),
    .A2(_0675_),
    .B1(_0684_),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[13][1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0770_));
 sky130_fd_sc_hd__a311o_1 _3919_ (.A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[10][1] ),
    .A2(_0666_),
    .A3(_0667_),
    .B1(_0769_),
    .C1(_0770_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0771_));
 sky130_fd_sc_hd__nor3_4 _3920_ (.A(_0766_),
    .B(_0768_),
    .C(_0771_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0772_));
 sky130_fd_sc_hd__mux4_1 _3921_ (.A0(\i_tinyqv.cpu.imm[17] ),
    .A1(\i_tinyqv.cpu.imm[21] ),
    .A2(\i_tinyqv.cpu.imm[25] ),
    .A3(\i_tinyqv.cpu.imm[29] ),
    .S0(_0608_),
    .S1(_0614_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0773_));
 sky130_fd_sc_hd__a21o_1 _3922_ (.A1(\i_tinyqv.cpu.i_core.imm_lo[1] ),
    .A2(_0615_),
    .B1(\i_tinyqv.cpu.counter[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0774_));
 sky130_fd_sc_hd__and3_1 _3923_ (.A(_0614_),
    .B(_0608_),
    .C(\i_tinyqv.cpu.imm[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0775_));
 sky130_fd_sc_hd__a221o_1 _3924_ (.A1(\i_tinyqv.cpu.i_core.imm_lo[5] ),
    .A2(_0748_),
    .B1(_0690_),
    .B2(\i_tinyqv.cpu.i_core.imm_lo[9] ),
    .C1(_0775_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0776_));
 sky130_fd_sc_hd__o22a_2 _3925_ (.A1(_0611_),
    .A2(_0773_),
    .B1(_0774_),
    .B2(_0776_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0777_));
 sky130_fd_sc_hd__nand2_1 _3926_ (.A(_0698_),
    .B(_0777_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0778_));
 sky130_fd_sc_hd__o21a_1 _3927_ (.A1(_0698_),
    .A2(_0772_),
    .B1(_0778_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0779_));
 sky130_fd_sc_hd__xor2_1 _3928_ (.A(_0658_),
    .B(_0779_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0780_));
 sky130_fd_sc_hd__nand2_1 _3929_ (.A(_0763_),
    .B(_0780_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0781_));
 sky130_fd_sc_hd__nor2_1 _3930_ (.A(_0763_),
    .B(_0780_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0782_));
 sky130_fd_sc_hd__a21oi_2 _3931_ (.A1(_0747_),
    .A2(_0781_),
    .B1(_0782_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0783_));
 sky130_fd_sc_hd__clkbuf_4 _3932_ (.A(\i_tinyqv.cpu.instr_data_start[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0784_));
 sky130_fd_sc_hd__a22o_1 _3933_ (.A1(net85),
    .A2(_0615_),
    .B1(_0617_),
    .B2(\i_tinyqv.cpu.instr_data_start[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0785_));
 sky130_fd_sc_hd__a221o_1 _3934_ (.A1(\i_tinyqv.cpu.instr_data_start[6] ),
    .A2(_0619_),
    .B1(_0690_),
    .B2(\i_tinyqv.cpu.instr_data_start[10] ),
    .C1(_0785_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0786_));
 sky130_fd_sc_hd__a22o_1 _3935_ (.A1(\i_tinyqv.cpu.instr_data_start[22] ),
    .A2(_0610_),
    .B1(_0786_),
    .B2(_0752_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0787_));
 sky130_fd_sc_hd__a21oi_1 _3936_ (.A1(_0784_),
    .A2(_0613_),
    .B1(_0787_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0788_));
 sky130_fd_sc_hd__a22o_1 _3937_ (.A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[10][2] ),
    .A2(_0646_),
    .B1(_0637_),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[11][2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0789_));
 sky130_fd_sc_hd__a22o_1 _3938_ (.A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[6][2] ),
    .A2(_0639_),
    .B1(net62),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[13][2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0790_));
 sky130_fd_sc_hd__and4_1 _3939_ (.A(_0611_),
    .B(_0690_),
    .C(_0732_),
    .D(_0733_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0791_));
 sky130_fd_sc_hd__a22o_1 _3940_ (.A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[1][2] ),
    .A2(_0648_),
    .B1(net48),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[14][2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0792_));
 sky130_fd_sc_hd__or4_4 _3941_ (.A(_0789_),
    .B(_0790_),
    .C(_0791_),
    .D(_0792_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0793_));
 sky130_fd_sc_hd__a22o_1 _3942_ (.A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[8][2] ),
    .A2(net27),
    .B1(net26),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[2][2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0794_));
 sky130_fd_sc_hd__a22o_1 _3943_ (.A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[15][2] ),
    .A2(_0633_),
    .B1(_0631_),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[12][2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0795_));
 sky130_fd_sc_hd__a22o_1 _3944_ (.A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[5][2] ),
    .A2(_0645_),
    .B1(_0642_),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[9][2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0796_));
 sky130_fd_sc_hd__a2111o_2 _3945_ (.A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[7][2] ),
    .A2(_0649_),
    .B1(_0794_),
    .C1(_0795_),
    .D1(_0796_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0797_));
 sky130_fd_sc_hd__nor2_4 _3946_ (.A(_0793_),
    .B(_0797_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0798_));
 sky130_fd_sc_hd__mux2_1 _3947_ (.A0(_0788_),
    .A1(_0798_),
    .S(_0654_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0799_));
 sky130_fd_sc_hd__a22o_1 _3948_ (.A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[12][2] ),
    .A2(_0674_),
    .B1(_0678_),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[7][2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0800_));
 sky130_fd_sc_hd__a221o_1 _3949_ (.A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[15][2] ),
    .A2(_0677_),
    .B1(_0684_),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[13][2] ),
    .C1(_0800_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0801_));
 sky130_fd_sc_hd__a32o_1 _3950_ (.A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[2][2] ),
    .A2(_0667_),
    .A3(_0670_),
    .B1(net24),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[1][2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0802_));
 sky130_fd_sc_hd__a221o_1 _3951_ (.A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[11][2] ),
    .A2(_0664_),
    .B1(_0680_),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[9][2] ),
    .C1(_0802_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0803_));
 sky130_fd_sc_hd__and4_1 _3952_ (.A(_0611_),
    .B(_0620_),
    .C(_0711_),
    .D(_0670_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0804_));
 sky130_fd_sc_hd__a32o_1 _3953_ (.A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[10][2] ),
    .A2(_0666_),
    .A3(_0667_),
    .B1(_0681_),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[6][2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0805_));
 sky130_fd_sc_hd__a22o_1 _3954_ (.A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[8][2] ),
    .A2(net25),
    .B1(_0675_),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[5][2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0806_));
 sky130_fd_sc_hd__a2111o_1 _3955_ (.A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[14][2] ),
    .A2(_0668_),
    .B1(_0804_),
    .C1(_0805_),
    .D1(_0806_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0807_));
 sky130_fd_sc_hd__nor3_1 _3956_ (.A(_0801_),
    .B(_0803_),
    .C(_0807_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0808_));
 sky130_fd_sc_hd__a22o_1 _3957_ (.A1(\i_tinyqv.cpu.imm[22] ),
    .A2(_0619_),
    .B1(_0690_),
    .B2(\i_tinyqv.cpu.imm[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0809_));
 sky130_fd_sc_hd__a221o_1 _3958_ (.A1(\i_tinyqv.cpu.imm[18] ),
    .A2(_0615_),
    .B1(_0617_),
    .B2(\i_tinyqv.cpu.imm[30] ),
    .C1(_0809_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0810_));
 sky130_fd_sc_hd__a22o_1 _3959_ (.A1(\i_tinyqv.cpu.imm[14] ),
    .A2(_0617_),
    .B1(_0619_),
    .B2(\i_tinyqv.cpu.i_core.imm_lo[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0811_));
 sky130_fd_sc_hd__a221o_1 _3960_ (.A1(\i_tinyqv.cpu.i_core.imm_lo[2] ),
    .A2(_0615_),
    .B1(_0690_),
    .B2(\i_tinyqv.cpu.i_core.imm_lo[10] ),
    .C1(\i_tinyqv.cpu.counter[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0812_));
 sky130_fd_sc_hd__or2_1 _3961_ (.A(_0811_),
    .B(_0812_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0813_));
 sky130_fd_sc_hd__o21ai_2 _3962_ (.A1(_0752_),
    .A2(_0810_),
    .B1(_0813_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0814_));
 sky130_fd_sc_hd__mux2_1 _3963_ (.A0(net16),
    .A1(_0814_),
    .S(_0698_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0815_));
 sky130_fd_sc_hd__xor2_1 _3964_ (.A(_0658_),
    .B(_0815_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0816_));
 sky130_fd_sc_hd__or2_1 _3965_ (.A(net86),
    .B(_0816_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0817_));
 sky130_fd_sc_hd__nand2_1 _3966_ (.A(net86),
    .B(_0816_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0818_));
 sky130_fd_sc_hd__nand2_1 _3967_ (.A(_0817_),
    .B(_0818_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0819_));
 sky130_fd_sc_hd__nand2_1 _3968_ (.A(net80),
    .B(_0700_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0820_));
 sky130_fd_sc_hd__o211ai_2 _3969_ (.A1(_0783_),
    .A2(_0819_),
    .B1(_0820_),
    .C1(_0817_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0821_));
 sky130_fd_sc_hd__or2b_4 _3970_ (.A(_0655_),
    .B_N(_0699_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0822_));
 sky130_fd_sc_hd__or2b_1 _3971_ (.A(_0699_),
    .B_N(_0655_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0823_));
 sky130_fd_sc_hd__nand2_2 _3972_ (.A(_0822_),
    .B(_0823_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0824_));
 sky130_fd_sc_hd__a21oi_1 _3973_ (.A1(_0656_),
    .A2(_0824_),
    .B1(net141),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0825_));
 sky130_fd_sc_hd__a21o_1 _3974_ (.A1(_0701_),
    .A2(_0821_),
    .B1(_0825_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0826_));
 sky130_fd_sc_hd__and2_1 _3975_ (.A(_0799_),
    .B(_0815_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0827_));
 sky130_fd_sc_hd__nor2_1 _3976_ (.A(_0799_),
    .B(_0815_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0828_));
 sky130_fd_sc_hd__nor2_1 _3977_ (.A(_0708_),
    .B(net79),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0829_));
 sky130_fd_sc_hd__xor2_1 _3978_ (.A(_0742_),
    .B(_0829_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0830_));
 sky130_fd_sc_hd__xnor2_1 _3979_ (.A(_0763_),
    .B(_0779_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0831_));
 sky130_fd_sc_hd__o211a_1 _3980_ (.A1(_0827_),
    .A2(_0828_),
    .B1(_0830_),
    .C1(_0831_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0832_));
 sky130_fd_sc_hd__o21a_1 _3981_ (.A1(\i_tinyqv.cpu.i_core.cmp ),
    .A2(_0744_),
    .B1(_0824_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0833_));
 sky130_fd_sc_hd__a21oi_1 _3982_ (.A1(_0832_),
    .A2(_0833_),
    .B1(_0656_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0834_));
 sky130_fd_sc_hd__a211o_1 _3983_ (.A1(_0656_),
    .A2(_0820_),
    .B1(_0834_),
    .C1(net141),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0835_));
 sky130_fd_sc_hd__nand2_1 _3984_ (.A(_0826_),
    .B(_0835_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\i_tinyqv.cpu.i_core.cmp_out ));
 sky130_fd_sc_hd__nor2_1 _3985_ (.A(\i_tinyqv.cpu.is_store ),
    .B(\i_tinyqv.cpu.is_load ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0836_));
 sky130_fd_sc_hd__o21a_1 _3986_ (.A1(\i_tinyqv.cpu.no_write_in_progress ),
    .A2(_0836_),
    .B1(\i_tinyqv.cpu.debug_instr_valid ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0837_));
 sky130_fd_sc_hd__clkbuf_8 _3987_ (.A(_0608_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0838_));
 sky130_fd_sc_hd__and2_1 _3988_ (.A(\i_tinyqv.cpu.counter[4] ),
    .B(_0614_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0839_));
 sky130_fd_sc_hd__buf_2 _3989_ (.A(_0839_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0840_));
 sky130_fd_sc_hd__nand2_2 _3990_ (.A(_0838_),
    .B(_0840_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0841_));
 sky130_fd_sc_hd__inv_2 _3991_ (.A(\i_tinyqv.cpu.i_core.cycle[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0842_));
 sky130_fd_sc_hd__inv_2 _3992_ (.A(\i_tinyqv.cpu.alu_op[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0843_));
 sky130_fd_sc_hd__inv_2 _3993_ (.A(\i_tinyqv.cpu.alu_op[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0844_));
 sky130_fd_sc_hd__and2_1 _3994_ (.A(_0844_),
    .B(\i_tinyqv.cpu.alu_op[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0845_));
 sky130_fd_sc_hd__and2_2 _3995_ (.A(\i_tinyqv.cpu.alu_op[1] ),
    .B(\i_tinyqv.cpu.alu_op[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0846_));
 sky130_fd_sc_hd__a211o_2 _3996_ (.A1(_0843_),
    .A2(\i_tinyqv.cpu.alu_op[1] ),
    .B1(_0845_),
    .C1(_0846_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0847_));
 sky130_fd_sc_hd__nor2_1 _3997_ (.A(_0842_),
    .B(_0847_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0848_));
 sky130_fd_sc_hd__o21ai_2 _3998_ (.A1(\i_tinyqv.cpu.is_alu_reg ),
    .A2(\i_tinyqv.cpu.is_alu_imm ),
    .B1(_0653_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0849_));
 sky130_fd_sc_hd__a211o_1 _3999_ (.A1(_0842_),
    .A2(_0847_),
    .B1(_0849_),
    .C1(\i_tinyqv.cpu.i_core.cycle[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0850_));
 sky130_fd_sc_hd__and3_1 _4000_ (.A(\i_tinyqv.cpu.debug_instr_valid ),
    .B(\i_tinyqv.cpu.is_load ),
    .C(\i_tinyqv.cpu.no_write_in_progress ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0851_));
 sky130_fd_sc_hd__nand2_1 _4001_ (.A(\i_tinyqv.cpu.debug_instr_valid ),
    .B(\i_tinyqv.cpu.is_auipc ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0852_));
 sky130_fd_sc_hd__nor2_1 _4002_ (.A(\i_tinyqv.cpu.i_core.is_interrupt ),
    .B(\i_tinyqv.cpu.is_branch ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0853_));
 sky130_fd_sc_hd__nand2_4 _4003_ (.A(\i_tinyqv.cpu.is_store ),
    .B(\i_tinyqv.cpu.no_write_in_progress ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0854_));
 sky130_fd_sc_hd__nand2_2 _4004_ (.A(\i_tinyqv.cpu.debug_instr_valid ),
    .B(\i_tinyqv.cpu.is_system ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0855_));
 sky130_fd_sc_hd__and4_1 _4005_ (.A(_0852_),
    .B(_0853_),
    .C(_0854_),
    .D(_0855_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0856_));
 sky130_fd_sc_hd__nand2_1 _4006_ (.A(\i_tinyqv.cpu.debug_instr_valid ),
    .B(\i_tinyqv.cpu.is_lui ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0857_));
 sky130_fd_sc_hd__o21ai_4 _4007_ (.A1(\i_tinyqv.cpu.is_jal ),
    .A2(\i_tinyqv.cpu.is_jalr ),
    .B1(\i_tinyqv.cpu.debug_instr_valid ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0858_));
 sky130_fd_sc_hd__nand4_1 _4008_ (.A(_0837_),
    .B(_0856_),
    .C(_0857_),
    .D(_0858_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0859_));
 sky130_fd_sc_hd__a31o_1 _4009_ (.A1(\i_tinyqv.cpu.i_core.load_done ),
    .A2(_0849_),
    .A3(_0851_),
    .B1(_0859_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0860_));
 sky130_fd_sc_hd__o21ba_1 _4010_ (.A1(_0848_),
    .A2(_0850_),
    .B1_N(_0860_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0861_));
 sky130_fd_sc_hd__or2_1 _4011_ (.A(_0841_),
    .B(_0861_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0862_));
 sky130_fd_sc_hd__inv_2 _4012_ (.A(_0862_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0863_));
 sky130_fd_sc_hd__o21a_1 _4013_ (.A1(net127),
    .A2(_0837_),
    .B1(_0863_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0029_));
 sky130_fd_sc_hd__inv_2 _4014_ (.A(\i_tinyqv.mem.qspi_data_byte_idx[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0864_));
 sky130_fd_sc_hd__or3_4 _4015_ (.A(\i_tinyqv.cpu.data_addr[27] ),
    .B(\i_tinyqv.cpu.data_addr[26] ),
    .C(\i_tinyqv.cpu.data_addr[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0865_));
 sky130_fd_sc_hd__a21o_1 _4016_ (.A1(\i_tinyqv.cpu.data_read_n[1] ),
    .A2(\i_tinyqv.cpu.data_write_n[1] ),
    .B1(_0865_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0866_));
 sky130_fd_sc_hd__xnor2_1 _4017_ (.A(_0864_),
    .B(_0866_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0867_));
 sky130_fd_sc_hd__clkbuf_4 _4018_ (.A(\i_tinyqv.mem.qspi_data_byte_idx[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0868_));
 sky130_fd_sc_hd__a21oi_2 _4019_ (.A1(\i_tinyqv.cpu.data_read_n[0] ),
    .A2(\i_tinyqv.cpu.data_write_n[0] ),
    .B1(_0866_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0869_));
 sky130_fd_sc_hd__and2_1 _4020_ (.A(_0868_),
    .B(_0869_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0870_));
 sky130_fd_sc_hd__nor2_1 _4021_ (.A(_0868_),
    .B(_0869_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0871_));
 sky130_fd_sc_hd__nor3_1 _4022_ (.A(_0867_),
    .B(_0870_),
    .C(_0871_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0872_));
 sky130_fd_sc_hd__and2_1 _4023_ (.A(\i_tinyqv.mem.q_ctrl.data_req ),
    .B(_0872_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0873_));
 sky130_fd_sc_hd__clkbuf_1 _4024_ (.A(_0873_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0082_));
 sky130_fd_sc_hd__mux2_1 _4025_ (.A0(\i_uart_tx.txd_reg ),
    .A1(\gpio_out[0] ),
    .S(\gpio_out_sel[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0874_));
 sky130_fd_sc_hd__buf_4 _4026_ (.A(_0874_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[0]));
 sky130_fd_sc_hd__mux2_2 _4027_ (.A0(\i_spi.spi_select ),
    .A1(\debug_rd_r[2] ),
    .S(debug_register_data),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0875_));
 sky130_fd_sc_hd__mux2_1 _4028_ (.A0(_0875_),
    .A1(\gpio_out[4] ),
    .S(\gpio_out_sel[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0876_));
 sky130_fd_sc_hd__clkbuf_4 _4029_ (.A(_0876_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[4]));
 sky130_fd_sc_hd__and2_2 _4030_ (.A(_0852_),
    .B(_0849_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0877_));
 sky130_fd_sc_hd__nand2_2 _4031_ (.A(\i_tinyqv.cpu.data_ready_core ),
    .B(_0851_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0878_));
 sky130_fd_sc_hd__and2_1 _4032_ (.A(_0653_),
    .B(\i_tinyqv.cpu.is_lui ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0879_));
 sky130_fd_sc_hd__clkbuf_2 _4033_ (.A(_0879_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0880_));
 sky130_fd_sc_hd__buf_2 _4034_ (.A(\i_tinyqv.cpu.instr_data_start[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0881_));
 sky130_fd_sc_hd__buf_2 _4035_ (.A(\i_tinyqv.cpu.instr_data_start[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0882_));
 sky130_fd_sc_hd__buf_2 _4036_ (.A(\i_tinyqv.cpu.instr_data_start[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0883_));
 sky130_fd_sc_hd__buf_2 _4037_ (.A(\i_tinyqv.cpu.instr_data_start[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0884_));
 sky130_fd_sc_hd__and2_1 _4038_ (.A(\i_tinyqv.cpu.instr_len[2] ),
    .B(\i_tinyqv.cpu.pc[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0885_));
 sky130_fd_sc_hd__nor2_1 _4039_ (.A(\i_tinyqv.cpu.instr_len[2] ),
    .B(\i_tinyqv.cpu.pc[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0886_));
 sky130_fd_sc_hd__nor2_4 _4040_ (.A(_0885_),
    .B(_0886_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0887_));
 sky130_fd_sc_hd__a31o_2 _4041_ (.A1(\i_tinyqv.cpu.instr_len[1] ),
    .A2(_0749_),
    .A3(_0887_),
    .B1(_0885_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0888_));
 sky130_fd_sc_hd__and3_1 _4042_ (.A(\i_tinyqv.cpu.instr_data_start[4] ),
    .B(_0884_),
    .C(_0888_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0889_));
 sky130_fd_sc_hd__and2_1 _4043_ (.A(\i_tinyqv.cpu.instr_data_start[5] ),
    .B(_0889_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0890_));
 sky130_fd_sc_hd__and3_1 _4044_ (.A(\i_tinyqv.cpu.instr_data_start[7] ),
    .B(_0883_),
    .C(_0890_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0891_));
 sky130_fd_sc_hd__and2_1 _4045_ (.A(\i_tinyqv.cpu.instr_data_start[8] ),
    .B(_0891_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0892_));
 sky130_fd_sc_hd__and3_1 _4046_ (.A(\i_tinyqv.cpu.instr_data_start[10] ),
    .B(_0882_),
    .C(_0892_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0893_));
 sky130_fd_sc_hd__and2_1 _4047_ (.A(\i_tinyqv.cpu.instr_data_start[11] ),
    .B(_0893_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0894_));
 sky130_fd_sc_hd__and3_1 _4048_ (.A(\i_tinyqv.cpu.instr_data_start[13] ),
    .B(_0726_),
    .C(_0894_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0895_));
 sky130_fd_sc_hd__and2_1 _4049_ (.A(\i_tinyqv.cpu.instr_data_start[14] ),
    .B(_0895_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0896_));
 sky130_fd_sc_hd__and3_1 _4050_ (.A(\i_tinyqv.cpu.instr_data_start[16] ),
    .B(_0881_),
    .C(_0896_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0897_));
 sky130_fd_sc_hd__and2_1 _4051_ (.A(\i_tinyqv.cpu.instr_data_start[17] ),
    .B(_0897_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0898_));
 sky130_fd_sc_hd__and3_1 _4052_ (.A(\i_tinyqv.cpu.instr_data_start[19] ),
    .B(_0784_),
    .C(_0898_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0899_));
 sky130_fd_sc_hd__and2_1 _4053_ (.A(\i_tinyqv.cpu.instr_data_start[20] ),
    .B(_0899_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0900_));
 sky130_fd_sc_hd__nor2_1 _4054_ (.A(\i_tinyqv.cpu.instr_data_start[20] ),
    .B(_0899_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0901_));
 sky130_fd_sc_hd__nor2_1 _4055_ (.A(_0900_),
    .B(_0901_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0902_));
 sky130_fd_sc_hd__nand2_1 _4056_ (.A(_0610_),
    .B(_0902_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0903_));
 sky130_fd_sc_hd__a21oi_1 _4057_ (.A1(_0884_),
    .A2(_0888_),
    .B1(\i_tinyqv.cpu.instr_data_start[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0904_));
 sky130_fd_sc_hd__or2_1 _4058_ (.A(_0889_),
    .B(_0904_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0905_));
 sky130_fd_sc_hd__xnor2_1 _4059_ (.A(_0726_),
    .B(_0894_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0906_));
 sky130_fd_sc_hd__clkbuf_8 _4060_ (.A(_0614_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0907_));
 sky130_fd_sc_hd__clkinv_4 _4061_ (.A(_0838_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0908_));
 sky130_fd_sc_hd__nand2_4 _4062_ (.A(_0907_),
    .B(_0908_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0909_));
 sky130_fd_sc_hd__nor2_1 _4063_ (.A(\i_tinyqv.cpu.instr_data_start[8] ),
    .B(_0891_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0910_));
 sky130_fd_sc_hd__or2_1 _4064_ (.A(_0892_),
    .B(_0910_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0911_));
 sky130_fd_sc_hd__or2_1 _4065_ (.A(_0909_),
    .B(_0911_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0912_));
 sky130_fd_sc_hd__o221a_1 _4066_ (.A1(_0609_),
    .A2(_0905_),
    .B1(_0906_),
    .B2(_0724_),
    .C1(_0912_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0913_));
 sky130_fd_sc_hd__a21oi_1 _4067_ (.A1(_0881_),
    .A2(_0896_),
    .B1(\i_tinyqv.cpu.instr_data_start[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0914_));
 sky130_fd_sc_hd__or2_1 _4068_ (.A(_0897_),
    .B(_0914_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0915_));
 sky130_fd_sc_hd__nand2_4 _4069_ (.A(_0688_),
    .B(_0689_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0916_));
 sky130_fd_sc_hd__o22a_1 _4070_ (.A1(_0688_),
    .A2(_0913_),
    .B1(_0915_),
    .B2(_0916_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0917_));
 sky130_fd_sc_hd__a21o_1 _4071_ (.A1(_0903_),
    .A2(_0917_),
    .B1(_0858_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0918_));
 sky130_fd_sc_hd__nor2_2 _4072_ (.A(_0656_),
    .B(\i_tinyqv.cpu.alu_op[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0919_));
 sky130_fd_sc_hd__nor2_2 _4073_ (.A(_0855_),
    .B(_0919_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0920_));
 sky130_fd_sc_hd__and2_1 _4074_ (.A(_0858_),
    .B(_0920_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0921_));
 sky130_fd_sc_hd__or4b_2 _4075_ (.A(\i_tinyqv.cpu.i_core.imm_lo[3] ),
    .B(\i_tinyqv.cpu.i_core.imm_lo[2] ),
    .C(\i_tinyqv.cpu.i_core.imm_lo[1] ),
    .D_N(\i_tinyqv.cpu.i_core.imm_lo[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0922_));
 sky130_fd_sc_hd__or3_1 _4076_ (.A(\i_tinyqv.cpu.i_core.imm_lo[7] ),
    .B(\i_tinyqv.cpu.i_core.imm_lo[5] ),
    .C(\i_tinyqv.cpu.i_core.imm_lo[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0923_));
 sky130_fd_sc_hd__or2_1 _4077_ (.A(\i_tinyqv.cpu.i_core.imm_lo[8] ),
    .B(\i_tinyqv.cpu.i_core.imm_lo[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0924_));
 sky130_fd_sc_hd__nand2_1 _4078_ (.A(\i_tinyqv.cpu.i_core.imm_lo[11] ),
    .B(\i_tinyqv.cpu.i_core.imm_lo[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0925_));
 sky130_fd_sc_hd__or4_1 _4079_ (.A(\i_tinyqv.cpu.i_core.imm_lo[6] ),
    .B(_0923_),
    .C(_0924_),
    .D(_0925_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0926_));
 sky130_fd_sc_hd__nor2_1 _4080_ (.A(_0922_),
    .B(_0926_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0927_));
 sky130_fd_sc_hd__or4b_1 _4081_ (.A(\i_tinyqv.cpu.i_core.imm_lo[3] ),
    .B(\i_tinyqv.cpu.i_core.imm_lo[2] ),
    .C(\i_tinyqv.cpu.i_core.imm_lo[0] ),
    .D_N(\i_tinyqv.cpu.i_core.imm_lo[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0928_));
 sky130_fd_sc_hd__nor2_1 _4082_ (.A(_0928_),
    .B(_0926_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0929_));
 sky130_fd_sc_hd__or4_1 _4083_ (.A(\i_tinyqv.cpu.i_core.imm_lo[3] ),
    .B(\i_tinyqv.cpu.i_core.imm_lo[2] ),
    .C(\i_tinyqv.cpu.i_core.imm_lo[1] ),
    .D(\i_tinyqv.cpu.i_core.imm_lo[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0930_));
 sky130_fd_sc_hd__nor2_1 _4084_ (.A(_0926_),
    .B(_0930_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0931_));
 sky130_fd_sc_hd__and4bb_1 _4085_ (.A_N(\i_tinyqv.cpu.i_core.imm_lo[11] ),
    .B_N(\i_tinyqv.cpu.i_core.imm_lo[10] ),
    .C(\i_tinyqv.cpu.i_core.imm_lo[8] ),
    .D(\i_tinyqv.cpu.i_core.imm_lo[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0932_));
 sky130_fd_sc_hd__or3b_2 _4086_ (.A(\i_tinyqv.cpu.i_core.imm_lo[6] ),
    .B(_0923_),
    .C_N(_0932_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0933_));
 sky130_fd_sc_hd__or2_1 _4087_ (.A(_0933_),
    .B(_0922_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0934_));
 sky130_fd_sc_hd__inv_2 _4088_ (.A(\i_tinyqv.cpu.i_core.mcause[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0935_));
 sky130_fd_sc_hd__nor3_1 _4089_ (.A(\i_tinyqv.cpu.i_core.imm_lo[7] ),
    .B(\i_tinyqv.cpu.i_core.imm_lo[5] ),
    .C(\i_tinyqv.cpu.i_core.imm_lo[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0936_));
 sky130_fd_sc_hd__nand3_2 _4090_ (.A(\i_tinyqv.cpu.i_core.imm_lo[6] ),
    .B(_0936_),
    .C(_0932_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0937_));
 sky130_fd_sc_hd__or3_1 _4091_ (.A(_0935_),
    .B(_0928_),
    .C(_0937_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0938_));
 sky130_fd_sc_hd__nand2_4 _4092_ (.A(_0752_),
    .B(_0748_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0939_));
 sky130_fd_sc_hd__a21oi_1 _4093_ (.A1(_0934_),
    .A2(_0938_),
    .B1(_0939_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0940_));
 sky130_fd_sc_hd__a221o_1 _4094_ (.A1(\i_tinyqv.cpu.i_core.i_instrret.data[0] ),
    .A2(_0929_),
    .B1(_0931_),
    .B2(\i_tinyqv.cpu.i_core.cycle_count[0] ),
    .C1(_0940_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0941_));
 sky130_fd_sc_hd__or4b_4 _4095_ (.A(\i_tinyqv.cpu.i_core.imm_lo[3] ),
    .B(\i_tinyqv.cpu.i_core.imm_lo[1] ),
    .C(\i_tinyqv.cpu.i_core.imm_lo[0] ),
    .D_N(\i_tinyqv.cpu.i_core.imm_lo[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0942_));
 sky130_fd_sc_hd__nor3_1 _4096_ (.A(_0916_),
    .B(_0937_),
    .C(_0942_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0943_));
 sky130_fd_sc_hd__nor3_4 _4097_ (.A(_0916_),
    .B(_0942_),
    .C(_0933_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0944_));
 sky130_fd_sc_hd__nor2_2 _4098_ (.A(_0688_),
    .B(_0907_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0945_));
 sky130_fd_sc_hd__nand2_2 _4099_ (.A(_0908_),
    .B(_0945_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0946_));
 sky130_fd_sc_hd__nor3_1 _4100_ (.A(_0946_),
    .B(_0928_),
    .C(_0937_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0947_));
 sky130_fd_sc_hd__nor3_1 _4101_ (.A(_0840_),
    .B(_0937_),
    .C(_0922_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0948_));
 sky130_fd_sc_hd__a22o_1 _4102_ (.A1(\i_tinyqv.cpu.i_core.mcause[0] ),
    .A2(_0947_),
    .B1(_0948_),
    .B2(\i_tinyqv.cpu.i_core.mepc[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0949_));
 sky130_fd_sc_hd__a221o_1 _4103_ (.A1(\i_tinyqv.cpu.i_core.mip[16] ),
    .A2(_0943_),
    .B1(_0944_),
    .B2(\i_tinyqv.cpu.i_core.mie[16] ),
    .C1(_0949_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0950_));
 sky130_fd_sc_hd__a211o_1 _4104_ (.A1(\i_tinyqv.cpu.i_core.cycle_count[3] ),
    .A2(_0927_),
    .B1(_0941_),
    .C1(_0950_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0951_));
 sky130_fd_sc_hd__a21oi_1 _4105_ (.A1(_0921_),
    .A2(_0951_),
    .B1(_0880_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0952_));
 sky130_fd_sc_hd__a22o_1 _4106_ (.A1(_0707_),
    .A2(_0880_),
    .B1(_0918_),
    .B2(_0952_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0953_));
 sky130_fd_sc_hd__nand2_1 _4107_ (.A(_0878_),
    .B(_0953_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0954_));
 sky130_fd_sc_hd__a211o_2 _4108_ (.A1(\i_tinyqv.cpu.i_core.mem_op[0] ),
    .A2(_0752_),
    .B1(_0945_),
    .C1(\i_tinyqv.cpu.i_core.mem_op[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0955_));
 sky130_fd_sc_hd__buf_2 _4109_ (.A(_0688_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0956_));
 sky130_fd_sc_hd__clkbuf_4 _4110_ (.A(_0865_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0957_));
 sky130_fd_sc_hd__a221o_1 _4111_ (.A1(\i_tinyqv.mem.data_from_read[16] ),
    .A2(_0689_),
    .B1(_0748_),
    .B2(\i_tinyqv.mem.data_from_read[20] ),
    .C1(_0957_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0958_));
 sky130_fd_sc_hd__or4_1 _4112_ (.A(\i_tinyqv.cpu.data_addr[24] ),
    .B(\i_tinyqv.cpu.data_addr[1] ),
    .C(\i_tinyqv.cpu.data_addr[7] ),
    .D(\i_tinyqv.cpu.data_addr[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0959_));
 sky130_fd_sc_hd__or4b_1 _4113_ (.A(\i_tinyqv.cpu.data_addr[0] ),
    .B(\i_tinyqv.cpu.data_addr[26] ),
    .C(\i_tinyqv.cpu.data_addr[25] ),
    .D_N(\i_tinyqv.cpu.data_addr[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0960_));
 sky130_fd_sc_hd__or2_1 _4114_ (.A(_0959_),
    .B(_0960_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0961_));
 sky130_fd_sc_hd__or4_1 _4115_ (.A(\i_tinyqv.cpu.data_addr[13] ),
    .B(\i_tinyqv.cpu.data_addr[12] ),
    .C(\i_tinyqv.cpu.data_addr[15] ),
    .D(\i_tinyqv.cpu.data_addr[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0962_));
 sky130_fd_sc_hd__or4_1 _4116_ (.A(\i_tinyqv.cpu.data_addr[9] ),
    .B(\i_tinyqv.cpu.data_addr[8] ),
    .C(\i_tinyqv.cpu.data_addr[11] ),
    .D(\i_tinyqv.cpu.data_addr[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0963_));
 sky130_fd_sc_hd__or4_1 _4117_ (.A(\i_tinyqv.cpu.data_addr[21] ),
    .B(\i_tinyqv.cpu.data_addr[20] ),
    .C(\i_tinyqv.cpu.data_addr[23] ),
    .D(\i_tinyqv.cpu.data_addr[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0964_));
 sky130_fd_sc_hd__or4_1 _4118_ (.A(\i_tinyqv.cpu.data_addr[17] ),
    .B(\i_tinyqv.cpu.data_addr[16] ),
    .C(\i_tinyqv.cpu.data_addr[19] ),
    .D(\i_tinyqv.cpu.data_addr[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0965_));
 sky130_fd_sc_hd__or4_2 _4119_ (.A(_0962_),
    .B(_0963_),
    .C(_0964_),
    .D(_0965_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0966_));
 sky130_fd_sc_hd__nor3_1 _4120_ (.A(\i_tinyqv.cpu.data_addr[5] ),
    .B(_0961_),
    .C(_0966_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0967_));
 sky130_fd_sc_hd__nand2_1 _4121_ (.A(\i_tinyqv.cpu.data_addr[2] ),
    .B(_0967_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0968_));
 sky130_fd_sc_hd__or3_4 _4122_ (.A(\i_tinyqv.cpu.data_addr[3] ),
    .B(_0961_),
    .C(_0966_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0969_));
 sky130_fd_sc_hd__and2b_1 _4123_ (.A_N(_0967_),
    .B(\i_tinyqv.cpu.data_addr[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0970_));
 sky130_fd_sc_hd__a21o_2 _4124_ (.A1(_0968_),
    .A2(_0969_),
    .B1(_0970_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0971_));
 sky130_fd_sc_hd__nor3_1 _4125_ (.A(\i_tinyqv.cpu.data_addr[27] ),
    .B(\i_tinyqv.cpu.data_addr[26] ),
    .C(\i_tinyqv.cpu.data_addr[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0972_));
 sky130_fd_sc_hd__and2_1 _4126_ (.A(_0907_),
    .B(net28),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0973_));
 sky130_fd_sc_hd__buf_4 _4127_ (.A(_0838_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0974_));
 sky130_fd_sc_hd__mux2_1 _4128_ (.A0(\i_tinyqv.mem.qspi_data_buf[24] ),
    .A1(\i_tinyqv.mem.qspi_data_buf[28] ),
    .S(_0974_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0975_));
 sky130_fd_sc_hd__mux2_1 _4129_ (.A0(\i_tinyqv.cpu.instr_data_in[8] ),
    .A1(\i_tinyqv.cpu.instr_data_in[12] ),
    .S(_0838_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0976_));
 sky130_fd_sc_hd__and2_1 _4130_ (.A(\i_tinyqv.mem.q_ctrl.data_ready ),
    .B(_0872_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0977_));
 sky130_fd_sc_hd__inv_2 _4131_ (.A(\i_tinyqv.mem.instr_active ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0978_));
 sky130_fd_sc_hd__o21a_4 _4132_ (.A1(\i_tinyqv.mem.qspi_write_done ),
    .A2(_0977_),
    .B1(_0978_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0979_));
 sky130_fd_sc_hd__mux2_1 _4133_ (.A0(_0975_),
    .A1(_0976_),
    .S(_0979_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0980_));
 sky130_fd_sc_hd__a22o_1 _4134_ (.A1(_0958_),
    .A2(_0971_),
    .B1(_0973_),
    .B2(_0980_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0981_));
 sky130_fd_sc_hd__and2_1 _4135_ (.A(_0752_),
    .B(_0971_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0982_));
 sky130_fd_sc_hd__or4_4 _4136_ (.A(\i_tinyqv.cpu.data_addr[4] ),
    .B(\i_tinyqv.cpu.data_addr[5] ),
    .C(_0961_),
    .D(_0966_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0983_));
 sky130_fd_sc_hd__inv_2 _4137_ (.A(\i_tinyqv.cpu.data_addr[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0984_));
 sky130_fd_sc_hd__or2_2 _4138_ (.A(_0984_),
    .B(_0969_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0985_));
 sky130_fd_sc_hd__nor2_2 _4139_ (.A(_0983_),
    .B(_0985_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0986_));
 sky130_fd_sc_hd__and2_1 _4140_ (.A(\i_tinyqv.cpu.data_addr[4] ),
    .B(_0967_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0987_));
 sky130_fd_sc_hd__or3_2 _4141_ (.A(\i_debug_uart_tx.fsm_state[3] ),
    .B(\i_debug_uart_tx.fsm_state[2] ),
    .C(\i_debug_uart_tx.fsm_state[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0988_));
 sky130_fd_sc_hd__or2_4 _4142_ (.A(\i_debug_uart_tx.fsm_state[0] ),
    .B(_0988_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0989_));
 sky130_fd_sc_hd__or3_4 _4143_ (.A(\i_uart_tx.fsm_state[3] ),
    .B(\i_uart_tx.fsm_state[2] ),
    .C(\i_uart_tx.fsm_state[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0990_));
 sky130_fd_sc_hd__nor2_4 _4144_ (.A(\i_uart_tx.fsm_state[0] ),
    .B(_0990_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0991_));
 sky130_fd_sc_hd__nor2_1 _4145_ (.A(_0985_),
    .B(_0991_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0992_));
 sky130_fd_sc_hd__a31o_1 _4146_ (.A1(\i_tinyqv.cpu.data_addr[2] ),
    .A2(_0969_),
    .A3(_0989_),
    .B1(_0992_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0993_));
 sky130_fd_sc_hd__a221o_1 _4147_ (.A1(net2),
    .A2(_0986_),
    .B1(_0987_),
    .B2(_0993_),
    .C1(_0974_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0994_));
 sky130_fd_sc_hd__inv_2 _4148_ (.A(_0969_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0995_));
 sky130_fd_sc_hd__and3_1 _4149_ (.A(_0984_),
    .B(_0995_),
    .C(_0987_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0996_));
 sky130_fd_sc_hd__clkbuf_4 _4150_ (.A(_0996_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0997_));
 sky130_fd_sc_hd__or2_2 _4151_ (.A(\i_tinyqv.cpu.data_addr[4] ),
    .B(_0967_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0998_));
 sky130_fd_sc_hd__or2_2 _4152_ (.A(\i_tinyqv.cpu.data_addr[2] ),
    .B(_0969_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0999_));
 sky130_fd_sc_hd__nor2_4 _4153_ (.A(_0998_),
    .B(_0999_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1000_));
 sky130_fd_sc_hd__nor2_4 _4154_ (.A(_0999_),
    .B(_0983_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1001_));
 sky130_fd_sc_hd__a22o_1 _4155_ (.A1(\i_spi.data[0] ),
    .A2(_1000_),
    .B1(_1001_),
    .B2(uo_out[0]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1002_));
 sky130_fd_sc_hd__nor3_1 _4156_ (.A(_0984_),
    .B(_0995_),
    .C(_0983_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1003_));
 sky130_fd_sc_hd__nor2_2 _4157_ (.A(_0998_),
    .B(_0985_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1004_));
 sky130_fd_sc_hd__a22o_1 _4158_ (.A1(\gpio_out_sel[0] ),
    .A2(_1003_),
    .B1(_1004_),
    .B2(\i_spi.busy ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1005_));
 sky130_fd_sc_hd__a211o_1 _4159_ (.A1(\i_uart_rx.recieved_data[0] ),
    .A2(_0997_),
    .B1(_1002_),
    .C1(_1005_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1006_));
 sky130_fd_sc_hd__a221o_1 _4160_ (.A1(net6),
    .A2(_0986_),
    .B1(_0997_),
    .B2(\i_uart_rx.recieved_data[4] ),
    .C1(_0908_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1007_));
 sky130_fd_sc_hd__a22o_1 _4161_ (.A1(\i_spi.data[4] ),
    .A2(_1000_),
    .B1(_1001_),
    .B2(uo_out[4]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1008_));
 sky130_fd_sc_hd__a211o_1 _4162_ (.A1(\gpio_out_sel[4] ),
    .A2(net14),
    .B1(_1007_),
    .C1(_1008_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1009_));
 sky130_fd_sc_hd__o211a_1 _4163_ (.A1(_0994_),
    .A2(_1006_),
    .B1(_1009_),
    .C1(_0945_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1010_));
 sky130_fd_sc_hd__mux2_1 _4164_ (.A0(\i_tinyqv.cpu.instr_data_in[0] ),
    .A1(\i_tinyqv.cpu.instr_data_in[4] ),
    .S(_0974_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1011_));
 sky130_fd_sc_hd__nand2_2 _4165_ (.A(_0869_),
    .B(_0979_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1012_));
 sky130_fd_sc_hd__mux2_1 _4166_ (.A0(_0976_),
    .A1(_1011_),
    .S(_1012_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1013_));
 sky130_fd_sc_hd__mux2_1 _4167_ (.A0(\i_tinyqv.mem.qspi_data_buf[8] ),
    .A1(\i_tinyqv.mem.qspi_data_buf[12] ),
    .S(_0838_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1014_));
 sky130_fd_sc_hd__inv_2 _4168_ (.A(_0866_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1015_));
 sky130_fd_sc_hd__and3_1 _4169_ (.A(\i_tinyqv.cpu.data_read_n[0] ),
    .B(\i_tinyqv.cpu.data_write_n[0] ),
    .C(_1015_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1016_));
 sky130_fd_sc_hd__nand2_4 _4170_ (.A(_0979_),
    .B(_1016_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1017_));
 sky130_fd_sc_hd__mux2_1 _4171_ (.A0(_0976_),
    .A1(_1014_),
    .S(_1017_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1018_));
 sky130_fd_sc_hd__mux2_1 _4172_ (.A0(_1013_),
    .A1(_1018_),
    .S(_0907_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1019_));
 sky130_fd_sc_hd__o22a_1 _4173_ (.A1(_0982_),
    .A2(_1010_),
    .B1(_1019_),
    .B2(_0957_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1020_));
 sky130_fd_sc_hd__a21o_1 _4174_ (.A1(_0956_),
    .A2(_0981_),
    .B1(_1020_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1021_));
 sky130_fd_sc_hd__inv_2 _4175_ (.A(_0955_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1022_));
 sky130_fd_sc_hd__a21o_1 _4176_ (.A1(\i_tinyqv.cpu.i_core.load_top_bit ),
    .A2(_1022_),
    .B1(_0878_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1023_));
 sky130_fd_sc_hd__a21o_1 _4177_ (.A1(_0955_),
    .A2(_1021_),
    .B1(_1023_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1024_));
 sky130_fd_sc_hd__nand2_1 _4178_ (.A(_0852_),
    .B(_0849_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1025_));
 sky130_fd_sc_hd__clkbuf_4 _4179_ (.A(_0946_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1026_));
 sky130_fd_sc_hd__clkbuf_4 _4180_ (.A(\i_tinyqv.cpu.alu_op[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1027_));
 sky130_fd_sc_hd__clkbuf_4 _4181_ (.A(_1027_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1028_));
 sky130_fd_sc_hd__clkbuf_4 _4182_ (.A(_1028_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1029_));
 sky130_fd_sc_hd__buf_2 _4183_ (.A(_1029_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1030_));
 sky130_fd_sc_hd__or2_4 _4184_ (.A(\i_tinyqv.cpu.i_core.cycle[1] ),
    .B(_0842_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1031_));
 sky130_fd_sc_hd__or4_1 _4185_ (.A(_1030_),
    .B(_0844_),
    .C(\i_tinyqv.cpu.alu_op[3] ),
    .D(_1031_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1032_));
 sky130_fd_sc_hd__nor2_1 _4186_ (.A(_1026_),
    .B(_1032_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1033_));
 sky130_fd_sc_hd__nor2_1 _4187_ (.A(_1033_),
    .B(_0877_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1034_));
 sky130_fd_sc_hd__a21o_1 _4188_ (.A1(\i_tinyqv.cpu.i_core.cmp ),
    .A2(_1025_),
    .B1(_1034_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1035_));
 sky130_fd_sc_hd__buf_4 _4189_ (.A(_1027_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1036_));
 sky130_fd_sc_hd__xnor2_1 _4190_ (.A(_0688_),
    .B(_1036_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1037_));
 sky130_fd_sc_hd__or2_1 _4191_ (.A(\i_tinyqv.cpu.i_core.i_shift.b[4] ),
    .B(_1037_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1038_));
 sky130_fd_sc_hd__xnor2_1 _4192_ (.A(_0907_),
    .B(_1027_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1039_));
 sky130_fd_sc_hd__xnor2_1 _4193_ (.A(\i_tinyqv.cpu.i_core.i_shift.b[3] ),
    .B(_1039_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1040_));
 sky130_fd_sc_hd__xnor2_1 _4194_ (.A(_0838_),
    .B(_1027_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1041_));
 sky130_fd_sc_hd__nand2_1 _4195_ (.A(\i_tinyqv.cpu.i_core.i_shift.b[2] ),
    .B(_1041_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1042_));
 sky130_fd_sc_hd__nor2_1 _4196_ (.A(_1040_),
    .B(_1042_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1043_));
 sky130_fd_sc_hd__a21o_1 _4197_ (.A1(\i_tinyqv.cpu.i_core.i_shift.b[3] ),
    .A2(_1039_),
    .B1(_1043_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1044_));
 sky130_fd_sc_hd__nand2_1 _4198_ (.A(\i_tinyqv.cpu.i_core.i_shift.b[4] ),
    .B(_1037_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1045_));
 sky130_fd_sc_hd__a21boi_2 _4199_ (.A1(_1038_),
    .A2(_1044_),
    .B1_N(_1045_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1046_));
 sky130_fd_sc_hd__and2_1 _4200_ (.A(_1040_),
    .B(_1042_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1047_));
 sky130_fd_sc_hd__or2_2 _4201_ (.A(_1043_),
    .B(_1047_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1048_));
 sky130_fd_sc_hd__mux4_1 _4202_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[31] ),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[30] ),
    .A2(\i_tinyqv.cpu.i_core.i_shift.a[0] ),
    .A3(\i_tinyqv.cpu.i_core.i_shift.a[1] ),
    .S0(\i_tinyqv.cpu.i_core.i_shift.adjusted_shift_amt[0] ),
    .S1(_1029_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1049_));
 sky130_fd_sc_hd__clkbuf_4 _4203_ (.A(\i_tinyqv.cpu.i_core.i_shift.adjusted_shift_amt[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1050_));
 sky130_fd_sc_hd__mux4_1 _4204_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[29] ),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[2] ),
    .A2(\i_tinyqv.cpu.i_core.i_shift.a[28] ),
    .A3(\i_tinyqv.cpu.i_core.i_shift.a[3] ),
    .S0(_1036_),
    .S1(_1050_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1051_));
 sky130_fd_sc_hd__mux2_1 _4205_ (.A0(_1049_),
    .A1(_1051_),
    .S(\i_tinyqv.cpu.i_core.i_shift.adjusted_shift_amt[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1052_));
 sky130_fd_sc_hd__mux4_1 _4206_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[27] ),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[26] ),
    .A2(\i_tinyqv.cpu.i_core.i_shift.a[4] ),
    .A3(\i_tinyqv.cpu.i_core.i_shift.a[5] ),
    .S0(\i_tinyqv.cpu.i_core.i_shift.adjusted_shift_amt[0] ),
    .S1(_1029_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1053_));
 sky130_fd_sc_hd__clkbuf_4 _4207_ (.A(\i_tinyqv.cpu.i_core.i_shift.a[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1054_));
 sky130_fd_sc_hd__mux4_1 _4208_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[25] ),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[24] ),
    .A2(\i_tinyqv.cpu.i_core.i_shift.a[6] ),
    .A3(_1054_),
    .S0(\i_tinyqv.cpu.i_core.i_shift.adjusted_shift_amt[0] ),
    .S1(_1029_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1055_));
 sky130_fd_sc_hd__mux2_1 _4209_ (.A0(_1053_),
    .A1(_1055_),
    .S(\i_tinyqv.cpu.i_core.i_shift.adjusted_shift_amt[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1056_));
 sky130_fd_sc_hd__or2_1 _4210_ (.A(\i_tinyqv.cpu.i_core.i_shift.b[2] ),
    .B(_1041_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1057_));
 sky130_fd_sc_hd__and2_2 _4211_ (.A(_1042_),
    .B(_1057_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1058_));
 sky130_fd_sc_hd__mux2_1 _4212_ (.A0(_1052_),
    .A1(_1056_),
    .S(_1058_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1059_));
 sky130_fd_sc_hd__buf_2 _4213_ (.A(\i_tinyqv.cpu.i_core.i_shift.a[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1060_));
 sky130_fd_sc_hd__mux2_1 _4214_ (.A0(_1060_),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[16] ),
    .S(_1028_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1061_));
 sky130_fd_sc_hd__mux2_1 _4215_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[14] ),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[17] ),
    .S(_1027_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1062_));
 sky130_fd_sc_hd__mux2_1 _4216_ (.A0(_1061_),
    .A1(_1062_),
    .S(_1050_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1063_));
 sky130_fd_sc_hd__mux2_1 _4217_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[13] ),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[18] ),
    .S(_1027_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1064_));
 sky130_fd_sc_hd__mux2_1 _4218_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[12] ),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[19] ),
    .S(_1027_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1065_));
 sky130_fd_sc_hd__mux2_1 _4219_ (.A0(_1064_),
    .A1(_1065_),
    .S(_1050_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1066_));
 sky130_fd_sc_hd__mux2_1 _4220_ (.A0(_1063_),
    .A1(_1066_),
    .S(\i_tinyqv.cpu.i_core.i_shift.adjusted_shift_amt[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1067_));
 sky130_fd_sc_hd__mux2_1 _4221_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[11] ),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[20] ),
    .S(_1028_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1068_));
 sky130_fd_sc_hd__mux2_1 _4222_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[10] ),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[21] ),
    .S(_1027_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1069_));
 sky130_fd_sc_hd__mux2_1 _4223_ (.A0(_1068_),
    .A1(_1069_),
    .S(_1050_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1070_));
 sky130_fd_sc_hd__mux2_1 _4224_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[9] ),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[22] ),
    .S(_1027_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1071_));
 sky130_fd_sc_hd__mux2_1 _4225_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[8] ),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[23] ),
    .S(_1027_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1072_));
 sky130_fd_sc_hd__mux2_1 _4226_ (.A0(_1071_),
    .A1(_1072_),
    .S(\i_tinyqv.cpu.i_core.i_shift.adjusted_shift_amt[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1073_));
 sky130_fd_sc_hd__mux2_1 _4227_ (.A0(_1070_),
    .A1(_1073_),
    .S(\i_tinyqv.cpu.i_core.i_shift.adjusted_shift_amt[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1074_));
 sky130_fd_sc_hd__mux2_1 _4228_ (.A0(_1067_),
    .A1(_1074_),
    .S(_1058_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1075_));
 sky130_fd_sc_hd__a21o_1 _4229_ (.A1(_1038_),
    .A2(_1045_),
    .B1(_1044_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1076_));
 sky130_fd_sc_hd__clkbuf_4 _4230_ (.A(_1076_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1077_));
 sky130_fd_sc_hd__mux2_1 _4231_ (.A0(_1059_),
    .A1(_1075_),
    .S(_1077_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1078_));
 sky130_fd_sc_hd__nand2_1 _4232_ (.A(_1048_),
    .B(_1078_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1079_));
 sky130_fd_sc_hd__buf_2 _4233_ (.A(_1058_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1080_));
 sky130_fd_sc_hd__mux2_1 _4234_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[3] ),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[28] ),
    .S(_1029_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1081_));
 sky130_fd_sc_hd__mux2_1 _4235_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[2] ),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[29] ),
    .S(_1036_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1082_));
 sky130_fd_sc_hd__clkbuf_4 _4236_ (.A(_1050_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1083_));
 sky130_fd_sc_hd__mux2_1 _4237_ (.A0(_1081_),
    .A1(_1082_),
    .S(_1083_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1084_));
 sky130_fd_sc_hd__mux2_1 _4238_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[1] ),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[30] ),
    .S(_1036_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1085_));
 sky130_fd_sc_hd__mux2_1 _4239_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[0] ),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[31] ),
    .S(_1036_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1086_));
 sky130_fd_sc_hd__mux2_1 _4240_ (.A0(_1085_),
    .A1(_1086_),
    .S(_1083_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1087_));
 sky130_fd_sc_hd__clkbuf_4 _4241_ (.A(\i_tinyqv.cpu.i_core.i_shift.adjusted_shift_amt[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1088_));
 sky130_fd_sc_hd__mux2_1 _4242_ (.A0(_1084_),
    .A1(_1087_),
    .S(_1088_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1089_));
 sky130_fd_sc_hd__nand2_1 _4243_ (.A(_1080_),
    .B(_1089_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1090_));
 sky130_fd_sc_hd__nand2_2 _4244_ (.A(_1042_),
    .B(_1057_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1091_));
 sky130_fd_sc_hd__buf_2 _4245_ (.A(_1091_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1092_));
 sky130_fd_sc_hd__mux2_1 _4246_ (.A0(_1054_),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[24] ),
    .S(_1036_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1093_));
 sky130_fd_sc_hd__mux2_1 _4247_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[6] ),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[25] ),
    .S(_1036_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1094_));
 sky130_fd_sc_hd__mux2_1 _4248_ (.A0(_1093_),
    .A1(_1094_),
    .S(_1083_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1095_));
 sky130_fd_sc_hd__mux2_1 _4249_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[5] ),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[26] ),
    .S(_1036_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1096_));
 sky130_fd_sc_hd__mux2_1 _4250_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[4] ),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[27] ),
    .S(_1029_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1097_));
 sky130_fd_sc_hd__mux2_1 _4251_ (.A0(_1096_),
    .A1(_1097_),
    .S(_1083_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1098_));
 sky130_fd_sc_hd__mux2_1 _4252_ (.A0(_1095_),
    .A1(_1098_),
    .S(_1088_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1099_));
 sky130_fd_sc_hd__nand2_1 _4253_ (.A(_1092_),
    .B(_1099_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1100_));
 sky130_fd_sc_hd__mux2_1 _4254_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[23] ),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[8] ),
    .S(_1028_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1101_));
 sky130_fd_sc_hd__mux2_1 _4255_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[22] ),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[9] ),
    .S(_1028_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1102_));
 sky130_fd_sc_hd__clkbuf_4 _4256_ (.A(\i_tinyqv.cpu.i_core.i_shift.adjusted_shift_amt[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1103_));
 sky130_fd_sc_hd__mux2_1 _4257_ (.A0(_1101_),
    .A1(_1102_),
    .S(_1103_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1104_));
 sky130_fd_sc_hd__mux2_1 _4258_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[21] ),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[10] ),
    .S(_1028_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1105_));
 sky130_fd_sc_hd__mux2_1 _4259_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[20] ),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[11] ),
    .S(_1028_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1106_));
 sky130_fd_sc_hd__mux2_1 _4260_ (.A0(_1105_),
    .A1(_1106_),
    .S(_1103_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1107_));
 sky130_fd_sc_hd__clkbuf_4 _4261_ (.A(\i_tinyqv.cpu.i_core.i_shift.adjusted_shift_amt[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1108_));
 sky130_fd_sc_hd__mux2_1 _4262_ (.A0(_1104_),
    .A1(_1107_),
    .S(_1108_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1109_));
 sky130_fd_sc_hd__mux2_1 _4263_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[19] ),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[12] ),
    .S(_1028_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1110_));
 sky130_fd_sc_hd__mux2_1 _4264_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[18] ),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[13] ),
    .S(_1028_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1111_));
 sky130_fd_sc_hd__mux2_1 _4265_ (.A0(_1110_),
    .A1(_1111_),
    .S(_1103_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1112_));
 sky130_fd_sc_hd__mux2_1 _4266_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[17] ),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[14] ),
    .S(_1028_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1113_));
 sky130_fd_sc_hd__mux2_1 _4267_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[16] ),
    .A1(_1060_),
    .S(_1036_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1114_));
 sky130_fd_sc_hd__mux2_1 _4268_ (.A0(_1113_),
    .A1(_1114_),
    .S(_1050_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1115_));
 sky130_fd_sc_hd__mux2_1 _4269_ (.A0(_1112_),
    .A1(_1115_),
    .S(_1108_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1116_));
 sky130_fd_sc_hd__a21o_1 _4270_ (.A1(_1080_),
    .A2(_1116_),
    .B1(_1076_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1117_));
 sky130_fd_sc_hd__a21oi_1 _4271_ (.A1(_1092_),
    .A2(_1109_),
    .B1(_1117_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1118_));
 sky130_fd_sc_hd__a311o_1 _4272_ (.A1(_1077_),
    .A2(_1090_),
    .A3(_1100_),
    .B1(_1118_),
    .C1(_1048_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1119_));
 sky130_fd_sc_hd__nand2_1 _4273_ (.A(\i_tinyqv.cpu.alu_op[3] ),
    .B(\i_tinyqv.cpu.i_core.i_shift.a[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1120_));
 sky130_fd_sc_hd__and2b_1 _4274_ (.A_N(_1046_),
    .B(_1120_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1121_));
 sky130_fd_sc_hd__a31o_1 _4275_ (.A1(_1046_),
    .A2(_1079_),
    .A3(_1119_),
    .B1(_1121_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1122_));
 sky130_fd_sc_hd__nand2_1 _4276_ (.A(_1030_),
    .B(_1122_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1123_));
 sky130_fd_sc_hd__nand2_4 _4277_ (.A(_0844_),
    .B(net69),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1124_));
 sky130_fd_sc_hd__nor2_2 _4278_ (.A(_1124_),
    .B(_1031_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1125_));
 sky130_fd_sc_hd__mux2_1 _4279_ (.A0(_1065_),
    .A1(_1068_),
    .S(_1103_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1126_));
 sky130_fd_sc_hd__mux2_1 _4280_ (.A0(_1069_),
    .A1(_1071_),
    .S(_1103_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1127_));
 sky130_fd_sc_hd__mux2_1 _4281_ (.A0(_1126_),
    .A1(_1127_),
    .S(_1088_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1128_));
 sky130_fd_sc_hd__nand2_1 _4282_ (.A(_1092_),
    .B(_1128_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1129_));
 sky130_fd_sc_hd__mux2_1 _4283_ (.A0(_1072_),
    .A1(_1093_),
    .S(_1103_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1130_));
 sky130_fd_sc_hd__mux2_1 _4284_ (.A0(_1094_),
    .A1(_1096_),
    .S(_1083_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1131_));
 sky130_fd_sc_hd__mux2_1 _4285_ (.A0(_1130_),
    .A1(_1131_),
    .S(_1088_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1132_));
 sky130_fd_sc_hd__nand2_1 _4286_ (.A(_1080_),
    .B(_1132_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1133_));
 sky130_fd_sc_hd__mux4_1 _4287_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[28] ),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[3] ),
    .A2(\i_tinyqv.cpu.i_core.i_shift.a[27] ),
    .A3(\i_tinyqv.cpu.i_core.i_shift.a[4] ),
    .S0(_1029_),
    .S1(_1103_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1134_));
 sky130_fd_sc_hd__mux4_1 _4288_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[26] ),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[25] ),
    .A2(\i_tinyqv.cpu.i_core.i_shift.a[5] ),
    .A3(\i_tinyqv.cpu.i_core.i_shift.a[6] ),
    .S0(\i_tinyqv.cpu.i_core.i_shift.adjusted_shift_amt[0] ),
    .S1(_1029_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1135_));
 sky130_fd_sc_hd__mux2_1 _4289_ (.A0(_1134_),
    .A1(_1135_),
    .S(_1108_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1136_));
 sky130_fd_sc_hd__mux2_1 _4290_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[24] ),
    .A1(_1054_),
    .S(_1036_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1137_));
 sky130_fd_sc_hd__mux2_1 _4291_ (.A0(_1137_),
    .A1(_1101_),
    .S(_1050_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1138_));
 sky130_fd_sc_hd__mux2_1 _4292_ (.A0(_1102_),
    .A1(_1105_),
    .S(_1050_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1139_));
 sky130_fd_sc_hd__mux2_1 _4293_ (.A0(_1138_),
    .A1(_1139_),
    .S(\i_tinyqv.cpu.i_core.i_shift.adjusted_shift_amt[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1140_));
 sky130_fd_sc_hd__a21o_1 _4294_ (.A1(_1080_),
    .A2(_1140_),
    .B1(_1076_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1141_));
 sky130_fd_sc_hd__a21oi_1 _4295_ (.A1(_1091_),
    .A2(_1136_),
    .B1(_1141_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1142_));
 sky130_fd_sc_hd__nor2_1 _4296_ (.A(_1043_),
    .B(_1047_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1143_));
 sky130_fd_sc_hd__a311o_1 _4297_ (.A1(_1077_),
    .A2(_1129_),
    .A3(_1133_),
    .B1(_1142_),
    .C1(_1143_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1144_));
 sky130_fd_sc_hd__mux2_1 _4298_ (.A0(_1097_),
    .A1(_1081_),
    .S(_1083_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1145_));
 sky130_fd_sc_hd__mux2_1 _4299_ (.A0(_1082_),
    .A1(_1085_),
    .S(_1083_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1146_));
 sky130_fd_sc_hd__mux2_1 _4300_ (.A0(_1145_),
    .A1(_1146_),
    .S(_1088_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1147_));
 sky130_fd_sc_hd__nand2_1 _4301_ (.A(_1092_),
    .B(_1147_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1148_));
 sky130_fd_sc_hd__clkbuf_4 _4302_ (.A(_1108_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1149_));
 sky130_fd_sc_hd__nor2_1 _4303_ (.A(_1083_),
    .B(_1086_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1150_));
 sky130_fd_sc_hd__a21oi_1 _4304_ (.A1(_1083_),
    .A2(_1120_),
    .B1(_1150_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1151_));
 sky130_fd_sc_hd__nor2_1 _4305_ (.A(_1088_),
    .B(_1151_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1152_));
 sky130_fd_sc_hd__a211o_1 _4306_ (.A1(_1149_),
    .A2(_1120_),
    .B1(_1091_),
    .C1(_1152_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1153_));
 sky130_fd_sc_hd__mux2_1 _4307_ (.A0(_1114_),
    .A1(_1061_),
    .S(_1103_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1154_));
 sky130_fd_sc_hd__mux2_1 _4308_ (.A0(_1062_),
    .A1(_1064_),
    .S(_1103_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1155_));
 sky130_fd_sc_hd__mux2_1 _4309_ (.A0(_1154_),
    .A1(_1155_),
    .S(_1108_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1156_));
 sky130_fd_sc_hd__mux2_1 _4310_ (.A0(_1106_),
    .A1(_1110_),
    .S(_1050_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1157_));
 sky130_fd_sc_hd__mux2_1 _4311_ (.A0(_1111_),
    .A1(_1113_),
    .S(_1050_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1158_));
 sky130_fd_sc_hd__mux2_1 _4312_ (.A0(_1157_),
    .A1(_1158_),
    .S(\i_tinyqv.cpu.i_core.i_shift.adjusted_shift_amt[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1159_));
 sky130_fd_sc_hd__a21o_1 _4313_ (.A1(_1091_),
    .A2(_1159_),
    .B1(_1076_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1160_));
 sky130_fd_sc_hd__a21oi_1 _4314_ (.A1(_1080_),
    .A2(_1156_),
    .B1(_1160_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1161_));
 sky130_fd_sc_hd__a311o_1 _4315_ (.A1(_1077_),
    .A2(_1148_),
    .A3(_1153_),
    .B1(_1161_),
    .C1(_1048_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1162_));
 sky130_fd_sc_hd__a31o_1 _4316_ (.A1(_1046_),
    .A2(_1144_),
    .A3(_1162_),
    .B1(_1121_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1163_));
 sky130_fd_sc_hd__nand2_1 _4317_ (.A(_0843_),
    .B(_1163_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1164_));
 sky130_fd_sc_hd__and3_1 _4318_ (.A(_1123_),
    .B(_1125_),
    .C(_1164_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1165_));
 sky130_fd_sc_hd__a21oi_4 _4319_ (.A1(net45),
    .A2(net64),
    .B1(_0842_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1166_));
 sky130_fd_sc_hd__clkbuf_4 _4320_ (.A(_1166_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1167_));
 sky130_fd_sc_hd__a21o_1 _4321_ (.A1(\i_tinyqv.cpu.i_core.i_shift.a[0] ),
    .A2(_1167_),
    .B1(\i_tinyqv.cpu.i_core.multiplier.accum[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1168_));
 sky130_fd_sc_hd__nand3_1 _4322_ (.A(\i_tinyqv.cpu.i_core.i_shift.a[0] ),
    .B(\i_tinyqv.cpu.i_core.multiplier.accum[0] ),
    .C(_1167_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1169_));
 sky130_fd_sc_hd__inv_2 _4323_ (.A(_0847_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1170_));
 sky130_fd_sc_hd__and2b_1 _4324_ (.A_N(_0746_),
    .B(_0743_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1171_));
 sky130_fd_sc_hd__nand2_1 _4325_ (.A(_1171_),
    .B(_0745_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1172_));
 sky130_fd_sc_hd__nand2_2 _4326_ (.A(_0843_),
    .B(_0919_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1173_));
 sky130_fd_sc_hd__o21ba_1 _4327_ (.A1(_1171_),
    .A2(_0745_),
    .B1_N(_1173_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1174_));
 sky130_fd_sc_hd__and3b_1 _4328_ (.A_N(net69),
    .B(_0656_),
    .C(_1030_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1175_));
 sky130_fd_sc_hd__o31a_1 _4329_ (.A1(_0742_),
    .A2(_0708_),
    .A3(net78),
    .B1(_1175_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1176_));
 sky130_fd_sc_hd__nand2_1 _4330_ (.A(_1030_),
    .B(_0919_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1177_));
 sky130_fd_sc_hd__and3_1 _4331_ (.A(_1029_),
    .B(_0656_),
    .C(\i_tinyqv.cpu.alu_op[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1178_));
 sky130_fd_sc_hd__o21a_1 _4332_ (.A1(_0708_),
    .A2(net79),
    .B1(_1178_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1179_));
 sky130_fd_sc_hd__a2bb2o_1 _4333_ (.A1_N(_0830_),
    .A2_N(_1177_),
    .B1(_1179_),
    .B2(_0742_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1180_));
 sky130_fd_sc_hd__a211o_1 _4334_ (.A1(_1172_),
    .A2(_1174_),
    .B1(_1176_),
    .C1(_1180_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1181_));
 sky130_fd_sc_hd__a32o_1 _4335_ (.A1(_0846_),
    .A2(_1168_),
    .A3(_1169_),
    .B1(_1170_),
    .B2(_1181_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1182_));
 sky130_fd_sc_hd__or3_1 _4336_ (.A(_1165_),
    .B(_1033_),
    .C(_1182_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1183_));
 sky130_fd_sc_hd__a32o_1 _4337_ (.A1(_0877_),
    .A2(_0954_),
    .A3(_1024_),
    .B1(_1035_),
    .B2(_1183_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1184_));
 sky130_fd_sc_hd__clkbuf_4 _4338_ (.A(_1184_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.debug_rd[0] ));
 sky130_fd_sc_hd__or2_1 _4339_ (.A(_0855_),
    .B(_0919_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1185_));
 sky130_fd_sc_hd__and4_1 _4340_ (.A(_0857_),
    .B(_0858_),
    .C(_0878_),
    .D(_1185_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1186_));
 sky130_fd_sc_hd__and3_1 _4341_ (.A(_0842_),
    .B(_0846_),
    .C(_1025_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1187_));
 sky130_fd_sc_hd__a21oi_4 _4342_ (.A1(_0877_),
    .A2(_1186_),
    .B1(_1187_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1188_));
 sky130_fd_sc_hd__and3_1 _4343_ (.A(\i_tinyqv.cpu.i_core.i_registers.rd[2] ),
    .B(\i_tinyqv.cpu.i_core.i_registers.rd[3] ),
    .C(_1188_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1189_));
 sky130_fd_sc_hd__and3_2 _4344_ (.A(\i_tinyqv.cpu.i_core.i_registers.rd[1] ),
    .B(\i_tinyqv.cpu.i_core.i_registers.rd[0] ),
    .C(_1189_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1190_));
 sky130_fd_sc_hd__mux2_1 _4345_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[15][0] ),
    .A1(\i_tinyqv.cpu.debug_rd[0] ),
    .S(_1190_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1191_));
 sky130_fd_sc_hd__clkbuf_1 _4346_ (.A(_1191_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0050_));
 sky130_fd_sc_hd__mux2_1 _4347_ (.A0(\i_uart_rx.uart_rts ),
    .A1(\gpio_out[1] ),
    .S(\gpio_out_sel[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1192_));
 sky130_fd_sc_hd__buf_4 _4348_ (.A(_1192_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[1]));
 sky130_fd_sc_hd__mux2_1 _4349_ (.A0(\i_spi.spi_clk_out ),
    .A1(\debug_rd_r[3] ),
    .S(debug_register_data),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1193_));
 sky130_fd_sc_hd__mux2_1 _4350_ (.A0(_1193_),
    .A1(\gpio_out[5] ),
    .S(\gpio_out_sel[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1194_));
 sky130_fd_sc_hd__clkbuf_4 _4351_ (.A(_1194_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[5]));
 sky130_fd_sc_hd__a22o_1 _4352_ (.A1(\i_tinyqv.cpu.i_core.mip[17] ),
    .A2(_0943_),
    .B1(_0944_),
    .B2(\i_tinyqv.cpu.i_core.mie[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1195_));
 sky130_fd_sc_hd__mux2_1 _4353_ (.A0(\i_tinyqv.cpu.i_core.time_hi[0] ),
    .A1(\i_tinyqv.cpu.i_core.cycle_count_wide[4] ),
    .S(_0841_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1196_));
 sky130_fd_sc_hd__a22o_1 _4354_ (.A1(\i_tinyqv.cpu.i_core.cycle_count[1] ),
    .A2(_0931_),
    .B1(_1196_),
    .B2(_0927_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1197_));
 sky130_fd_sc_hd__a221o_1 _4355_ (.A1(\i_tinyqv.cpu.i_core.mcause[1] ),
    .A2(_0947_),
    .B1(_0929_),
    .B2(\i_tinyqv.cpu.i_core.i_instrret.data[1] ),
    .C1(_1197_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1198_));
 sky130_fd_sc_hd__a211o_1 _4356_ (.A1(\i_tinyqv.cpu.i_core.mepc[1] ),
    .A2(net19),
    .B1(_1195_),
    .C1(_1198_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1199_));
 sky130_fd_sc_hd__a21oi_1 _4357_ (.A1(_0726_),
    .A2(_0894_),
    .B1(\i_tinyqv.cpu.instr_data_start[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1200_));
 sky130_fd_sc_hd__or2_1 _4358_ (.A(_0895_),
    .B(_1200_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1201_));
 sky130_fd_sc_hd__xor2_1 _4359_ (.A(_0882_),
    .B(_0892_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1202_));
 sky130_fd_sc_hd__inv_2 _4360_ (.A(_1202_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1203_));
 sky130_fd_sc_hd__nor2_1 _4361_ (.A(\i_tinyqv.cpu.instr_data_start[5] ),
    .B(_0889_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1204_));
 sky130_fd_sc_hd__or2_1 _4362_ (.A(_0890_),
    .B(_1204_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1205_));
 sky130_fd_sc_hd__nand2_2 _4363_ (.A(\i_tinyqv.cpu.instr_len[1] ),
    .B(\i_tinyqv.cpu.pc[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1206_));
 sky130_fd_sc_hd__or2_1 _4364_ (.A(\i_tinyqv.cpu.instr_len[1] ),
    .B(\i_tinyqv.cpu.pc[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1207_));
 sky130_fd_sc_hd__nand2_2 _4365_ (.A(_1206_),
    .B(_1207_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1208_));
 sky130_fd_sc_hd__a221o_1 _4366_ (.A1(_0748_),
    .A2(_1205_),
    .B1(_1208_),
    .B2(_0689_),
    .C1(_0688_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1209_));
 sky130_fd_sc_hd__a221o_1 _4367_ (.A1(_0617_),
    .A2(_1201_),
    .B1(_1203_),
    .B2(_0691_),
    .C1(_1209_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1210_));
 sky130_fd_sc_hd__xor2_1 _4368_ (.A(\i_tinyqv.cpu.instr_data_start[21] ),
    .B(_0900_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1211_));
 sky130_fd_sc_hd__nor2_1 _4369_ (.A(\i_tinyqv.cpu.instr_data_start[17] ),
    .B(_0897_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1212_));
 sky130_fd_sc_hd__or2_1 _4370_ (.A(_0898_),
    .B(_1212_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1213_));
 sky130_fd_sc_hd__o2bb2a_1 _4371_ (.A1_N(_0610_),
    .A2_N(_1211_),
    .B1(_1213_),
    .B2(_0916_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1214_));
 sky130_fd_sc_hd__a21oi_1 _4372_ (.A1(_1210_),
    .A2(_1214_),
    .B1(_0858_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1215_));
 sky130_fd_sc_hd__a211o_1 _4373_ (.A1(_0921_),
    .A2(_1199_),
    .B1(_1215_),
    .C1(_0880_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1216_));
 sky130_fd_sc_hd__o21ai_1 _4374_ (.A1(_0777_),
    .A2(_0857_),
    .B1(_1216_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1217_));
 sky130_fd_sc_hd__nand2_1 _4375_ (.A(_0878_),
    .B(_1217_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1218_));
 sky130_fd_sc_hd__a221o_1 _4376_ (.A1(\i_tinyqv.mem.data_from_read[17] ),
    .A2(_0689_),
    .B1(_0748_),
    .B2(\i_tinyqv.mem.data_from_read[21] ),
    .C1(_0957_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1219_));
 sky130_fd_sc_hd__mux2_1 _4377_ (.A0(\i_tinyqv.mem.qspi_data_buf[25] ),
    .A1(\i_tinyqv.mem.qspi_data_buf[29] ),
    .S(_0974_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1220_));
 sky130_fd_sc_hd__mux2_1 _4378_ (.A0(\i_tinyqv.cpu.instr_data_in[9] ),
    .A1(\i_tinyqv.cpu.instr_data_in[13] ),
    .S(_0838_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1221_));
 sky130_fd_sc_hd__mux2_1 _4379_ (.A0(_1220_),
    .A1(_1221_),
    .S(_0979_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1222_));
 sky130_fd_sc_hd__a22o_1 _4380_ (.A1(_0971_),
    .A2(_1219_),
    .B1(_1222_),
    .B2(_0973_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1223_));
 sky130_fd_sc_hd__a221o_1 _4381_ (.A1(\i_uart_rx.recieved_data[1] ),
    .A2(_0997_),
    .B1(uo_out[1]),
    .B2(_1001_),
    .C1(_0974_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1224_));
 sky130_fd_sc_hd__inv_2 _4382_ (.A(_0985_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1225_));
 sky130_fd_sc_hd__inv_2 _4383_ (.A(\i_uart_rx.fsm_state[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1226_));
 sky130_fd_sc_hd__nand3b_4 _4384_ (.A_N(\i_uart_rx.fsm_state[2] ),
    .B(\i_uart_rx.fsm_state[1] ),
    .C(\i_uart_rx.fsm_state[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1227_));
 sky130_fd_sc_hd__nor2_4 _4385_ (.A(_1226_),
    .B(_1227_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1228_));
 sky130_fd_sc_hd__a32o_1 _4386_ (.A1(_1225_),
    .A2(_0987_),
    .A3(_1228_),
    .B1(_1003_),
    .B2(\gpio_out_sel[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1229_));
 sky130_fd_sc_hd__a221o_1 _4387_ (.A1(\i_spi.data[1] ),
    .A2(_1000_),
    .B1(_0986_),
    .B2(net3),
    .C1(_1229_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1230_));
 sky130_fd_sc_hd__a22o_1 _4388_ (.A1(net7),
    .A2(_0986_),
    .B1(_1001_),
    .B2(uo_out[5]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1231_));
 sky130_fd_sc_hd__a221o_1 _4389_ (.A1(\i_spi.data[5] ),
    .A2(_1000_),
    .B1(_0997_),
    .B2(\i_uart_rx.recieved_data[5] ),
    .C1(_0908_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1232_));
 sky130_fd_sc_hd__a211o_1 _4390_ (.A1(\gpio_out_sel[5] ),
    .A2(net14),
    .B1(_1231_),
    .C1(_1232_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1233_));
 sky130_fd_sc_hd__o211a_1 _4391_ (.A1(_1224_),
    .A2(_1230_),
    .B1(_0945_),
    .C1(_1233_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1234_));
 sky130_fd_sc_hd__mux2_1 _4392_ (.A0(\i_tinyqv.cpu.instr_data_in[13] ),
    .A1(\i_tinyqv.mem.qspi_data_buf[13] ),
    .S(_1017_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1235_));
 sky130_fd_sc_hd__mux2_1 _4393_ (.A0(\i_tinyqv.cpu.instr_data_in[1] ),
    .A1(\i_tinyqv.cpu.instr_data_in[5] ),
    .S(_0838_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1236_));
 sky130_fd_sc_hd__mux2_1 _4394_ (.A0(_1221_),
    .A1(_1236_),
    .S(_1012_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1237_));
 sky130_fd_sc_hd__mux2_1 _4395_ (.A0(\i_tinyqv.cpu.instr_data_in[9] ),
    .A1(\i_tinyqv.mem.qspi_data_buf[9] ),
    .S(_1017_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1238_));
 sky130_fd_sc_hd__o22a_1 _4396_ (.A1(_0907_),
    .A2(_1237_),
    .B1(_1238_),
    .B2(_0909_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1239_));
 sky130_fd_sc_hd__o21a_1 _4397_ (.A1(_0724_),
    .A2(_1235_),
    .B1(_1239_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1240_));
 sky130_fd_sc_hd__o22a_1 _4398_ (.A1(_0982_),
    .A2(_1234_),
    .B1(_1240_),
    .B2(_0957_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1241_));
 sky130_fd_sc_hd__a21o_1 _4399_ (.A1(_0956_),
    .A2(_1223_),
    .B1(_1241_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1242_));
 sky130_fd_sc_hd__a21o_1 _4400_ (.A1(_0955_),
    .A2(_1242_),
    .B1(_1023_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1243_));
 sky130_fd_sc_hd__and3_1 _4401_ (.A(\i_tinyqv.cpu.i_core.i_shift.a[1] ),
    .B(\i_tinyqv.cpu.i_core.multiplier.accum[1] ),
    .C(_1166_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1244_));
 sky130_fd_sc_hd__a21oi_1 _4402_ (.A1(\i_tinyqv.cpu.i_core.i_shift.a[1] ),
    .A2(_1167_),
    .B1(\i_tinyqv.cpu.i_core.multiplier.accum[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1245_));
 sky130_fd_sc_hd__or2_1 _4403_ (.A(_1244_),
    .B(_1245_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1246_));
 sky130_fd_sc_hd__or2_1 _4404_ (.A(_1169_),
    .B(_1246_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1247_));
 sky130_fd_sc_hd__nand2_1 _4405_ (.A(_1169_),
    .B(_1246_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1248_));
 sky130_fd_sc_hd__nand2_1 _4406_ (.A(_1247_),
    .B(_1248_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1249_));
 sky130_fd_sc_hd__nor2_2 _4407_ (.A(_0842_),
    .B(net68),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1250_));
 sky130_fd_sc_hd__nand2_1 _4408_ (.A(\i_tinyqv.cpu.i_core.i_shift.a[0] ),
    .B(_1250_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1251_));
 sky130_fd_sc_hd__xor2_1 _4409_ (.A(_1249_),
    .B(_1251_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1252_));
 sky130_fd_sc_hd__or3b_1 _4410_ (.A(_0763_),
    .B(_0779_),
    .C_N(_1178_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1253_));
 sky130_fd_sc_hd__a21bo_1 _4411_ (.A1(_0763_),
    .A2(_0779_),
    .B1_N(_1175_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1254_));
 sky130_fd_sc_hd__a21oi_1 _4412_ (.A1(_0743_),
    .A2(_0745_),
    .B1(_0746_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1255_));
 sky130_fd_sc_hd__or2b_1 _4413_ (.A(_0782_),
    .B_N(_0781_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1256_));
 sky130_fd_sc_hd__or2_1 _4414_ (.A(_1255_),
    .B(_1256_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1257_));
 sky130_fd_sc_hd__a21oi_1 _4415_ (.A1(_1255_),
    .A2(_1256_),
    .B1(_1173_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1258_));
 sky130_fd_sc_hd__o2bb2a_1 _4416_ (.A1_N(_1257_),
    .A2_N(_1258_),
    .B1(_1177_),
    .B2(_0831_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1259_));
 sky130_fd_sc_hd__and3_1 _4417_ (.A(_1253_),
    .B(_1254_),
    .C(_1259_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1260_));
 sky130_fd_sc_hd__nor2_1 _4418_ (.A(_0846_),
    .B(_1260_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1261_));
 sky130_fd_sc_hd__mux2_1 _4419_ (.A0(_1098_),
    .A1(_1084_),
    .S(_1149_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1262_));
 sky130_fd_sc_hd__nand2_1 _4420_ (.A(_1092_),
    .B(_1262_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1263_));
 sky130_fd_sc_hd__nor2_1 _4421_ (.A(_1149_),
    .B(_1087_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1264_));
 sky130_fd_sc_hd__a211o_1 _4422_ (.A1(_1149_),
    .A2(_1120_),
    .B1(_1092_),
    .C1(_1264_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1265_));
 sky130_fd_sc_hd__mux2_1 _4423_ (.A0(_1107_),
    .A1(_1112_),
    .S(_1149_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1266_));
 sky130_fd_sc_hd__mux2_1 _4424_ (.A0(_1115_),
    .A1(_1063_),
    .S(_1088_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1267_));
 sky130_fd_sc_hd__a21o_1 _4425_ (.A1(_1080_),
    .A2(_1267_),
    .B1(_1077_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1268_));
 sky130_fd_sc_hd__a21oi_1 _4426_ (.A1(_1092_),
    .A2(_1266_),
    .B1(_1268_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1269_));
 sky130_fd_sc_hd__a311o_1 _4427_ (.A1(_1077_),
    .A2(_1263_),
    .A3(_1265_),
    .B1(_1269_),
    .C1(_1048_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1270_));
 sky130_fd_sc_hd__mux2_1 _4428_ (.A0(_1066_),
    .A1(_1070_),
    .S(_1149_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1271_));
 sky130_fd_sc_hd__nand2_1 _4429_ (.A(_1092_),
    .B(_1271_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1272_));
 sky130_fd_sc_hd__mux2_1 _4430_ (.A0(_1073_),
    .A1(_1095_),
    .S(_1149_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1273_));
 sky130_fd_sc_hd__nand2_1 _4431_ (.A(_1080_),
    .B(_1273_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1274_));
 sky130_fd_sc_hd__mux2_1 _4432_ (.A0(_1055_),
    .A1(_1104_),
    .S(_1149_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1275_));
 sky130_fd_sc_hd__mux2_1 _4433_ (.A0(_1051_),
    .A1(_1053_),
    .S(_1088_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1276_));
 sky130_fd_sc_hd__a21o_1 _4434_ (.A1(_1092_),
    .A2(_1276_),
    .B1(_1077_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1277_));
 sky130_fd_sc_hd__a21oi_1 _4435_ (.A1(_1080_),
    .A2(_1275_),
    .B1(_1277_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1278_));
 sky130_fd_sc_hd__a311o_1 _4436_ (.A1(_1077_),
    .A2(_1272_),
    .A3(_1274_),
    .B1(_1278_),
    .C1(_1143_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1279_));
 sky130_fd_sc_hd__a31oi_1 _4437_ (.A1(_1046_),
    .A2(_1270_),
    .A3(_1279_),
    .B1(_1121_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1280_));
 sky130_fd_sc_hd__mux4_1 _4438_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[30] ),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[1] ),
    .A2(\i_tinyqv.cpu.i_core.i_shift.a[29] ),
    .A3(\i_tinyqv.cpu.i_core.i_shift.a[2] ),
    .S0(_1029_),
    .S1(_1103_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1281_));
 sky130_fd_sc_hd__mux2_1 _4439_ (.A0(_1281_),
    .A1(_1134_),
    .S(_1108_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1282_));
 sky130_fd_sc_hd__mux2_1 _4440_ (.A0(_1135_),
    .A1(_1138_),
    .S(_1108_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1283_));
 sky130_fd_sc_hd__mux2_1 _4441_ (.A0(_1282_),
    .A1(_1283_),
    .S(_1058_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1284_));
 sky130_fd_sc_hd__mux2_1 _4442_ (.A0(_1155_),
    .A1(_1126_),
    .S(_1108_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1285_));
 sky130_fd_sc_hd__mux2_1 _4443_ (.A0(_1127_),
    .A1(_1130_),
    .S(_1108_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1286_));
 sky130_fd_sc_hd__mux2_1 _4444_ (.A0(_1285_),
    .A1(_1286_),
    .S(_1058_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1287_));
 sky130_fd_sc_hd__mux2_1 _4445_ (.A0(_1284_),
    .A1(_1287_),
    .S(_1077_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1288_));
 sky130_fd_sc_hd__nand2_1 _4446_ (.A(_1048_),
    .B(_1288_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1289_));
 sky130_fd_sc_hd__mux2_1 _4447_ (.A0(_1146_),
    .A1(_1151_),
    .S(_1149_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1290_));
 sky130_fd_sc_hd__nand2_1 _4448_ (.A(_1080_),
    .B(_1290_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1291_));
 sky130_fd_sc_hd__mux2_1 _4449_ (.A0(_1131_),
    .A1(_1145_),
    .S(_1088_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1292_));
 sky130_fd_sc_hd__nand2_1 _4450_ (.A(_1092_),
    .B(_1292_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1293_));
 sky130_fd_sc_hd__mux2_1 _4451_ (.A0(_1158_),
    .A1(_1154_),
    .S(_1088_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1294_));
 sky130_fd_sc_hd__mux2_1 _4452_ (.A0(_1139_),
    .A1(_1157_),
    .S(_1108_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1295_));
 sky130_fd_sc_hd__a21o_1 _4453_ (.A1(_1091_),
    .A2(_1295_),
    .B1(_1076_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1296_));
 sky130_fd_sc_hd__a21oi_1 _4454_ (.A1(_1080_),
    .A2(_1294_),
    .B1(_1296_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1297_));
 sky130_fd_sc_hd__a311o_1 _4455_ (.A1(_1077_),
    .A2(_1291_),
    .A3(_1293_),
    .B1(_1297_),
    .C1(_1048_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1298_));
 sky130_fd_sc_hd__a31o_1 _4456_ (.A1(_1046_),
    .A2(_1289_),
    .A3(_1298_),
    .B1(_1121_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1299_));
 sky130_fd_sc_hd__nand2_1 _4457_ (.A(_1030_),
    .B(_1299_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1300_));
 sky130_fd_sc_hd__o211a_1 _4458_ (.A1(_1030_),
    .A2(_1280_),
    .B1(_1300_),
    .C1(_1125_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1301_));
 sky130_fd_sc_hd__a211o_1 _4459_ (.A1(_0846_),
    .A2(_1252_),
    .B1(_1261_),
    .C1(_1301_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1302_));
 sky130_fd_sc_hd__a32o_2 _4460_ (.A1(_0877_),
    .A2(_1218_),
    .A3(_1243_),
    .B1(_1034_),
    .B2(_1302_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1303_));
 sky130_fd_sc_hd__buf_2 _4461_ (.A(_1303_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.debug_rd[1] ));
 sky130_fd_sc_hd__mux2_1 _4462_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[15][1] ),
    .A1(\i_tinyqv.cpu.debug_rd[1] ),
    .S(_1190_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1304_));
 sky130_fd_sc_hd__clkbuf_1 _4463_ (.A(_1304_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0051_));
 sky130_fd_sc_hd__mux2_1 _4464_ (.A0(\i_spi.spi_dc ),
    .A1(\debug_rd_r[0] ),
    .S(debug_register_data),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1305_));
 sky130_fd_sc_hd__mux2_1 _4465_ (.A0(_1305_),
    .A1(\gpio_out[2] ),
    .S(\gpio_out_sel[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1306_));
 sky130_fd_sc_hd__buf_4 _4466_ (.A(_1306_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[2]));
 sky130_fd_sc_hd__mux2_1 _4467_ (.A0(\i_debug_uart_tx.txd_reg ),
    .A1(\gpio_out[6] ),
    .S(\gpio_out_sel[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1307_));
 sky130_fd_sc_hd__clkbuf_4 _4468_ (.A(_1307_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[6]));
 sky130_fd_sc_hd__inv_2 _4469_ (.A(_1244_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1308_));
 sky130_fd_sc_hd__o21a_2 _4470_ (.A1(_0793_),
    .A2(_0797_),
    .B1(\i_tinyqv.cpu.i_core.cycle[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1309_));
 sky130_fd_sc_hd__and2_1 _4471_ (.A(\i_tinyqv.cpu.i_core.i_shift.a[0] ),
    .B(_1309_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1310_));
 sky130_fd_sc_hd__inv_2 _4472_ (.A(\i_tinyqv.cpu.i_core.i_shift.a[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1311_));
 sky130_fd_sc_hd__and2_2 _4473_ (.A(net44),
    .B(net65),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1312_));
 sky130_fd_sc_hd__or2_2 _4474_ (.A(_0842_),
    .B(_1312_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1313_));
 sky130_fd_sc_hd__nor2_1 _4475_ (.A(_1311_),
    .B(_1313_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1314_));
 sky130_fd_sc_hd__or3b_2 _4476_ (.A(_1311_),
    .B(_1313_),
    .C_N(_1310_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1315_));
 sky130_fd_sc_hd__o21a_1 _4477_ (.A1(_1310_),
    .A2(_1314_),
    .B1(_1315_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1316_));
 sky130_fd_sc_hd__xnor2_1 _4478_ (.A(\i_tinyqv.cpu.i_core.multiplier.accum[2] ),
    .B(_1316_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1317_));
 sky130_fd_sc_hd__xnor2_1 _4479_ (.A(_1308_),
    .B(_1317_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1318_));
 sky130_fd_sc_hd__nand2_1 _4480_ (.A(\i_tinyqv.cpu.i_core.i_shift.a[1] ),
    .B(_1250_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1319_));
 sky130_fd_sc_hd__xor2_1 _4481_ (.A(_1318_),
    .B(_1319_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1320_));
 sky130_fd_sc_hd__o21ai_1 _4482_ (.A1(_1249_),
    .A2(_1251_),
    .B1(_1247_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1321_));
 sky130_fd_sc_hd__nand2_1 _4483_ (.A(_1320_),
    .B(_1321_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1322_));
 sky130_fd_sc_hd__or2_1 _4484_ (.A(_1320_),
    .B(_1321_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1323_));
 sky130_fd_sc_hd__or2_1 _4485_ (.A(_0783_),
    .B(_0819_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1324_));
 sky130_fd_sc_hd__a21oi_1 _4486_ (.A1(_0783_),
    .A2(_0819_),
    .B1(_1173_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1325_));
 sky130_fd_sc_hd__nand2_1 _4487_ (.A(_1324_),
    .B(_1325_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1326_));
 sky130_fd_sc_hd__o21ba_1 _4488_ (.A1(_0828_),
    .A2(_1177_),
    .B1_N(_1175_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1327_));
 sky130_fd_sc_hd__o2bb2a_1 _4489_ (.A1_N(_0828_),
    .A2_N(_1178_),
    .B1(_1327_),
    .B2(_0827_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1328_));
 sky130_fd_sc_hd__a21oi_1 _4490_ (.A1(_1326_),
    .A2(_1328_),
    .B1(_0847_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1329_));
 sky130_fd_sc_hd__a311o_1 _4491_ (.A1(_0846_),
    .A2(_1322_),
    .A3(_1323_),
    .B1(_1125_),
    .C1(_1329_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1330_));
 sky130_fd_sc_hd__o21ai_1 _4492_ (.A1(_1030_),
    .A2(_1299_),
    .B1(_1125_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1331_));
 sky130_fd_sc_hd__a21o_1 _4493_ (.A1(_1030_),
    .A2(_1280_),
    .B1(_1331_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1332_));
 sky130_fd_sc_hd__and3_1 _4494_ (.A(\i_tinyqv.cpu.instr_data_start[22] ),
    .B(\i_tinyqv.cpu.instr_data_start[21] ),
    .C(_0900_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1333_));
 sky130_fd_sc_hd__a21oi_1 _4495_ (.A1(\i_tinyqv.cpu.instr_data_start[21] ),
    .A2(_0900_),
    .B1(\i_tinyqv.cpu.instr_data_start[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1334_));
 sky130_fd_sc_hd__nor2_1 _4496_ (.A(_1333_),
    .B(_1334_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1335_));
 sky130_fd_sc_hd__nand2_1 _4497_ (.A(_0610_),
    .B(_1335_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1336_));
 sky130_fd_sc_hd__nor2_1 _4498_ (.A(\i_tinyqv.cpu.instr_data_start[14] ),
    .B(_0895_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1337_));
 sky130_fd_sc_hd__nor2_1 _4499_ (.A(_0896_),
    .B(_1337_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1338_));
 sky130_fd_sc_hd__xnor2_4 _4500_ (.A(_0887_),
    .B(_1206_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1339_));
 sky130_fd_sc_hd__xnor2_1 _4501_ (.A(_0883_),
    .B(_0890_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1340_));
 sky130_fd_sc_hd__a21oi_1 _4502_ (.A1(_0882_),
    .A2(_0892_),
    .B1(\i_tinyqv.cpu.instr_data_start[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1341_));
 sky130_fd_sc_hd__or2_1 _4503_ (.A(_0893_),
    .B(_1341_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1342_));
 sky130_fd_sc_hd__o22ai_1 _4504_ (.A1(_0609_),
    .A2(_1340_),
    .B1(_1342_),
    .B2(_0909_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1343_));
 sky130_fd_sc_hd__a221o_1 _4505_ (.A1(_0617_),
    .A2(_1338_),
    .B1(_1339_),
    .B2(_0689_),
    .C1(_1343_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1344_));
 sky130_fd_sc_hd__xnor2_1 _4506_ (.A(_0784_),
    .B(_0898_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1345_));
 sky130_fd_sc_hd__o2bb2a_1 _4507_ (.A1_N(_0752_),
    .A2_N(_1344_),
    .B1(_1345_),
    .B2(_0916_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1346_));
 sky130_fd_sc_hd__a21o_1 _4508_ (.A1(_1336_),
    .A2(_1346_),
    .B1(_0858_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1347_));
 sky130_fd_sc_hd__or2_2 _4509_ (.A(_0933_),
    .B(_0930_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1348_));
 sky130_fd_sc_hd__nor2_1 _4510_ (.A(_0946_),
    .B(_1348_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1349_));
 sky130_fd_sc_hd__a21oi_1 _4511_ (.A1(_0946_),
    .A2(_0841_),
    .B1(_0934_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1350_));
 sky130_fd_sc_hd__mux2_1 _4512_ (.A0(\i_tinyqv.cpu.i_core.time_hi[1] ),
    .A1(\i_tinyqv.cpu.i_core.cycle_count_wide[5] ),
    .S(_0841_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1351_));
 sky130_fd_sc_hd__a22o_1 _4513_ (.A1(\i_tinyqv.cpu.i_core.cycle_count[2] ),
    .A2(_0931_),
    .B1(_1351_),
    .B2(_0927_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1352_));
 sky130_fd_sc_hd__a211o_1 _4514_ (.A1(\i_tinyqv.cpu.i_core.i_instrret.data[2] ),
    .A2(_0929_),
    .B1(_1350_),
    .C1(_1352_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1353_));
 sky130_fd_sc_hd__a221o_1 _4515_ (.A1(\i_tinyqv.cpu.i_core.mepc[2] ),
    .A2(net19),
    .B1(_1349_),
    .B2(\i_tinyqv.cpu.i_core.mstatus_mte ),
    .C1(_1353_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1354_));
 sky130_fd_sc_hd__a221o_1 _4516_ (.A1(\i_tinyqv.cpu.i_core.mie[18] ),
    .A2(_0944_),
    .B1(_1228_),
    .B2(net15),
    .C1(_1354_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1355_));
 sky130_fd_sc_hd__a21oi_1 _4517_ (.A1(_0921_),
    .A2(_1355_),
    .B1(_0880_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1356_));
 sky130_fd_sc_hd__a22o_1 _4518_ (.A1(_0814_),
    .A2(_0880_),
    .B1(_1347_),
    .B2(_1356_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1357_));
 sky130_fd_sc_hd__a221o_1 _4519_ (.A1(\i_tinyqv.mem.data_from_read[18] ),
    .A2(_0689_),
    .B1(_0748_),
    .B2(\i_tinyqv.mem.data_from_read[22] ),
    .C1(_0957_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1358_));
 sky130_fd_sc_hd__mux2_1 _4520_ (.A0(\i_tinyqv.mem.qspi_data_buf[26] ),
    .A1(\i_tinyqv.mem.qspi_data_buf[30] ),
    .S(_0974_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1359_));
 sky130_fd_sc_hd__mux2_1 _4521_ (.A0(\i_tinyqv.cpu.instr_data_in[10] ),
    .A1(\i_tinyqv.cpu.instr_data_in[14] ),
    .S(_0838_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1360_));
 sky130_fd_sc_hd__mux2_1 _4522_ (.A0(_1359_),
    .A1(_1360_),
    .S(_0979_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1361_));
 sky130_fd_sc_hd__a22o_1 _4523_ (.A1(_0971_),
    .A2(_1358_),
    .B1(_1361_),
    .B2(_0973_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1362_));
 sky130_fd_sc_hd__and2_1 _4524_ (.A(_1001_),
    .B(uo_out[6]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1363_));
 sky130_fd_sc_hd__a221o_1 _4525_ (.A1(net8),
    .A2(_0986_),
    .B1(net14),
    .B2(\gpio_out_sel[6] ),
    .C1(_1363_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1364_));
 sky130_fd_sc_hd__a221o_1 _4526_ (.A1(\i_spi.data[6] ),
    .A2(_1000_),
    .B1(_0997_),
    .B2(\i_uart_rx.recieved_data[6] ),
    .C1(_0908_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1365_));
 sky130_fd_sc_hd__a221o_1 _4527_ (.A1(\i_uart_rx.recieved_data[2] ),
    .A2(_0996_),
    .B1(net14),
    .B2(\gpio_out_sel[2] ),
    .C1(_0974_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1366_));
 sky130_fd_sc_hd__a22o_1 _4528_ (.A1(\i_spi.data[2] ),
    .A2(_1000_),
    .B1(_1001_),
    .B2(uo_out[2]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1367_));
 sky130_fd_sc_hd__a211o_1 _4529_ (.A1(net4),
    .A2(_0986_),
    .B1(_1366_),
    .C1(_1367_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1368_));
 sky130_fd_sc_hd__o211a_1 _4530_ (.A1(_1364_),
    .A2(_1365_),
    .B1(_1368_),
    .C1(_0945_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1369_));
 sky130_fd_sc_hd__mux2_1 _4531_ (.A0(\i_tinyqv.cpu.instr_data_in[14] ),
    .A1(\i_tinyqv.mem.qspi_data_buf[14] ),
    .S(_1017_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1370_));
 sky130_fd_sc_hd__mux2_1 _4532_ (.A0(\i_tinyqv.cpu.instr_data_in[10] ),
    .A1(\i_tinyqv.mem.qspi_data_buf[10] ),
    .S(_1017_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1371_));
 sky130_fd_sc_hd__mux2_1 _4533_ (.A0(\i_tinyqv.cpu.instr_data_in[2] ),
    .A1(\i_tinyqv.cpu.instr_data_in[6] ),
    .S(_0838_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1372_));
 sky130_fd_sc_hd__mux2_1 _4534_ (.A0(_1360_),
    .A1(_1372_),
    .S(_1012_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1373_));
 sky130_fd_sc_hd__o22a_1 _4535_ (.A1(_0909_),
    .A2(_1371_),
    .B1(_1373_),
    .B2(_0907_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1374_));
 sky130_fd_sc_hd__o21a_1 _4536_ (.A1(_0724_),
    .A2(_1370_),
    .B1(_1374_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1375_));
 sky130_fd_sc_hd__o22a_1 _4537_ (.A1(_0982_),
    .A2(_1369_),
    .B1(_1375_),
    .B2(_0957_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1376_));
 sky130_fd_sc_hd__a21oi_1 _4538_ (.A1(_0956_),
    .A2(_1362_),
    .B1(_1376_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1377_));
 sky130_fd_sc_hd__o21ba_1 _4539_ (.A1(_1022_),
    .A2(_1377_),
    .B1_N(_1023_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1378_));
 sky130_fd_sc_hd__a21oi_1 _4540_ (.A1(_0878_),
    .A2(_1357_),
    .B1(_1378_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1379_));
 sky130_fd_sc_hd__a32o_2 _4541_ (.A1(_1034_),
    .A2(_1330_),
    .A3(_1332_),
    .B1(_1379_),
    .B2(_0877_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1380_));
 sky130_fd_sc_hd__buf_4 _4542_ (.A(_1380_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.debug_rd[2] ));
 sky130_fd_sc_hd__mux2_1 _4543_ (.A0(net104),
    .A1(\i_tinyqv.cpu.debug_rd[2] ),
    .S(_1190_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1381_));
 sky130_fd_sc_hd__clkbuf_1 _4544_ (.A(_1381_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0052_));
 sky130_fd_sc_hd__mux2_1 _4545_ (.A0(\i_spi.data[7] ),
    .A1(\debug_rd_r[1] ),
    .S(debug_register_data),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1382_));
 sky130_fd_sc_hd__mux2_1 _4546_ (.A0(_1382_),
    .A1(\gpio_out[3] ),
    .S(\gpio_out_sel[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1383_));
 sky130_fd_sc_hd__clkbuf_4 _4547_ (.A(_1383_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[3]));
 sky130_fd_sc_hd__inv_2 _4548_ (.A(net7),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1384_));
 sky130_fd_sc_hd__inv_2 _4549_ (.A(\i_tinyqv.cpu.data_continue ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1385_));
 sky130_fd_sc_hd__nand2_2 _4550_ (.A(_0688_),
    .B(_0907_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1386_));
 sky130_fd_sc_hd__nor2_2 _4551_ (.A(_0908_),
    .B(_1386_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1387_));
 sky130_fd_sc_hd__inv_2 _4552_ (.A(\i_tinyqv.cpu.i_core.mem_op[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1388_));
 sky130_fd_sc_hd__a21oi_1 _4553_ (.A1(_0826_),
    .A2(_0835_),
    .B1(_1388_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1389_));
 sky130_fd_sc_hd__nand2_4 _4554_ (.A(_0653_),
    .B(\i_tinyqv.cpu.is_branch ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1390_));
 sky130_fd_sc_hd__a31o_1 _4555_ (.A1(_1388_),
    .A2(_0826_),
    .A3(_0835_),
    .B1(_1390_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1391_));
 sky130_fd_sc_hd__nor2_2 _4556_ (.A(_0855_),
    .B(_1173_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1392_));
 sky130_fd_sc_hd__nand3_1 _4557_ (.A(\i_tinyqv.cpu.i_core.imm_lo[8] ),
    .B(\i_tinyqv.cpu.i_core.imm_lo[9] ),
    .C(_1392_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1393_));
 sky130_fd_sc_hd__nor2_1 _4558_ (.A(\i_tinyqv.cpu.i_core.imm_lo[8] ),
    .B(\i_tinyqv.cpu.i_core.imm_lo[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1394_));
 sky130_fd_sc_hd__a21oi_2 _4559_ (.A1(_1394_),
    .A2(_1392_),
    .B1(\i_tinyqv.cpu.i_core.is_interrupt ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1395_));
 sky130_fd_sc_hd__and3_1 _4560_ (.A(_0858_),
    .B(_1393_),
    .C(_1395_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1396_));
 sky130_fd_sc_hd__o21ai_2 _4561_ (.A1(_1389_),
    .A2(_1391_),
    .B1(_1396_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1397_));
 sky130_fd_sc_hd__and2_4 _4562_ (.A(_1387_),
    .B(_1397_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1398_));
 sky130_fd_sc_hd__buf_8 _4563_ (.A(_1398_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1399_));
 sky130_fd_sc_hd__clkinv_4 _4564_ (.A(\i_tinyqv.cpu.i_core.i_cycles.rstn ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1400_));
 sky130_fd_sc_hd__a22o_1 _4565_ (.A1(\i_tinyqv.cpu.i_core.mie[16] ),
    .A2(\i_tinyqv.cpu.i_core.mip[16] ),
    .B1(\i_tinyqv.cpu.i_core.mip[17] ),
    .B2(\i_tinyqv.cpu.i_core.mie[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1401_));
 sky130_fd_sc_hd__a21oi_1 _4566_ (.A1(\i_tinyqv.cpu.i_core.mie[18] ),
    .A2(_1228_),
    .B1(_1401_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1402_));
 sky130_fd_sc_hd__nand2_1 _4567_ (.A(\i_tinyqv.cpu.i_core.mie[19] ),
    .B(_0991_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1403_));
 sky130_fd_sc_hd__a21bo_1 _4568_ (.A1(_1402_),
    .A2(_1403_),
    .B1_N(\i_tinyqv.cpu.i_core.mstatus_mie ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1404_));
 sky130_fd_sc_hd__nor2_1 _4569_ (.A(_0862_),
    .B(_1404_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1405_));
 sky130_fd_sc_hd__buf_2 _4570_ (.A(\i_tinyqv.cpu.instr_write_offset[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1406_));
 sky130_fd_sc_hd__inv_2 _4571_ (.A(_0749_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1407_));
 sky130_fd_sc_hd__mux2_4 _4572_ (.A0(_1407_),
    .A1(_1208_),
    .S(_0653_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1408_));
 sky130_fd_sc_hd__buf_4 _4573_ (.A(_1408_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1409_));
 sky130_fd_sc_hd__inv_2 _4574_ (.A(\i_tinyqv.cpu.debug_instr_valid ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1410_));
 sky130_fd_sc_hd__or2_2 _4575_ (.A(\i_tinyqv.cpu.debug_instr_valid ),
    .B(\i_tinyqv.cpu.pc[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1411_));
 sky130_fd_sc_hd__o21a_4 _4576_ (.A1(_1410_),
    .A2(_1339_),
    .B1(_1411_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1412_));
 sky130_fd_sc_hd__mux2_1 _4577_ (.A0(\i_tinyqv.cpu.instr_data[0][0] ),
    .A1(\i_tinyqv.cpu.instr_data[2][0] ),
    .S(net36),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1413_));
 sky130_fd_sc_hd__clkbuf_4 _4578_ (.A(_1412_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1414_));
 sky130_fd_sc_hd__inv_2 _4579_ (.A(_1208_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1415_));
 sky130_fd_sc_hd__mux2_4 _4580_ (.A0(_0749_),
    .A1(_1415_),
    .S(_0653_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1416_));
 sky130_fd_sc_hd__o21ai_2 _4581_ (.A1(_1410_),
    .A2(net325),
    .B1(_1411_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1417_));
 sky130_fd_sc_hd__or2_1 _4582_ (.A(\i_tinyqv.cpu.instr_data[3][0] ),
    .B(_1417_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1418_));
 sky130_fd_sc_hd__o211a_1 _4583_ (.A1(\i_tinyqv.cpu.instr_data[1][0] ),
    .A2(_1414_),
    .B1(_1416_),
    .C1(_1418_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1419_));
 sky130_fd_sc_hd__a21oi_4 _4584_ (.A1(_1409_),
    .A2(_1413_),
    .B1(_1419_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1420_));
 sky130_fd_sc_hd__or2_1 _4585_ (.A(\i_tinyqv.cpu.instr_data[1][1] ),
    .B(_1414_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1421_));
 sky130_fd_sc_hd__buf_2 _4586_ (.A(_1417_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1422_));
 sky130_fd_sc_hd__or2_2 _4587_ (.A(\i_tinyqv.cpu.instr_data[3][1] ),
    .B(_1422_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1423_));
 sky130_fd_sc_hd__or2_1 _4588_ (.A(\i_tinyqv.cpu.instr_data[0][1] ),
    .B(net36),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1424_));
 sky130_fd_sc_hd__o211a_1 _4589_ (.A1(\i_tinyqv.cpu.instr_data[2][1] ),
    .A2(_1422_),
    .B1(_1408_),
    .C1(_1424_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1425_));
 sky130_fd_sc_hd__a31oi_4 _4590_ (.A1(_1416_),
    .A2(_1421_),
    .A3(_1423_),
    .B1(_1425_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1426_));
 sky130_fd_sc_hd__or2_2 _4591_ (.A(_1420_),
    .B(_1426_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1427_));
 sky130_fd_sc_hd__nand2_1 _4592_ (.A(_0653_),
    .B(_0888_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1428_));
 sky130_fd_sc_hd__xnor2_1 _4593_ (.A(\i_tinyqv.cpu.instr_write_offset[3] ),
    .B(_1428_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1429_));
 sky130_fd_sc_hd__a21o_1 _4594_ (.A1(\i_tinyqv.cpu.instr_write_offset[2] ),
    .A2(_1422_),
    .B1(_1429_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1430_));
 sky130_fd_sc_hd__o31a_1 _4595_ (.A1(_1406_),
    .A2(_1409_),
    .A3(_1427_),
    .B1(_1430_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1431_));
 sky130_fd_sc_hd__buf_4 _4596_ (.A(_1409_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1432_));
 sky130_fd_sc_hd__or2_1 _4597_ (.A(\i_tinyqv.cpu.instr_write_offset[2] ),
    .B(_1422_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1433_));
 sky130_fd_sc_hd__o21a_1 _4598_ (.A1(_1406_),
    .A2(_1409_),
    .B1(_1433_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1434_));
 sky130_fd_sc_hd__a2bb2o_1 _4599_ (.A1_N(_1430_),
    .A2_N(_1434_),
    .B1(_1433_),
    .B2(_1429_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1435_));
 sky130_fd_sc_hd__a31o_1 _4600_ (.A1(_1406_),
    .A2(_1432_),
    .A3(_1427_),
    .B1(_1435_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1436_));
 sky130_fd_sc_hd__inv_2 _4601_ (.A(\i_tinyqv.cpu.was_early_branch ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1437_));
 sky130_fd_sc_hd__o21ai_2 _4602_ (.A1(_1431_),
    .A2(_1436_),
    .B1(_1437_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1438_));
 sky130_fd_sc_hd__nand2_1 _4603_ (.A(_0837_),
    .B(_0863_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1439_));
 sky130_fd_sc_hd__or3_2 _4604_ (.A(\i_tinyqv.cpu.additional_mem_ops[2] ),
    .B(\i_tinyqv.cpu.additional_mem_ops[1] ),
    .C(\i_tinyqv.cpu.additional_mem_ops[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1440_));
 sky130_fd_sc_hd__or2_1 _4605_ (.A(_1439_),
    .B(_1440_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1441_));
 sky130_fd_sc_hd__buf_2 _4606_ (.A(_1441_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1442_));
 sky130_fd_sc_hd__o21ai_1 _4607_ (.A1(_0653_),
    .A2(_0841_),
    .B1(_1442_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1443_));
 sky130_fd_sc_hd__or4b_1 _4608_ (.A(_1400_),
    .B(_1405_),
    .C(_1438_),
    .D_N(_1443_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1444_));
 sky130_fd_sc_hd__or2_1 _4609_ (.A(\i_tinyqv.cpu.instr_data[3][3] ),
    .B(_1422_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1445_));
 sky130_fd_sc_hd__o21a_1 _4610_ (.A1(\i_tinyqv.cpu.instr_data[1][3] ),
    .A2(_1414_),
    .B1(_1416_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1446_));
 sky130_fd_sc_hd__mux2_1 _4611_ (.A0(\i_tinyqv.cpu.instr_data[0][3] ),
    .A1(\i_tinyqv.cpu.instr_data[2][3] ),
    .S(_1412_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1447_));
 sky130_fd_sc_hd__a22o_1 _4612_ (.A1(_1445_),
    .A2(_1446_),
    .B1(_1447_),
    .B2(_1408_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1448_));
 sky130_fd_sc_hd__clkbuf_4 _4613_ (.A(_1414_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1449_));
 sky130_fd_sc_hd__mux2_1 _4614_ (.A0(\i_tinyqv.cpu.instr_data[1][5] ),
    .A1(\i_tinyqv.cpu.instr_data[3][5] ),
    .S(_1449_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1450_));
 sky130_fd_sc_hd__mux2_1 _4615_ (.A0(\i_tinyqv.cpu.instr_data[0][5] ),
    .A1(\i_tinyqv.cpu.instr_data[2][5] ),
    .S(_1449_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1451_));
 sky130_fd_sc_hd__mux2_2 _4616_ (.A0(_1450_),
    .A1(_1451_),
    .S(_1409_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1452_));
 sky130_fd_sc_hd__mux2_1 _4617_ (.A0(\i_tinyqv.cpu.instr_data[1][6] ),
    .A1(\i_tinyqv.cpu.instr_data[3][6] ),
    .S(_1414_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1453_));
 sky130_fd_sc_hd__mux2_1 _4618_ (.A0(\i_tinyqv.cpu.instr_data[0][6] ),
    .A1(\i_tinyqv.cpu.instr_data[2][6] ),
    .S(_1414_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1454_));
 sky130_fd_sc_hd__mux2_2 _4619_ (.A0(_1453_),
    .A1(_1454_),
    .S(_1409_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1455_));
 sky130_fd_sc_hd__nand2_1 _4620_ (.A(_1452_),
    .B(_1455_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1456_));
 sky130_fd_sc_hd__or2_1 _4621_ (.A(\i_tinyqv.cpu.instr_data[3][2] ),
    .B(_1422_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1457_));
 sky130_fd_sc_hd__o21a_1 _4622_ (.A1(\i_tinyqv.cpu.instr_data[1][2] ),
    .A2(_1414_),
    .B1(_1416_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1458_));
 sky130_fd_sc_hd__mux2_1 _4623_ (.A0(\i_tinyqv.cpu.instr_data[0][2] ),
    .A1(\i_tinyqv.cpu.instr_data[2][2] ),
    .S(_1412_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1459_));
 sky130_fd_sc_hd__a22o_4 _4624_ (.A1(_1457_),
    .A2(_1458_),
    .B1(_1459_),
    .B2(_1408_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1460_));
 sky130_fd_sc_hd__buf_4 _4625_ (.A(_1416_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1461_));
 sky130_fd_sc_hd__mux2_1 _4626_ (.A0(\i_tinyqv.cpu.instr_data[1][4] ),
    .A1(\i_tinyqv.cpu.instr_data[3][4] ),
    .S(_1414_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1462_));
 sky130_fd_sc_hd__or2_1 _4627_ (.A(\i_tinyqv.cpu.instr_data[2][4] ),
    .B(_1422_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1463_));
 sky130_fd_sc_hd__o211a_1 _4628_ (.A1(\i_tinyqv.cpu.instr_data[0][4] ),
    .A2(_1414_),
    .B1(_1409_),
    .C1(_1463_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1464_));
 sky130_fd_sc_hd__a21oi_1 _4629_ (.A1(_1461_),
    .A2(_1462_),
    .B1(_1464_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1465_));
 sky130_fd_sc_hd__and3b_1 _4630_ (.A_N(_1456_),
    .B(_1460_),
    .C(_1465_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1466_));
 sky130_fd_sc_hd__nand2_1 _4631_ (.A(_1448_),
    .B(_1466_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1467_));
 sky130_fd_sc_hd__a31o_2 _4632_ (.A1(_1461_),
    .A2(_1421_),
    .A3(_1423_),
    .B1(_1425_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1468_));
 sky130_fd_sc_hd__or2_1 _4633_ (.A(_1420_),
    .B(_1468_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1469_));
 sky130_fd_sc_hd__mux2_2 _4634_ (.A0(\i_tinyqv.cpu.instr_data[1][13] ),
    .A1(\i_tinyqv.cpu.instr_data[3][13] ),
    .S(net36),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1470_));
 sky130_fd_sc_hd__or2_1 _4635_ (.A(\i_tinyqv.cpu.instr_data[2][13] ),
    .B(_1417_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1471_));
 sky130_fd_sc_hd__o211a_1 _4636_ (.A1(\i_tinyqv.cpu.instr_data[0][13] ),
    .A2(_1414_),
    .B1(_1408_),
    .C1(_1471_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1472_));
 sky130_fd_sc_hd__a21oi_4 _4637_ (.A1(_1461_),
    .A2(_1470_),
    .B1(_1472_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1473_));
 sky130_fd_sc_hd__mux2_1 _4638_ (.A0(\i_tinyqv.cpu.instr_data[1][14] ),
    .A1(\i_tinyqv.cpu.instr_data[3][14] ),
    .S(net322),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1474_));
 sky130_fd_sc_hd__mux2_1 _4639_ (.A0(\i_tinyqv.cpu.instr_data[0][14] ),
    .A1(\i_tinyqv.cpu.instr_data[2][14] ),
    .S(net322),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1475_));
 sky130_fd_sc_hd__mux2_4 _4640_ (.A0(_1474_),
    .A1(_1475_),
    .S(_1408_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1476_));
 sky130_fd_sc_hd__or2_2 _4641_ (.A(_1473_),
    .B(_1476_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1477_));
 sky130_fd_sc_hd__nor2_2 _4642_ (.A(_1469_),
    .B(_1477_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1478_));
 sky130_fd_sc_hd__o21ba_1 _4643_ (.A1(_1427_),
    .A2(_1467_),
    .B1_N(_1478_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1479_));
 sky130_fd_sc_hd__nor3_4 _4644_ (.A(_1399_),
    .B(_1444_),
    .C(_1479_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1480_));
 sky130_fd_sc_hd__a21o_1 _4645_ (.A1(_1416_),
    .A2(_1470_),
    .B1(_1472_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1481_));
 sky130_fd_sc_hd__or2_1 _4646_ (.A(_1481_),
    .B(_1476_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1482_));
 sky130_fd_sc_hd__buf_4 _4647_ (.A(_1482_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1483_));
 sky130_fd_sc_hd__mux2_1 _4648_ (.A0(\i_tinyqv.cpu.instr_data[1][15] ),
    .A1(\i_tinyqv.cpu.instr_data[3][15] ),
    .S(net35),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1484_));
 sky130_fd_sc_hd__mux2_1 _4649_ (.A0(\i_tinyqv.cpu.instr_data[0][15] ),
    .A1(\i_tinyqv.cpu.instr_data[2][15] ),
    .S(net34),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1485_));
 sky130_fd_sc_hd__mux2_4 _4650_ (.A0(_1484_),
    .A1(_1485_),
    .S(_1408_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1486_));
 sky130_fd_sc_hd__nand2_1 _4651_ (.A(_1420_),
    .B(_1486_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1487_));
 sky130_fd_sc_hd__or2_1 _4652_ (.A(_1426_),
    .B(_1487_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1488_));
 sky130_fd_sc_hd__or2_1 _4653_ (.A(_1483_),
    .B(_1488_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1489_));
 sky130_fd_sc_hd__clkbuf_2 _4654_ (.A(_1489_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1490_));
 sky130_fd_sc_hd__a21o_2 _4655_ (.A1(_1416_),
    .A2(_1462_),
    .B1(_1464_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1491_));
 sky130_fd_sc_hd__or2_1 _4656_ (.A(_1448_),
    .B(_1460_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1492_));
 sky130_fd_sc_hd__or3_4 _4657_ (.A(_1455_),
    .B(_1491_),
    .C(_1492_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1493_));
 sky130_fd_sc_hd__or2_1 _4658_ (.A(_1452_),
    .B(_1493_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1494_));
 sky130_fd_sc_hd__or2_4 _4659_ (.A(_1490_),
    .B(_1494_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1495_));
 sky130_fd_sc_hd__mux2_1 _4660_ (.A0(\i_tinyqv.cpu.instr_data[1][10] ),
    .A1(\i_tinyqv.cpu.instr_data[3][10] ),
    .S(_1449_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1496_));
 sky130_fd_sc_hd__mux2_1 _4661_ (.A0(\i_tinyqv.cpu.instr_data[0][10] ),
    .A1(\i_tinyqv.cpu.instr_data[2][10] ),
    .S(_1449_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1497_));
 sky130_fd_sc_hd__mux2_1 _4662_ (.A0(_1496_),
    .A1(_1497_),
    .S(_1409_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1498_));
 sky130_fd_sc_hd__mux2_1 _4663_ (.A0(\i_tinyqv.cpu.instr_data[1][9] ),
    .A1(\i_tinyqv.cpu.instr_data[3][9] ),
    .S(_1449_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1499_));
 sky130_fd_sc_hd__mux2_1 _4664_ (.A0(\i_tinyqv.cpu.instr_data[0][9] ),
    .A1(\i_tinyqv.cpu.instr_data[2][9] ),
    .S(_1449_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1500_));
 sky130_fd_sc_hd__mux2_2 _4665_ (.A0(_1499_),
    .A1(_1500_),
    .S(_1409_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1501_));
 sky130_fd_sc_hd__or2_1 _4666_ (.A(_1498_),
    .B(_1501_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1502_));
 sky130_fd_sc_hd__mux2_1 _4667_ (.A0(\i_tinyqv.cpu.instr_data[1][12] ),
    .A1(\i_tinyqv.cpu.instr_data[3][12] ),
    .S(_1449_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1503_));
 sky130_fd_sc_hd__clkbuf_4 _4668_ (.A(_1449_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1504_));
 sky130_fd_sc_hd__or2_1 _4669_ (.A(\i_tinyqv.cpu.instr_data[2][12] ),
    .B(_1422_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1505_));
 sky130_fd_sc_hd__o211a_1 _4670_ (.A1(\i_tinyqv.cpu.instr_data[0][12] ),
    .A2(_1504_),
    .B1(_1409_),
    .C1(_1505_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1506_));
 sky130_fd_sc_hd__a21oi_4 _4671_ (.A1(_1461_),
    .A2(_1503_),
    .B1(_1506_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1507_));
 sky130_fd_sc_hd__mux2_1 _4672_ (.A0(\i_tinyqv.cpu.instr_data[1][7] ),
    .A1(\i_tinyqv.cpu.instr_data[3][7] ),
    .S(_1449_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1508_));
 sky130_fd_sc_hd__mux2_1 _4673_ (.A0(\i_tinyqv.cpu.instr_data[0][7] ),
    .A1(\i_tinyqv.cpu.instr_data[2][7] ),
    .S(_1449_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1509_));
 sky130_fd_sc_hd__mux2_4 _4674_ (.A0(_1508_),
    .A1(_1509_),
    .S(_1432_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1510_));
 sky130_fd_sc_hd__nand2_1 _4675_ (.A(_1507_),
    .B(_1510_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1511_));
 sky130_fd_sc_hd__mux2_1 _4676_ (.A0(\i_tinyqv.cpu.instr_data[1][8] ),
    .A1(\i_tinyqv.cpu.instr_data[3][8] ),
    .S(_1504_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1512_));
 sky130_fd_sc_hd__mux2_1 _4677_ (.A0(\i_tinyqv.cpu.instr_data[0][8] ),
    .A1(\i_tinyqv.cpu.instr_data[2][8] ),
    .S(_1504_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1513_));
 sky130_fd_sc_hd__mux2_4 _4678_ (.A0(_1512_),
    .A1(_1513_),
    .S(_1432_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1514_));
 sky130_fd_sc_hd__or4_4 _4679_ (.A(_1495_),
    .B(_1502_),
    .C(_1511_),
    .D(_1514_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1515_));
 sky130_fd_sc_hd__nor3_4 _4680_ (.A(_1399_),
    .B(_1444_),
    .C(_1515_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1516_));
 sky130_fd_sc_hd__a31o_1 _4681_ (.A1(_1437_),
    .A2(_1387_),
    .A3(net33),
    .B1(\i_tinyqv.cpu.instr_fetch_running ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1517_));
 sky130_fd_sc_hd__and3_1 _4682_ (.A(_0864_),
    .B(\i_tinyqv.mem.qspi_data_byte_idx[0] ),
    .C(\i_tinyqv.mem.q_ctrl.data_ready ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1518_));
 sky130_fd_sc_hd__and4_1 _4683_ (.A(\i_tinyqv.cpu.instr_fetch_running ),
    .B(\i_tinyqv.mem.instr_active ),
    .C(\i_tinyqv.cpu.instr_write_offset[1] ),
    .D(_1518_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1519_));
 sky130_fd_sc_hd__a31o_1 _4684_ (.A1(\i_tinyqv.cpu.instr_fetch_running ),
    .A2(\i_tinyqv.mem.instr_active ),
    .A3(_1518_),
    .B1(_1406_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1520_));
 sky130_fd_sc_hd__or2b_1 _4685_ (.A(_1519_),
    .B_N(_1520_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1521_));
 sky130_fd_sc_hd__nand2_1 _4686_ (.A(\i_tinyqv.cpu.instr_write_offset[2] ),
    .B(_1519_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1522_));
 sky130_fd_sc_hd__or2_1 _4687_ (.A(\i_tinyqv.cpu.instr_write_offset[2] ),
    .B(_1519_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1523_));
 sky130_fd_sc_hd__nand2_1 _4688_ (.A(_1522_),
    .B(_1523_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1524_));
 sky130_fd_sc_hd__o2bb2a_1 _4689_ (.A1_N(_0749_),
    .A2_N(_1521_),
    .B1(_1524_),
    .B2(net60),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1525_));
 sky130_fd_sc_hd__or3b_1 _4690_ (.A(_1439_),
    .B(_1440_),
    .C_N(_0888_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1526_));
 sky130_fd_sc_hd__xnor2_1 _4691_ (.A(\i_tinyqv.cpu.instr_write_offset[3] ),
    .B(_1522_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1527_));
 sky130_fd_sc_hd__xnor2_1 _4692_ (.A(_1526_),
    .B(_1527_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1528_));
 sky130_fd_sc_hd__a21boi_1 _4693_ (.A1(net60),
    .A2(_1524_),
    .B1_N(_1528_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1529_));
 sky130_fd_sc_hd__o211ai_2 _4694_ (.A1(_0749_),
    .A2(_1521_),
    .B1(_1525_),
    .C1(_1529_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1530_));
 sky130_fd_sc_hd__and2_1 _4695_ (.A(_0864_),
    .B(\i_tinyqv.mem.qspi_data_byte_idx[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1531_));
 sky130_fd_sc_hd__or4b_4 _4696_ (.A(_0978_),
    .B(_1530_),
    .C(\i_tinyqv.mem.q_ctrl.data_ready ),
    .D_N(_1531_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1532_));
 sky130_fd_sc_hd__and2_1 _4697_ (.A(\i_tinyqv.cpu.instr_fetch_started ),
    .B(_1532_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1533_));
 sky130_fd_sc_hd__or4_4 _4698_ (.A(_1480_),
    .B(_1516_),
    .C(_1517_),
    .D(_1533_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1534_));
 sky130_fd_sc_hd__inv_2 _4699_ (.A(_1518_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1535_));
 sky130_fd_sc_hd__a41o_2 _4700_ (.A1(\i_tinyqv.cpu.data_read_n[1] ),
    .A2(\i_tinyqv.cpu.data_read_n[0] ),
    .A3(\i_tinyqv.cpu.data_write_n[1] ),
    .A4(\i_tinyqv.cpu.data_write_n[0] ),
    .B1(_0865_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1536_));
 sky130_fd_sc_hd__a21o_1 _4701_ (.A1(_1535_),
    .A2(_1530_),
    .B1(_1536_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1537_));
 sky130_fd_sc_hd__o211a_1 _4702_ (.A1(\i_tinyqv.mem.q_ctrl.data_ready ),
    .A2(\i_tinyqv.mem.q_ctrl.data_req ),
    .B1(_1385_),
    .C1(_0872_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1538_));
 sky130_fd_sc_hd__or3_1 _4703_ (.A(\i_tinyqv.mem.q_ctrl.fsm_state[2] ),
    .B(\i_tinyqv.mem.q_ctrl.fsm_state[1] ),
    .C(\i_tinyqv.mem.q_ctrl.fsm_state[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1539_));
 sky130_fd_sc_hd__clkbuf_4 _4704_ (.A(_1539_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1540_));
 sky130_fd_sc_hd__or2_2 _4705_ (.A(\i_tinyqv.mem.qspi_write_done ),
    .B(_1540_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1541_));
 sky130_fd_sc_hd__o21ai_1 _4706_ (.A1(\i_tinyqv.mem.instr_active ),
    .A2(_1538_),
    .B1(_1541_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1542_));
 sky130_fd_sc_hd__a31o_4 _4707_ (.A1(\i_tinyqv.mem.instr_active ),
    .A2(_1534_),
    .A3(_1537_),
    .B1(_1542_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1543_));
 sky130_fd_sc_hd__inv_2 _4708_ (.A(net6),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1544_));
 sky130_fd_sc_hd__mux4_2 _4709_ (.A0(_1385_),
    .A1(_0946_),
    .A2(_1543_),
    .A3(_1532_),
    .S0(net5),
    .S1(_1544_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1545_));
 sky130_fd_sc_hd__buf_6 _4710_ (.A(_1516_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1546_));
 sky130_fd_sc_hd__mux4_1 _4711_ (.A0(_1188_),
    .A1(_1480_),
    .A2(_1546_),
    .A3(_1399_),
    .S0(net6),
    .S1(net5),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1547_));
 sky130_fd_sc_hd__nor2_1 _4712_ (.A(_1384_),
    .B(_1547_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1548_));
 sky130_fd_sc_hd__a211oi_2 _4713_ (.A1(_1384_),
    .A2(_1545_),
    .B1(_1548_),
    .C1(net8),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1549_));
 sky130_fd_sc_hd__or2_1 _4714_ (.A(_1480_),
    .B(_1546_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1550_));
 sky130_fd_sc_hd__or2_2 _4715_ (.A(_1550_),
    .B(_1517_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1551_));
 sky130_fd_sc_hd__buf_4 _4716_ (.A(_1518_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1552_));
 sky130_fd_sc_hd__nand2_1 _4717_ (.A(\i_tinyqv.mem.instr_active ),
    .B(_1552_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1553_));
 sky130_fd_sc_hd__mux4_1 _4718_ (.A0(_1551_),
    .A1(_1553_),
    .A2(_1410_),
    .A3(_1442_),
    .S0(net6),
    .S1(net5),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1554_));
 sky130_fd_sc_hd__inv_2 _4719_ (.A(_1404_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1555_));
 sky130_fd_sc_hd__or2_2 _4720_ (.A(_0865_),
    .B(_0979_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1556_));
 sky130_fd_sc_hd__a21oi_4 _4721_ (.A1(\i_tinyqv.cpu.data_write_n[1] ),
    .A2(\i_tinyqv.cpu.data_write_n[0] ),
    .B1(net28),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1557_));
 sky130_fd_sc_hd__a21oi_2 _4722_ (.A1(\i_tinyqv.cpu.data_read_n[1] ),
    .A2(\i_tinyqv.cpu.data_read_n[0] ),
    .B1(net28),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1558_));
 sky130_fd_sc_hd__mux4_1 _4723_ (.A0(_1555_),
    .A1(_1556_),
    .A2(_1557_),
    .A3(_1558_),
    .S0(net5),
    .S1(net6),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1559_));
 sky130_fd_sc_hd__o21ai_1 _4724_ (.A1(net7),
    .A2(_1559_),
    .B1(net8),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1560_));
 sky130_fd_sc_hd__a21oi_1 _4725_ (.A1(net7),
    .A2(_1554_),
    .B1(_1560_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1561_));
 sky130_fd_sc_hd__or2b_1 _4726_ (.A(\gpio_out[7] ),
    .B_N(\gpio_out_sel[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1562_));
 sky130_fd_sc_hd__o31a_4 _4727_ (.A1(\gpio_out_sel[7] ),
    .A2(_1549_),
    .A3(_1561_),
    .B1(_1562_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[7]));
 sky130_fd_sc_hd__nand2_2 _4728_ (.A(_0656_),
    .B(\i_tinyqv.cpu.alu_op[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1563_));
 sky130_fd_sc_hd__and2b_1 _4729_ (.A_N(_0823_),
    .B(_1178_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1564_));
 sky130_fd_sc_hd__nand2_1 _4730_ (.A(_0817_),
    .B(_1324_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1565_));
 sky130_fd_sc_hd__nand2_1 _4731_ (.A(_0701_),
    .B(_0820_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1566_));
 sky130_fd_sc_hd__xor2_1 _4732_ (.A(_1565_),
    .B(_1566_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1567_));
 sky130_fd_sc_hd__o22ai_1 _4733_ (.A1(_0824_),
    .A2(_1177_),
    .B1(_1567_),
    .B2(_1173_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1568_));
 sky130_fd_sc_hd__a211o_1 _4734_ (.A1(_0822_),
    .A2(_1175_),
    .B1(_1564_),
    .C1(_1568_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1569_));
 sky130_fd_sc_hd__and2_1 _4735_ (.A(\i_tinyqv.cpu.i_core.multiplier.accum[2] ),
    .B(_1316_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1570_));
 sky130_fd_sc_hd__o311a_1 _4736_ (.A1(_0636_),
    .A2(_0641_),
    .A3(net71),
    .B1(\i_tinyqv.cpu.i_core.i_shift.a[0] ),
    .C1(\i_tinyqv.cpu.i_core.cycle[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1571_));
 sky130_fd_sc_hd__o211a_1 _4737_ (.A1(net76),
    .A2(_0797_),
    .B1(\i_tinyqv.cpu.i_core.cycle[0] ),
    .C1(\i_tinyqv.cpu.i_core.i_shift.a[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1572_));
 sky130_fd_sc_hd__xnor2_2 _4738_ (.A(_1571_),
    .B(_1572_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1573_));
 sky130_fd_sc_hd__nand2_1 _4739_ (.A(\i_tinyqv.cpu.i_core.i_shift.a[3] ),
    .B(_1166_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1574_));
 sky130_fd_sc_hd__xor2_2 _4740_ (.A(_1573_),
    .B(_1574_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1575_));
 sky130_fd_sc_hd__xnor2_2 _4741_ (.A(_1315_),
    .B(_1575_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1576_));
 sky130_fd_sc_hd__xor2_2 _4742_ (.A(\i_tinyqv.cpu.i_core.multiplier.accum[3] ),
    .B(_1576_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1577_));
 sky130_fd_sc_hd__xnor2_2 _4743_ (.A(_1570_),
    .B(_1577_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1578_));
 sky130_fd_sc_hd__nand2_1 _4744_ (.A(\i_tinyqv.cpu.i_core.i_shift.a[2] ),
    .B(_1250_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1579_));
 sky130_fd_sc_hd__xor2_1 _4745_ (.A(_1578_),
    .B(_1579_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1580_));
 sky130_fd_sc_hd__or2_1 _4746_ (.A(_1308_),
    .B(_1317_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1581_));
 sky130_fd_sc_hd__o21ai_1 _4747_ (.A1(_1318_),
    .A2(_1319_),
    .B1(_1581_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1582_));
 sky130_fd_sc_hd__xor2_1 _4748_ (.A(_1580_),
    .B(_1582_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1583_));
 sky130_fd_sc_hd__xor2_1 _4749_ (.A(_1322_),
    .B(net82),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1584_));
 sky130_fd_sc_hd__nor2_1 _4750_ (.A(_1563_),
    .B(_1584_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1585_));
 sky130_fd_sc_hd__a211o_1 _4751_ (.A1(_1563_),
    .A2(_1569_),
    .B1(_1585_),
    .C1(_1125_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1586_));
 sky130_fd_sc_hd__mux2_1 _4752_ (.A0(_1122_),
    .A1(_1163_),
    .S(_1030_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1587_));
 sky130_fd_sc_hd__nand2_1 _4753_ (.A(_1125_),
    .B(_1587_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1588_));
 sky130_fd_sc_hd__clkbuf_4 _4754_ (.A(_0617_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1589_));
 sky130_fd_sc_hd__xnor2_1 _4755_ (.A(_0881_),
    .B(_0896_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1590_));
 sky130_fd_sc_hd__xor2_1 _4756_ (.A(_0884_),
    .B(_0888_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1591_));
 sky130_fd_sc_hd__a21oi_1 _4757_ (.A1(_0883_),
    .A2(_0890_),
    .B1(\i_tinyqv.cpu.instr_data_start[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1592_));
 sky130_fd_sc_hd__or2_1 _4758_ (.A(_0891_),
    .B(_1592_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1593_));
 sky130_fd_sc_hd__a2bb2o_1 _4759_ (.A1_N(_0612_),
    .A2_N(_1591_),
    .B1(_0748_),
    .B2(_1593_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1594_));
 sky130_fd_sc_hd__nor2_1 _4760_ (.A(\i_tinyqv.cpu.instr_data_start[11] ),
    .B(_0893_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1595_));
 sky130_fd_sc_hd__nor2_1 _4761_ (.A(_0894_),
    .B(_1595_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1596_));
 sky130_fd_sc_hd__nor2_1 _4762_ (.A(_0909_),
    .B(_1596_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1597_));
 sky130_fd_sc_hd__a2111o_1 _4763_ (.A1(_1589_),
    .A2(_1590_),
    .B1(_1594_),
    .C1(_1597_),
    .D1(_0688_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1598_));
 sky130_fd_sc_hd__xor2_1 _4764_ (.A(\i_tinyqv.cpu.instr_data_start[23] ),
    .B(_1333_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1599_));
 sky130_fd_sc_hd__a21oi_1 _4765_ (.A1(_0784_),
    .A2(_0898_),
    .B1(\i_tinyqv.cpu.instr_data_start[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1600_));
 sky130_fd_sc_hd__or2_1 _4766_ (.A(_0899_),
    .B(_1600_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1601_));
 sky130_fd_sc_hd__o2bb2a_1 _4767_ (.A1_N(_0610_),
    .A2_N(_1599_),
    .B1(_1601_),
    .B2(_0916_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1602_));
 sky130_fd_sc_hd__a21o_1 _4768_ (.A1(_1598_),
    .A2(_1602_),
    .B1(_0858_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1603_));
 sky130_fd_sc_hd__clkbuf_4 _4769_ (.A(_0841_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1604_));
 sky130_fd_sc_hd__nor2_1 _4770_ (.A(_1604_),
    .B(_0938_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1605_));
 sky130_fd_sc_hd__a221o_1 _4771_ (.A1(\i_tinyqv.cpu.i_core.mie[19] ),
    .A2(_0944_),
    .B1(net19),
    .B2(\i_tinyqv.cpu.i_core.mepc[3] ),
    .C1(_1605_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1606_));
 sky130_fd_sc_hd__mux2_1 _4772_ (.A0(\i_tinyqv.cpu.i_core.time_hi[2] ),
    .A1(\i_tinyqv.cpu.i_core.cycle_count_wide[6] ),
    .S(_1604_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1607_));
 sky130_fd_sc_hd__a22o_1 _4773_ (.A1(\i_tinyqv.cpu.i_core.cycle_count[3] ),
    .A2(_0931_),
    .B1(_1607_),
    .B2(_0927_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1608_));
 sky130_fd_sc_hd__nor2_1 _4774_ (.A(_0939_),
    .B(_1348_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1609_));
 sky130_fd_sc_hd__a22o_1 _4775_ (.A1(\i_tinyqv.cpu.i_core.mcause[3] ),
    .A2(_0947_),
    .B1(_1349_),
    .B2(\i_tinyqv.cpu.i_core.mstatus_mie ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1610_));
 sky130_fd_sc_hd__a221o_1 _4776_ (.A1(net15),
    .A2(_0991_),
    .B1(_1609_),
    .B2(\i_tinyqv.cpu.i_core.mstatus_mpie ),
    .C1(_1610_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1611_));
 sky130_fd_sc_hd__a2111o_1 _4777_ (.A1(\i_tinyqv.cpu.i_core.i_instrret.data[3] ),
    .A2(_0929_),
    .B1(_1606_),
    .C1(_1608_),
    .D1(_1611_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1612_));
 sky130_fd_sc_hd__a21oi_1 _4778_ (.A1(_0921_),
    .A2(_1612_),
    .B1(_0880_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1613_));
 sky130_fd_sc_hd__a22o_1 _4779_ (.A1(_0697_),
    .A2(_0880_),
    .B1(_1603_),
    .B2(_1613_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1614_));
 sky130_fd_sc_hd__mux2_1 _4780_ (.A0(\i_tinyqv.cpu.instr_data_in[15] ),
    .A1(\i_tinyqv.cpu.instr_data_in[7] ),
    .S(_1012_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1615_));
 sky130_fd_sc_hd__a22o_1 _4781_ (.A1(\i_spi.data[7] ),
    .A2(_1000_),
    .B1(_0986_),
    .B2(net9),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1616_));
 sky130_fd_sc_hd__a221o_1 _4782_ (.A1(\i_uart_rx.recieved_data[7] ),
    .A2(_0997_),
    .B1(net14),
    .B2(\gpio_out_sel[7] ),
    .C1(_1616_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1617_));
 sky130_fd_sc_hd__a211o_1 _4783_ (.A1(_1001_),
    .A2(uo_out[7]),
    .B1(_1617_),
    .C1(_0971_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1618_));
 sky130_fd_sc_hd__buf_2 _4784_ (.A(_0748_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1619_));
 sky130_fd_sc_hd__o211a_1 _4785_ (.A1(_0957_),
    .A2(_1615_),
    .B1(_1618_),
    .C1(_1619_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1620_));
 sky130_fd_sc_hd__mux2_1 _4786_ (.A0(\i_tinyqv.cpu.instr_data_in[15] ),
    .A1(\i_tinyqv.mem.qspi_data_buf[15] ),
    .S(_1017_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1621_));
 sky130_fd_sc_hd__mux2_1 _4787_ (.A0(\i_tinyqv.cpu.instr_data_in[11] ),
    .A1(\i_tinyqv.mem.qspi_data_buf[11] ),
    .S(_1017_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1622_));
 sky130_fd_sc_hd__mux2_1 _4788_ (.A0(_1621_),
    .A1(_1622_),
    .S(_0908_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1623_));
 sky130_fd_sc_hd__o211a_1 _4789_ (.A1(_0957_),
    .A2(_1623_),
    .B1(_0971_),
    .C1(_0907_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1624_));
 sky130_fd_sc_hd__a31o_1 _4790_ (.A1(\i_tinyqv.cpu.instr_data_in[11] ),
    .A2(_0869_),
    .A3(_0979_),
    .B1(_0865_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1625_));
 sky130_fd_sc_hd__a21o_1 _4791_ (.A1(\i_tinyqv.cpu.instr_data_in[3] ),
    .A2(_1012_),
    .B1(_1625_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1626_));
 sky130_fd_sc_hd__a22o_1 _4792_ (.A1(\gpio_out_sel[3] ),
    .A2(net14),
    .B1(uo_out[3]),
    .B2(_1001_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1627_));
 sky130_fd_sc_hd__a221o_1 _4793_ (.A1(\i_spi.data[3] ),
    .A2(_1000_),
    .B1(_0986_),
    .B2(net5),
    .C1(_1627_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1628_));
 sky130_fd_sc_hd__a211o_1 _4794_ (.A1(\i_uart_rx.recieved_data[3] ),
    .A2(_0997_),
    .B1(_1628_),
    .C1(_0971_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1629_));
 sky130_fd_sc_hd__a31o_1 _4795_ (.A1(_0689_),
    .A2(_1626_),
    .A3(_1629_),
    .B1(_0956_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1630_));
 sky130_fd_sc_hd__mux4_1 _4796_ (.A0(\i_tinyqv.mem.qspi_data_buf[27] ),
    .A1(\i_tinyqv.mem.qspi_data_buf[31] ),
    .A2(\i_tinyqv.cpu.instr_data_in[11] ),
    .A3(\i_tinyqv.cpu.instr_data_in[15] ),
    .S0(_0974_),
    .S1(_0979_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1631_));
 sky130_fd_sc_hd__a221o_1 _4797_ (.A1(\i_tinyqv.mem.data_from_read[19] ),
    .A2(_0689_),
    .B1(_0748_),
    .B2(\i_tinyqv.mem.data_from_read[23] ),
    .C1(_0865_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1632_));
 sky130_fd_sc_hd__o211a_1 _4798_ (.A1(_0970_),
    .A2(_0969_),
    .B1(_1632_),
    .C1(_0968_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1633_));
 sky130_fd_sc_hd__a211o_1 _4799_ (.A1(_0973_),
    .A2(_1631_),
    .B1(_1633_),
    .C1(_0752_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1634_));
 sky130_fd_sc_hd__o31a_1 _4800_ (.A1(_1620_),
    .A2(_1624_),
    .A3(_1630_),
    .B1(_1634_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1635_));
 sky130_fd_sc_hd__a21oi_2 _4801_ (.A1(_0955_),
    .A2(_1635_),
    .B1(_1023_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1636_));
 sky130_fd_sc_hd__a211oi_2 _4802_ (.A1(_0878_),
    .A2(_1614_),
    .B1(_1636_),
    .C1(_1025_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1637_));
 sky130_fd_sc_hd__a31o_4 _4803_ (.A1(_1034_),
    .A2(_1586_),
    .A3(_1588_),
    .B1(_1637_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1638_));
 sky130_fd_sc_hd__buf_6 _4804_ (.A(_1638_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.debug_rd[3] ));
 sky130_fd_sc_hd__mux2_1 _4805_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[15][3] ),
    .A1(net32),
    .S(_1190_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1639_));
 sky130_fd_sc_hd__clkbuf_1 _4806_ (.A(_1639_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0053_));
 sky130_fd_sc_hd__inv_2 _4807_ (.A(\i_tinyqv.cpu.i_core.i_registers.rd[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1640_));
 sky130_fd_sc_hd__and2_1 _4808_ (.A(\i_tinyqv.cpu.i_core.i_registers.rd[1] ),
    .B(_1640_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1641_));
 sky130_fd_sc_hd__and2_2 _4809_ (.A(_1189_),
    .B(_1641_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1642_));
 sky130_fd_sc_hd__mux2_1 _4810_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[14][0] ),
    .A1(\i_tinyqv.cpu.debug_rd[0] ),
    .S(_1642_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1643_));
 sky130_fd_sc_hd__clkbuf_1 _4811_ (.A(_1643_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0046_));
 sky130_fd_sc_hd__mux2_1 _4812_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[14][1] ),
    .A1(\i_tinyqv.cpu.debug_rd[1] ),
    .S(_1642_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1644_));
 sky130_fd_sc_hd__clkbuf_1 _4813_ (.A(_1644_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0047_));
 sky130_fd_sc_hd__mux2_1 _4814_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[14][2] ),
    .A1(\i_tinyqv.cpu.debug_rd[2] ),
    .S(_1642_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1645_));
 sky130_fd_sc_hd__clkbuf_1 _4815_ (.A(_1645_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0048_));
 sky130_fd_sc_hd__mux2_1 _4816_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[14][3] ),
    .A1(net32),
    .S(_1642_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1646_));
 sky130_fd_sc_hd__clkbuf_1 _4817_ (.A(_1646_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0049_));
 sky130_fd_sc_hd__nor2_1 _4818_ (.A(\i_tinyqv.cpu.i_core.i_registers.rd[1] ),
    .B(_1640_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1647_));
 sky130_fd_sc_hd__and2_2 _4819_ (.A(_1189_),
    .B(_1647_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1648_));
 sky130_fd_sc_hd__mux2_1 _4820_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[13][0] ),
    .A1(\i_tinyqv.cpu.debug_rd[0] ),
    .S(_1648_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1649_));
 sky130_fd_sc_hd__clkbuf_1 _4821_ (.A(_1649_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0042_));
 sky130_fd_sc_hd__mux2_1 _4822_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[13][1] ),
    .A1(\i_tinyqv.cpu.debug_rd[1] ),
    .S(_1648_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1650_));
 sky130_fd_sc_hd__clkbuf_1 _4823_ (.A(_1650_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0043_));
 sky130_fd_sc_hd__mux2_1 _4824_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[13][2] ),
    .A1(\i_tinyqv.cpu.debug_rd[2] ),
    .S(_1648_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1651_));
 sky130_fd_sc_hd__clkbuf_1 _4825_ (.A(_1651_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0044_));
 sky130_fd_sc_hd__mux2_1 _4826_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[13][3] ),
    .A1(\i_tinyqv.cpu.debug_rd[3] ),
    .S(_1648_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1652_));
 sky130_fd_sc_hd__clkbuf_1 _4827_ (.A(_1652_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0045_));
 sky130_fd_sc_hd__and3b_2 _4828_ (.A_N(\i_tinyqv.cpu.i_core.i_registers.rd[1] ),
    .B(_1640_),
    .C(_1189_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1653_));
 sky130_fd_sc_hd__mux2_1 _4829_ (.A0(net215),
    .A1(\i_tinyqv.cpu.debug_rd[0] ),
    .S(_1653_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1654_));
 sky130_fd_sc_hd__clkbuf_1 _4830_ (.A(_1654_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0038_));
 sky130_fd_sc_hd__mux2_1 _4831_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[12][1] ),
    .A1(\i_tinyqv.cpu.debug_rd[1] ),
    .S(_1653_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1655_));
 sky130_fd_sc_hd__clkbuf_1 _4832_ (.A(_1655_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0039_));
 sky130_fd_sc_hd__mux2_1 _4833_ (.A0(net103),
    .A1(\i_tinyqv.cpu.debug_rd[2] ),
    .S(_1653_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1656_));
 sky130_fd_sc_hd__clkbuf_1 _4834_ (.A(_1656_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0040_));
 sky130_fd_sc_hd__mux2_1 _4835_ (.A0(net101),
    .A1(net32),
    .S(_1653_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1657_));
 sky130_fd_sc_hd__clkbuf_1 _4836_ (.A(_1657_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0041_));
 sky130_fd_sc_hd__and3b_1 _4837_ (.A_N(\i_tinyqv.cpu.i_core.i_registers.rd[2] ),
    .B(\i_tinyqv.cpu.i_core.i_registers.rd[3] ),
    .C(_1188_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1658_));
 sky130_fd_sc_hd__and3_2 _4838_ (.A(\i_tinyqv.cpu.i_core.i_registers.rd[1] ),
    .B(\i_tinyqv.cpu.i_core.i_registers.rd[0] ),
    .C(_1658_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1659_));
 sky130_fd_sc_hd__mux2_1 _4839_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[11][0] ),
    .A1(\i_tinyqv.cpu.debug_rd[0] ),
    .S(_1659_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1660_));
 sky130_fd_sc_hd__clkbuf_1 _4840_ (.A(_1660_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0034_));
 sky130_fd_sc_hd__mux2_1 _4841_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[11][1] ),
    .A1(\i_tinyqv.cpu.debug_rd[1] ),
    .S(_1659_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1661_));
 sky130_fd_sc_hd__clkbuf_1 _4842_ (.A(_1661_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0035_));
 sky130_fd_sc_hd__mux2_1 _4843_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[11][2] ),
    .A1(\i_tinyqv.cpu.debug_rd[2] ),
    .S(_1659_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1662_));
 sky130_fd_sc_hd__clkbuf_1 _4844_ (.A(_1662_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0036_));
 sky130_fd_sc_hd__mux2_1 _4845_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[11][3] ),
    .A1(\i_tinyqv.cpu.debug_rd[3] ),
    .S(_1659_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1663_));
 sky130_fd_sc_hd__clkbuf_1 _4846_ (.A(_1663_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0037_));
 sky130_fd_sc_hd__and2_2 _4847_ (.A(_1641_),
    .B(_1658_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1664_));
 sky130_fd_sc_hd__mux2_1 _4848_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[10][0] ),
    .A1(\i_tinyqv.cpu.debug_rd[0] ),
    .S(_1664_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1665_));
 sky130_fd_sc_hd__clkbuf_1 _4849_ (.A(_1665_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0030_));
 sky130_fd_sc_hd__mux2_1 _4850_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[10][1] ),
    .A1(\i_tinyqv.cpu.debug_rd[1] ),
    .S(_1664_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1666_));
 sky130_fd_sc_hd__clkbuf_1 _4851_ (.A(_1666_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0031_));
 sky130_fd_sc_hd__mux2_1 _4852_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[10][2] ),
    .A1(\i_tinyqv.cpu.debug_rd[2] ),
    .S(_1664_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1667_));
 sky130_fd_sc_hd__clkbuf_1 _4853_ (.A(_1667_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0032_));
 sky130_fd_sc_hd__mux2_1 _4854_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[10][3] ),
    .A1(\i_tinyqv.cpu.debug_rd[3] ),
    .S(_1664_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1668_));
 sky130_fd_sc_hd__clkbuf_1 _4855_ (.A(_1668_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0033_));
 sky130_fd_sc_hd__and2_2 _4856_ (.A(_1647_),
    .B(_1658_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1669_));
 sky130_fd_sc_hd__mux2_1 _4857_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[9][0] ),
    .A1(\i_tinyqv.cpu.debug_rd[0] ),
    .S(_1669_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1670_));
 sky130_fd_sc_hd__clkbuf_1 _4858_ (.A(_1670_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0078_));
 sky130_fd_sc_hd__mux2_1 _4859_ (.A0(net254),
    .A1(\i_tinyqv.cpu.debug_rd[1] ),
    .S(_1669_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1671_));
 sky130_fd_sc_hd__clkbuf_1 _4860_ (.A(_1671_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0079_));
 sky130_fd_sc_hd__mux2_1 _4861_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[9][2] ),
    .A1(\i_tinyqv.cpu.debug_rd[2] ),
    .S(_1669_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1672_));
 sky130_fd_sc_hd__clkbuf_1 _4862_ (.A(_1672_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0080_));
 sky130_fd_sc_hd__mux2_1 _4863_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[9][3] ),
    .A1(\i_tinyqv.cpu.debug_rd[3] ),
    .S(_1669_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1673_));
 sky130_fd_sc_hd__clkbuf_1 _4864_ (.A(_1673_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0081_));
 sky130_fd_sc_hd__and3b_2 _4865_ (.A_N(\i_tinyqv.cpu.i_core.i_registers.rd[1] ),
    .B(_1640_),
    .C(_1658_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1674_));
 sky130_fd_sc_hd__mux2_1 _4866_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[8][0] ),
    .A1(\i_tinyqv.cpu.debug_rd[0] ),
    .S(_1674_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1675_));
 sky130_fd_sc_hd__clkbuf_1 _4867_ (.A(_1675_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0074_));
 sky130_fd_sc_hd__mux2_1 _4868_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[8][1] ),
    .A1(\i_tinyqv.cpu.debug_rd[1] ),
    .S(_1674_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1676_));
 sky130_fd_sc_hd__clkbuf_1 _4869_ (.A(_1676_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0075_));
 sky130_fd_sc_hd__mux2_1 _4870_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[8][2] ),
    .A1(\i_tinyqv.cpu.debug_rd[2] ),
    .S(_1674_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1677_));
 sky130_fd_sc_hd__clkbuf_1 _4871_ (.A(_1677_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0076_));
 sky130_fd_sc_hd__mux2_1 _4872_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[8][3] ),
    .A1(net32),
    .S(_1674_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1678_));
 sky130_fd_sc_hd__clkbuf_1 _4873_ (.A(_1678_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0077_));
 sky130_fd_sc_hd__nand3_2 _4874_ (.A(\i_tinyqv.cpu.i_core.i_registers.rd[1] ),
    .B(\i_tinyqv.cpu.i_core.i_registers.rd[0] ),
    .C(\i_tinyqv.cpu.i_core.i_registers.rd[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1679_));
 sky130_fd_sc_hd__nor3b_2 _4875_ (.A(_1679_),
    .B(\i_tinyqv.cpu.i_core.i_registers.rd[3] ),
    .C_N(_1188_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1680_));
 sky130_fd_sc_hd__mux2_1 _4876_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[7][0] ),
    .A1(\i_tinyqv.cpu.debug_rd[0] ),
    .S(_1680_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1681_));
 sky130_fd_sc_hd__clkbuf_1 _4877_ (.A(_1681_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0070_));
 sky130_fd_sc_hd__mux2_1 _4878_ (.A0(net216),
    .A1(\i_tinyqv.cpu.debug_rd[1] ),
    .S(_1680_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1682_));
 sky130_fd_sc_hd__clkbuf_1 _4879_ (.A(_1682_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0071_));
 sky130_fd_sc_hd__mux2_1 _4880_ (.A0(net150),
    .A1(\i_tinyqv.cpu.debug_rd[2] ),
    .S(_1680_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1683_));
 sky130_fd_sc_hd__clkbuf_1 _4881_ (.A(_1683_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0072_));
 sky130_fd_sc_hd__mux2_1 _4882_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[7][3] ),
    .A1(\i_tinyqv.cpu.debug_rd[3] ),
    .S(_1680_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1684_));
 sky130_fd_sc_hd__clkbuf_1 _4883_ (.A(_1684_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0073_));
 sky130_fd_sc_hd__and4b_2 _4884_ (.A_N(\i_tinyqv.cpu.i_core.i_registers.rd[3] ),
    .B(_1188_),
    .C(_1641_),
    .D(\i_tinyqv.cpu.i_core.i_registers.rd[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1685_));
 sky130_fd_sc_hd__mux2_1 _4885_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[6][0] ),
    .A1(_1184_),
    .S(_1685_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1686_));
 sky130_fd_sc_hd__clkbuf_1 _4886_ (.A(_1686_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0066_));
 sky130_fd_sc_hd__mux2_1 _4887_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[6][1] ),
    .A1(_1303_),
    .S(_1685_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1687_));
 sky130_fd_sc_hd__clkbuf_1 _4888_ (.A(_1687_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0067_));
 sky130_fd_sc_hd__mux2_1 _4889_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[6][2] ),
    .A1(_1380_),
    .S(_1685_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1688_));
 sky130_fd_sc_hd__clkbuf_1 _4890_ (.A(_1688_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0068_));
 sky130_fd_sc_hd__mux2_1 _4891_ (.A0(net152),
    .A1(_1638_),
    .S(_1685_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1689_));
 sky130_fd_sc_hd__clkbuf_1 _4892_ (.A(_1689_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0069_));
 sky130_fd_sc_hd__and4b_2 _4893_ (.A_N(\i_tinyqv.cpu.i_core.i_registers.rd[3] ),
    .B(_1188_),
    .C(_1647_),
    .D(\i_tinyqv.cpu.i_core.i_registers.rd[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1690_));
 sky130_fd_sc_hd__mux2_1 _4894_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[5][0] ),
    .A1(_1184_),
    .S(_1690_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1691_));
 sky130_fd_sc_hd__clkbuf_1 _4895_ (.A(_1691_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0062_));
 sky130_fd_sc_hd__mux2_1 _4896_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[5][1] ),
    .A1(_1303_),
    .S(_1690_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1692_));
 sky130_fd_sc_hd__clkbuf_1 _4897_ (.A(_1692_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0063_));
 sky130_fd_sc_hd__mux2_1 _4898_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[5][2] ),
    .A1(_1380_),
    .S(_1690_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1693_));
 sky130_fd_sc_hd__clkbuf_1 _4899_ (.A(_1693_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0064_));
 sky130_fd_sc_hd__mux2_1 _4900_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[5][3] ),
    .A1(_1638_),
    .S(_1690_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1694_));
 sky130_fd_sc_hd__clkbuf_1 _4901_ (.A(_1694_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0065_));
 sky130_fd_sc_hd__nor2_1 _4902_ (.A(\i_tinyqv.cpu.i_core.i_registers.rd[2] ),
    .B(\i_tinyqv.cpu.i_core.i_registers.rd[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1695_));
 sky130_fd_sc_hd__and3_2 _4903_ (.A(_1188_),
    .B(_1641_),
    .C(_1695_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1696_));
 sky130_fd_sc_hd__mux2_1 _4904_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[2][0] ),
    .A1(_1184_),
    .S(_1696_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1697_));
 sky130_fd_sc_hd__clkbuf_1 _4905_ (.A(_1697_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0058_));
 sky130_fd_sc_hd__mux2_1 _4906_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[2][1] ),
    .A1(_1303_),
    .S(_1696_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1698_));
 sky130_fd_sc_hd__clkbuf_1 _4907_ (.A(_1698_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0059_));
 sky130_fd_sc_hd__mux2_1 _4908_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[2][2] ),
    .A1(_1380_),
    .S(_1696_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1699_));
 sky130_fd_sc_hd__clkbuf_1 _4909_ (.A(_1699_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0060_));
 sky130_fd_sc_hd__mux2_1 _4910_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[2][3] ),
    .A1(_1638_),
    .S(_1696_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1700_));
 sky130_fd_sc_hd__clkbuf_1 _4911_ (.A(_1700_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0061_));
 sky130_fd_sc_hd__and3_2 _4912_ (.A(_1188_),
    .B(_1647_),
    .C(_1695_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1701_));
 sky130_fd_sc_hd__mux2_1 _4913_ (.A0(net198),
    .A1(_1184_),
    .S(_1701_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1702_));
 sky130_fd_sc_hd__clkbuf_1 _4914_ (.A(_1702_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0054_));
 sky130_fd_sc_hd__mux2_1 _4915_ (.A0(net268),
    .A1(_1303_),
    .S(_1701_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1703_));
 sky130_fd_sc_hd__clkbuf_1 _4916_ (.A(_1703_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0055_));
 sky130_fd_sc_hd__mux2_1 _4917_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[1][2] ),
    .A1(_1380_),
    .S(_1701_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1704_));
 sky130_fd_sc_hd__clkbuf_1 _4918_ (.A(_1704_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0056_));
 sky130_fd_sc_hd__mux2_1 _4919_ (.A0(\i_tinyqv.cpu.i_core.i_registers.reg_access[1][3] ),
    .A1(_1638_),
    .S(_1701_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1705_));
 sky130_fd_sc_hd__clkbuf_1 _4920_ (.A(_1705_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0057_));
 sky130_fd_sc_hd__clkbuf_4 _4921_ (.A(\i_tinyqv.mem.q_ctrl.fsm_state[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1706_));
 sky130_fd_sc_hd__buf_2 _4922_ (.A(\i_tinyqv.mem.q_ctrl.fsm_state[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1707_));
 sky130_fd_sc_hd__or2b_2 _4923_ (.A(_1707_),
    .B_N(\i_tinyqv.mem.q_ctrl.fsm_state[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1708_));
 sky130_fd_sc_hd__nor2_4 _4924_ (.A(_1706_),
    .B(_1708_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1709_));
 sky130_fd_sc_hd__and3b_1 _4925_ (.A_N(\i_tinyqv.mem.q_ctrl.fsm_state[1] ),
    .B(\i_tinyqv.mem.q_ctrl.fsm_state[0] ),
    .C(\i_tinyqv.mem.q_ctrl.fsm_state[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1710_));
 sky130_fd_sc_hd__buf_2 _4926_ (.A(_1710_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1711_));
 sky130_fd_sc_hd__clkbuf_4 _4927_ (.A(\i_tinyqv.cpu.instr_data_in[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1712_));
 sky130_fd_sc_hd__clkbuf_4 _4928_ (.A(\i_tinyqv.mem.q_ctrl.is_writing ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1713_));
 sky130_fd_sc_hd__or2b_1 _4929_ (.A(\i_tinyqv.mem.q_ctrl.fsm_state[1] ),
    .B_N(_1707_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1714_));
 sky130_fd_sc_hd__or2_1 _4930_ (.A(_1706_),
    .B(_1714_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1715_));
 sky130_fd_sc_hd__nor3_1 _4931_ (.A(_1713_),
    .B(\i_tinyqv.mem.q_ctrl.nibbles_remaining[0] ),
    .C(_1715_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1716_));
 sky130_fd_sc_hd__a221o_4 _4932_ (.A1(\i_tinyqv.mem.q_ctrl.addr[20] ),
    .A2(_1709_),
    .B1(_1711_),
    .B2(_1712_),
    .C1(_1716_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uio_out[1]));
 sky130_fd_sc_hd__buf_2 _4933_ (.A(\i_tinyqv.cpu.instr_data_in[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1717_));
 sky130_fd_sc_hd__a2bb2o_1 _4934_ (.A1_N(\i_tinyqv.mem.q_ctrl.nibbles_remaining[0] ),
    .A2_N(_1715_),
    .B1(_1709_),
    .B2(\i_tinyqv.mem.q_ctrl.addr[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1718_));
 sky130_fd_sc_hd__o21a_1 _4935_ (.A1(_1706_),
    .A2(_1708_),
    .B1(_1714_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1719_));
 sky130_fd_sc_hd__a211o_4 _4936_ (.A1(_1717_),
    .A2(_1711_),
    .B1(_1718_),
    .C1(_1719_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uio_out[2]));
 sky130_fd_sc_hd__buf_2 _4937_ (.A(\i_tinyqv.cpu.instr_data_in[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1720_));
 sky130_fd_sc_hd__a22o_4 _4938_ (.A1(\i_tinyqv.mem.q_ctrl.addr[22] ),
    .A2(_1709_),
    .B1(_1711_),
    .B2(_1720_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uio_out[4]));
 sky130_fd_sc_hd__buf_2 _4939_ (.A(\i_tinyqv.cpu.instr_data_in[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1721_));
 sky130_fd_sc_hd__a221o_1 _4940_ (.A1(_1706_),
    .A2(_1721_),
    .B1(\i_tinyqv.mem.q_ctrl.addr[23] ),
    .B2(_1709_),
    .C1(_1719_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1722_));
 sky130_fd_sc_hd__or2_1 _4941_ (.A(_1716_),
    .B(_1722_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1723_));
 sky130_fd_sc_hd__clkbuf_4 _4942_ (.A(_1723_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uio_out[5]));
 sky130_fd_sc_hd__and2_1 _4943_ (.A(\i_tinyqv.mem.q_ctrl.spi_data_oe[0] ),
    .B(net1),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1724_));
 sky130_fd_sc_hd__clkbuf_4 _4944_ (.A(_1724_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uio_oe[5]));
 sky130_fd_sc_hd__clkbuf_4 _4945_ (.A(_1557_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1725_));
 sky130_fd_sc_hd__and2_1 _4946_ (.A(_1001_),
    .B(_1725_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1726_));
 sky130_fd_sc_hd__clkbuf_4 _4947_ (.A(_1726_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1727_));
 sky130_fd_sc_hd__buf_4 _4948_ (.A(\i_debug_uart_tx.resetn ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1728_));
 sky130_fd_sc_hd__clkbuf_4 _4949_ (.A(_1728_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1729_));
 sky130_fd_sc_hd__nand2_2 _4950_ (.A(_1001_),
    .B(_1725_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1730_));
 sky130_fd_sc_hd__and3_1 _4951_ (.A(_1729_),
    .B(\gpio_out[0] ),
    .C(_1730_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1731_));
 sky130_fd_sc_hd__a21o_1 _4952_ (.A1(net117),
    .A2(_1727_),
    .B1(_1731_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0000_));
 sky130_fd_sc_hd__and3_1 _4953_ (.A(_1729_),
    .B(\gpio_out[1] ),
    .C(_1730_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1732_));
 sky130_fd_sc_hd__a21o_1 _4954_ (.A1(net97),
    .A2(_1727_),
    .B1(_1732_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0001_));
 sky130_fd_sc_hd__and3_1 _4955_ (.A(_1729_),
    .B(\gpio_out[2] ),
    .C(_1730_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1733_));
 sky130_fd_sc_hd__a21o_1 _4956_ (.A1(net98),
    .A2(_1727_),
    .B1(_1733_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0002_));
 sky130_fd_sc_hd__and3_1 _4957_ (.A(_1729_),
    .B(\gpio_out[3] ),
    .C(_1730_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1734_));
 sky130_fd_sc_hd__a21o_1 _4958_ (.A1(net197),
    .A2(_1727_),
    .B1(_1734_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0003_));
 sky130_fd_sc_hd__and3_1 _4959_ (.A(_1729_),
    .B(\gpio_out[4] ),
    .C(_1730_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1735_));
 sky130_fd_sc_hd__a21o_1 _4960_ (.A1(net238),
    .A2(_1727_),
    .B1(_1735_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0004_));
 sky130_fd_sc_hd__and3_1 _4961_ (.A(_1729_),
    .B(\gpio_out[5] ),
    .C(_1730_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1736_));
 sky130_fd_sc_hd__a21o_1 _4962_ (.A1(\i_debug_uart_tx.uart_tx_data[5] ),
    .A2(_1727_),
    .B1(_1736_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0005_));
 sky130_fd_sc_hd__buf_2 _4963_ (.A(_1728_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1737_));
 sky130_fd_sc_hd__and3_1 _4964_ (.A(_1737_),
    .B(\gpio_out[6] ),
    .C(_1730_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1738_));
 sky130_fd_sc_hd__a21o_1 _4965_ (.A1(net234),
    .A2(_1727_),
    .B1(_1738_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0006_));
 sky130_fd_sc_hd__and3_1 _4966_ (.A(_1737_),
    .B(\gpio_out[7] ),
    .C(_1730_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1739_));
 sky130_fd_sc_hd__a21o_1 _4967_ (.A1(\i_debug_uart_tx.uart_tx_data[7] ),
    .A2(_1727_),
    .B1(_1739_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0007_));
 sky130_fd_sc_hd__and2_1 _4968_ (.A(net14),
    .B(_1725_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1740_));
 sky130_fd_sc_hd__buf_2 _4969_ (.A(_1740_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1741_));
 sky130_fd_sc_hd__nand2_2 _4970_ (.A(net14),
    .B(_1725_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1742_));
 sky130_fd_sc_hd__and3_1 _4971_ (.A(_1737_),
    .B(\gpio_out_sel[0] ),
    .C(_1742_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1743_));
 sky130_fd_sc_hd__a21o_1 _4972_ (.A1(net117),
    .A2(_1741_),
    .B1(_1743_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0008_));
 sky130_fd_sc_hd__and3_1 _4973_ (.A(_1737_),
    .B(\gpio_out_sel[1] ),
    .C(_1742_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1744_));
 sky130_fd_sc_hd__a21o_1 _4974_ (.A1(net97),
    .A2(_1741_),
    .B1(_1744_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0009_));
 sky130_fd_sc_hd__and3_1 _4975_ (.A(_1737_),
    .B(\gpio_out_sel[2] ),
    .C(_1742_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1745_));
 sky130_fd_sc_hd__a21o_1 _4976_ (.A1(net98),
    .A2(_1741_),
    .B1(_1745_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0010_));
 sky130_fd_sc_hd__and3_1 _4977_ (.A(_1737_),
    .B(\gpio_out_sel[3] ),
    .C(_1742_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1746_));
 sky130_fd_sc_hd__a21o_1 _4978_ (.A1(net197),
    .A2(_1741_),
    .B1(_1746_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0011_));
 sky130_fd_sc_hd__and3_1 _4979_ (.A(_1737_),
    .B(\gpio_out_sel[4] ),
    .C(_1742_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1747_));
 sky130_fd_sc_hd__a21o_1 _4980_ (.A1(net238),
    .A2(_1741_),
    .B1(_1747_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0012_));
 sky130_fd_sc_hd__and3_1 _4981_ (.A(_1737_),
    .B(\gpio_out_sel[5] ),
    .C(_1742_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1748_));
 sky130_fd_sc_hd__a21o_1 _4982_ (.A1(net237),
    .A2(_1741_),
    .B1(_1748_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0013_));
 sky130_fd_sc_hd__and3_1 _4983_ (.A(_1737_),
    .B(\gpio_out_sel[6] ),
    .C(_1742_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1749_));
 sky130_fd_sc_hd__a21o_1 _4984_ (.A1(net234),
    .A2(_1741_),
    .B1(_1749_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0014_));
 sky130_fd_sc_hd__mux2_1 _4985_ (.A0(_1544_),
    .A1(\gpio_out_sel[7] ),
    .S(_1728_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1750_));
 sky130_fd_sc_hd__mux2_1 _4986_ (.A0(\i_debug_uart_tx.uart_tx_data[7] ),
    .A1(_1750_),
    .S(_1742_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1751_));
 sky130_fd_sc_hd__clkbuf_1 _4987_ (.A(_1751_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0015_));
 sky130_fd_sc_hd__buf_4 _4988_ (.A(\i_tinyqv.cpu.i_core.i_cycles.rstn ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1752_));
 sky130_fd_sc_hd__buf_4 _4989_ (.A(_1752_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1753_));
 sky130_fd_sc_hd__inv_2 _4990_ (.A(\i_tinyqv.cpu.no_write_in_progress ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1754_));
 sky130_fd_sc_hd__or2_2 _4991_ (.A(\i_tinyqv.cpu.i_core.cycle[1] ),
    .B(\i_tinyqv.cpu.i_core.cycle[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1755_));
 sky130_fd_sc_hd__or4_1 _4992_ (.A(_1410_),
    .B(_1754_),
    .C(_1604_),
    .D(_1755_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1756_));
 sky130_fd_sc_hd__or2_1 _4993_ (.A(_0836_),
    .B(_1756_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1757_));
 sky130_fd_sc_hd__buf_4 _4994_ (.A(_1757_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1758_));
 sky130_fd_sc_hd__nand2_1 _4995_ (.A(\i_tinyqv.cpu.is_load ),
    .B(_1442_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1759_));
 sky130_fd_sc_hd__nor2_1 _4996_ (.A(_1758_),
    .B(_1759_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1760_));
 sky130_fd_sc_hd__nor2_2 _4997_ (.A(_0836_),
    .B(_1756_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1761_));
 sky130_fd_sc_hd__and2_1 _4998_ (.A(\i_tinyqv.cpu.is_store ),
    .B(_1761_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1762_));
 sky130_fd_sc_hd__or2_1 _4999_ (.A(_1762_),
    .B(_1760_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1763_));
 sky130_fd_sc_hd__mux2_1 _5000_ (.A0(\i_tinyqv.cpu.data_continue ),
    .A1(_1440_),
    .S(_1763_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1764_));
 sky130_fd_sc_hd__o21a_1 _5001_ (.A1(_1753_),
    .A2(_1760_),
    .B1(_1764_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0028_));
 sky130_fd_sc_hd__or2b_1 _5002_ (.A(_1315_),
    .B_N(_1575_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1765_));
 sky130_fd_sc_hd__nand2_1 _5003_ (.A(\i_tinyqv.cpu.i_core.multiplier.accum[3] ),
    .B(_1576_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1766_));
 sky130_fd_sc_hd__o211a_1 _5004_ (.A1(net76),
    .A2(_0797_),
    .B1(\i_tinyqv.cpu.i_core.cycle[0] ),
    .C1(\i_tinyqv.cpu.i_core.i_shift.a[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1767_));
 sky130_fd_sc_hd__o311a_1 _5005_ (.A1(_0636_),
    .A2(_0641_),
    .A3(net72),
    .B1(\i_tinyqv.cpu.i_core.i_shift.a[1] ),
    .C1(\i_tinyqv.cpu.i_core.cycle[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1768_));
 sky130_fd_sc_hd__xnor2_1 _5006_ (.A(_1767_),
    .B(_1768_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1769_));
 sky130_fd_sc_hd__and2_1 _5007_ (.A(\i_tinyqv.cpu.i_core.i_shift.a[4] ),
    .B(_1166_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1770_));
 sky130_fd_sc_hd__xnor2_1 _5008_ (.A(_1769_),
    .B(_1770_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1771_));
 sky130_fd_sc_hd__nand2_1 _5009_ (.A(_1571_),
    .B(_1572_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1772_));
 sky130_fd_sc_hd__o21ai_1 _5010_ (.A1(_1573_),
    .A2(_1574_),
    .B1(_1772_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1773_));
 sky130_fd_sc_hd__xor2_1 _5011_ (.A(_1771_),
    .B(_1773_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1774_));
 sky130_fd_sc_hd__xnor2_1 _5012_ (.A(\i_tinyqv.cpu.i_core.multiplier.accum[4] ),
    .B(_1774_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1775_));
 sky130_fd_sc_hd__a21o_1 _5013_ (.A1(_1765_),
    .A2(_1766_),
    .B1(_1775_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1776_));
 sky130_fd_sc_hd__nand3_1 _5014_ (.A(_1765_),
    .B(_1766_),
    .C(_1775_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1777_));
 sky130_fd_sc_hd__nand2_1 _5015_ (.A(_1776_),
    .B(_1777_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1778_));
 sky130_fd_sc_hd__nand2_1 _5016_ (.A(\i_tinyqv.cpu.i_core.i_shift.a[3] ),
    .B(_1250_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1779_));
 sky130_fd_sc_hd__xor2_2 _5017_ (.A(_1778_),
    .B(_1779_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1780_));
 sky130_fd_sc_hd__nand2_1 _5018_ (.A(_1570_),
    .B(_1577_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1781_));
 sky130_fd_sc_hd__o21ai_2 _5019_ (.A1(_1578_),
    .A2(_1579_),
    .B1(_1781_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1782_));
 sky130_fd_sc_hd__xor2_2 _5020_ (.A(_1780_),
    .B(_1782_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1783_));
 sky130_fd_sc_hd__and2_1 _5021_ (.A(_1580_),
    .B(_1582_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1784_));
 sky130_fd_sc_hd__a31o_1 _5022_ (.A1(_1320_),
    .A2(_1321_),
    .A3(_1583_),
    .B1(_1784_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1785_));
 sky130_fd_sc_hd__xor2_1 _5023_ (.A(_1783_),
    .B(_1785_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0016_));
 sky130_fd_sc_hd__and2_1 _5024_ (.A(_1780_),
    .B(_1782_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1786_));
 sky130_fd_sc_hd__a21o_1 _5025_ (.A1(_1783_),
    .A2(_1785_),
    .B1(_1786_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1787_));
 sky130_fd_sc_hd__or2_1 _5026_ (.A(_1778_),
    .B(_1779_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1788_));
 sky130_fd_sc_hd__o31a_2 _5027_ (.A1(_0636_),
    .A2(_0641_),
    .A3(net73),
    .B1(\i_tinyqv.cpu.i_core.cycle[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1789_));
 sky130_fd_sc_hd__a22oi_1 _5028_ (.A1(\i_tinyqv.cpu.i_core.i_shift.a[3] ),
    .A2(_1309_),
    .B1(_1789_),
    .B2(\i_tinyqv.cpu.i_core.i_shift.a[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1790_));
 sky130_fd_sc_hd__a31o_1 _5029_ (.A1(\i_tinyqv.cpu.i_core.i_shift.a[3] ),
    .A2(_1767_),
    .A3(_1789_),
    .B1(_1790_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1791_));
 sky130_fd_sc_hd__nand2_1 _5030_ (.A(\i_tinyqv.cpu.i_core.i_shift.a[5] ),
    .B(_1166_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1792_));
 sky130_fd_sc_hd__xor2_1 _5031_ (.A(_1791_),
    .B(_1792_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1793_));
 sky130_fd_sc_hd__and2b_1 _5032_ (.A_N(_1769_),
    .B(_1770_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1794_));
 sky130_fd_sc_hd__a21o_1 _5033_ (.A1(_1767_),
    .A2(_1768_),
    .B1(_1794_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1795_));
 sky130_fd_sc_hd__xor2_1 _5034_ (.A(_1793_),
    .B(_1795_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1796_));
 sky130_fd_sc_hd__xnor2_1 _5035_ (.A(\i_tinyqv.cpu.i_core.multiplier.accum[5] ),
    .B(_1796_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1797_));
 sky130_fd_sc_hd__and2_1 _5036_ (.A(_1771_),
    .B(_1773_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1798_));
 sky130_fd_sc_hd__a21o_1 _5037_ (.A1(\i_tinyqv.cpu.i_core.multiplier.accum[4] ),
    .A2(_1774_),
    .B1(_1798_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1799_));
 sky130_fd_sc_hd__xor2_1 _5038_ (.A(_1797_),
    .B(_1799_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1800_));
 sky130_fd_sc_hd__nand2_1 _5039_ (.A(\i_tinyqv.cpu.i_core.i_shift.a[4] ),
    .B(_1250_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1801_));
 sky130_fd_sc_hd__xnor2_1 _5040_ (.A(_1800_),
    .B(_1801_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1802_));
 sky130_fd_sc_hd__and3_1 _5041_ (.A(_1776_),
    .B(_1788_),
    .C(_1802_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1803_));
 sky130_fd_sc_hd__a21oi_1 _5042_ (.A1(_1776_),
    .A2(_1788_),
    .B1(_1802_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1804_));
 sky130_fd_sc_hd__or2_1 _5043_ (.A(_1803_),
    .B(_1804_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1805_));
 sky130_fd_sc_hd__xnor2_1 _5044_ (.A(_1787_),
    .B(_1805_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0019_));
 sky130_fd_sc_hd__nand2_1 _5045_ (.A(\i_tinyqv.cpu.i_core.i_shift.a[3] ),
    .B(_1789_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1806_));
 sky130_fd_sc_hd__nand2_1 _5046_ (.A(\i_tinyqv.cpu.i_core.i_shift.a[4] ),
    .B(_1309_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1807_));
 sky130_fd_sc_hd__or2_1 _5047_ (.A(_1806_),
    .B(_1807_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1808_));
 sky130_fd_sc_hd__nand2_1 _5048_ (.A(_1806_),
    .B(_1807_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1809_));
 sky130_fd_sc_hd__nand2_1 _5049_ (.A(_1808_),
    .B(_1809_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1810_));
 sky130_fd_sc_hd__nand2_1 _5050_ (.A(\i_tinyqv.cpu.i_core.i_shift.a[6] ),
    .B(_1166_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1811_));
 sky130_fd_sc_hd__xor2_1 _5051_ (.A(_1810_),
    .B(_1811_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1812_));
 sky130_fd_sc_hd__buf_2 _5052_ (.A(_1789_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1813_));
 sky130_fd_sc_hd__nor2_1 _5053_ (.A(_1791_),
    .B(_1792_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1814_));
 sky130_fd_sc_hd__a31o_1 _5054_ (.A1(\i_tinyqv.cpu.i_core.i_shift.a[3] ),
    .A2(_1767_),
    .A3(_1813_),
    .B1(_1814_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1815_));
 sky130_fd_sc_hd__xor2_1 _5055_ (.A(_1812_),
    .B(_1815_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1816_));
 sky130_fd_sc_hd__xnor2_1 _5056_ (.A(\i_tinyqv.cpu.i_core.multiplier.accum[6] ),
    .B(_1816_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1817_));
 sky130_fd_sc_hd__and2_1 _5057_ (.A(_1793_),
    .B(_1795_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1818_));
 sky130_fd_sc_hd__a21o_1 _5058_ (.A1(\i_tinyqv.cpu.i_core.multiplier.accum[5] ),
    .A2(_1796_),
    .B1(_1818_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1819_));
 sky130_fd_sc_hd__xor2_1 _5059_ (.A(_1817_),
    .B(_1819_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1820_));
 sky130_fd_sc_hd__nand2_1 _5060_ (.A(\i_tinyqv.cpu.i_core.i_shift.a[5] ),
    .B(_1250_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1821_));
 sky130_fd_sc_hd__xor2_1 _5061_ (.A(_1820_),
    .B(_1821_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1822_));
 sky130_fd_sc_hd__and2b_1 _5062_ (.A_N(_1797_),
    .B(_1799_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1823_));
 sky130_fd_sc_hd__o21ba_1 _5063_ (.A1(_1800_),
    .A2(_1801_),
    .B1_N(_1823_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1824_));
 sky130_fd_sc_hd__xnor2_1 _5064_ (.A(_1822_),
    .B(_1824_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1825_));
 sky130_fd_sc_hd__a211o_1 _5065_ (.A1(_1783_),
    .A2(_1785_),
    .B1(_1804_),
    .C1(_1786_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1826_));
 sky130_fd_sc_hd__and3b_1 _5066_ (.A_N(_1803_),
    .B(_1825_),
    .C(_1826_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1827_));
 sky130_fd_sc_hd__and2b_1 _5067_ (.A_N(_1803_),
    .B(_1826_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1828_));
 sky130_fd_sc_hd__nor2_1 _5068_ (.A(_1825_),
    .B(_1828_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1829_));
 sky130_fd_sc_hd__nor2_1 _5069_ (.A(_1827_),
    .B(_1829_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0020_));
 sky130_fd_sc_hd__and2b_1 _5070_ (.A_N(_1824_),
    .B(_1822_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1830_));
 sky130_fd_sc_hd__nand2_1 _5071_ (.A(\i_tinyqv.cpu.i_core.i_shift.a[5] ),
    .B(_1789_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1831_));
 sky130_fd_sc_hd__or2_1 _5072_ (.A(_1807_),
    .B(_1831_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1832_));
 sky130_fd_sc_hd__a22o_1 _5073_ (.A1(\i_tinyqv.cpu.i_core.i_shift.a[5] ),
    .A2(_1309_),
    .B1(_1789_),
    .B2(\i_tinyqv.cpu.i_core.i_shift.a[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1833_));
 sky130_fd_sc_hd__nand2_1 _5074_ (.A(_1832_),
    .B(_1833_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1834_));
 sky130_fd_sc_hd__nand2_1 _5075_ (.A(_1054_),
    .B(_1167_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1835_));
 sky130_fd_sc_hd__xor2_1 _5076_ (.A(_1834_),
    .B(_1835_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1836_));
 sky130_fd_sc_hd__o21ai_1 _5077_ (.A1(_1810_),
    .A2(_1811_),
    .B1(_1808_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1837_));
 sky130_fd_sc_hd__nand2_1 _5078_ (.A(_1836_),
    .B(_1837_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1838_));
 sky130_fd_sc_hd__or2_1 _5079_ (.A(_1836_),
    .B(_1837_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1839_));
 sky130_fd_sc_hd__and2_1 _5080_ (.A(_1838_),
    .B(_1839_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1840_));
 sky130_fd_sc_hd__xnor2_1 _5081_ (.A(\i_tinyqv.cpu.i_core.multiplier.accum[7] ),
    .B(_1840_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1841_));
 sky130_fd_sc_hd__and2_1 _5082_ (.A(_1812_),
    .B(_1815_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1842_));
 sky130_fd_sc_hd__a21o_1 _5083_ (.A1(\i_tinyqv.cpu.i_core.multiplier.accum[6] ),
    .A2(_1816_),
    .B1(_1842_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1843_));
 sky130_fd_sc_hd__xor2_1 _5084_ (.A(_1841_),
    .B(_1843_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1844_));
 sky130_fd_sc_hd__clkbuf_4 _5085_ (.A(_1250_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1845_));
 sky130_fd_sc_hd__nand2_1 _5086_ (.A(\i_tinyqv.cpu.i_core.i_shift.a[6] ),
    .B(_1845_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1846_));
 sky130_fd_sc_hd__xor2_1 _5087_ (.A(_1844_),
    .B(_1846_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1847_));
 sky130_fd_sc_hd__and2b_1 _5088_ (.A_N(_1817_),
    .B(_1819_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1848_));
 sky130_fd_sc_hd__o21ba_1 _5089_ (.A1(_1820_),
    .A2(_1821_),
    .B1_N(_1848_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1849_));
 sky130_fd_sc_hd__xnor2_1 _5090_ (.A(_1847_),
    .B(_1849_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1850_));
 sky130_fd_sc_hd__o21a_1 _5091_ (.A1(_1830_),
    .A2(_1827_),
    .B1(_1850_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1851_));
 sky130_fd_sc_hd__nor3_1 _5092_ (.A(_1830_),
    .B(_1827_),
    .C(_1850_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1852_));
 sky130_fd_sc_hd__nor2_1 _5093_ (.A(_1851_),
    .B(_1852_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0021_));
 sky130_fd_sc_hd__and2b_1 _5094_ (.A_N(_1849_),
    .B(_1847_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1853_));
 sky130_fd_sc_hd__inv_2 _5095_ (.A(\i_tinyqv.cpu.i_core.i_shift.a[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1854_));
 sky130_fd_sc_hd__nand2_1 _5096_ (.A(\i_tinyqv.cpu.i_core.i_shift.a[6] ),
    .B(_1309_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1855_));
 sky130_fd_sc_hd__xnor2_1 _5097_ (.A(_1831_),
    .B(_1855_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1856_));
 sky130_fd_sc_hd__or3_1 _5098_ (.A(_1854_),
    .B(_1313_),
    .C(_1856_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1857_));
 sky130_fd_sc_hd__o21ai_1 _5099_ (.A1(_1854_),
    .A2(_1313_),
    .B1(_1856_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1858_));
 sky130_fd_sc_hd__and2_1 _5100_ (.A(_1857_),
    .B(_1858_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1859_));
 sky130_fd_sc_hd__o21ai_1 _5101_ (.A1(_1834_),
    .A2(_1835_),
    .B1(_1832_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1860_));
 sky130_fd_sc_hd__xor2_1 _5102_ (.A(_1859_),
    .B(_1860_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1861_));
 sky130_fd_sc_hd__nand2_1 _5103_ (.A(\i_tinyqv.cpu.i_core.multiplier.accum[8] ),
    .B(_1861_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1862_));
 sky130_fd_sc_hd__or2_1 _5104_ (.A(\i_tinyqv.cpu.i_core.multiplier.accum[8] ),
    .B(_1861_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1863_));
 sky130_fd_sc_hd__nand2_1 _5105_ (.A(_1862_),
    .B(_1863_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1864_));
 sky130_fd_sc_hd__a21bo_1 _5106_ (.A1(\i_tinyqv.cpu.i_core.multiplier.accum[7] ),
    .A2(_1840_),
    .B1_N(_1838_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1865_));
 sky130_fd_sc_hd__xor2_1 _5107_ (.A(_1864_),
    .B(_1865_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1866_));
 sky130_fd_sc_hd__nand2_1 _5108_ (.A(_1054_),
    .B(_1845_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1867_));
 sky130_fd_sc_hd__xor2_1 _5109_ (.A(_1866_),
    .B(_1867_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1868_));
 sky130_fd_sc_hd__or2b_1 _5110_ (.A(_1841_),
    .B_N(_1843_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1869_));
 sky130_fd_sc_hd__o21ai_1 _5111_ (.A1(_1844_),
    .A2(_1846_),
    .B1(_1869_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1870_));
 sky130_fd_sc_hd__nand2_1 _5112_ (.A(_1868_),
    .B(_1870_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1871_));
 sky130_fd_sc_hd__or2_1 _5113_ (.A(_1868_),
    .B(_1870_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1872_));
 sky130_fd_sc_hd__and2_1 _5114_ (.A(_1871_),
    .B(_1872_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1873_));
 sky130_fd_sc_hd__o21ai_1 _5115_ (.A1(_1853_),
    .A2(_1851_),
    .B1(_1873_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1874_));
 sky130_fd_sc_hd__or3_1 _5116_ (.A(_1853_),
    .B(_1851_),
    .C(_1873_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1875_));
 sky130_fd_sc_hd__and2_1 _5117_ (.A(_1874_),
    .B(_1875_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1876_));
 sky130_fd_sc_hd__clkbuf_1 _5118_ (.A(_1876_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0022_));
 sky130_fd_sc_hd__nand2_1 _5119_ (.A(_1859_),
    .B(_1860_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1877_));
 sky130_fd_sc_hd__nand2_1 _5120_ (.A(\i_tinyqv.cpu.i_core.i_shift.a[7] ),
    .B(_1789_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1878_));
 sky130_fd_sc_hd__or2_1 _5121_ (.A(_1855_),
    .B(_1878_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1879_));
 sky130_fd_sc_hd__buf_2 _5122_ (.A(_1309_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1880_));
 sky130_fd_sc_hd__a22o_1 _5123_ (.A1(_1054_),
    .A2(_1880_),
    .B1(_1789_),
    .B2(\i_tinyqv.cpu.i_core.i_shift.a[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1881_));
 sky130_fd_sc_hd__nand2_1 _5124_ (.A(_1879_),
    .B(_1881_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1882_));
 sky130_fd_sc_hd__nand2_1 _5125_ (.A(\i_tinyqv.cpu.i_core.i_shift.a[9] ),
    .B(_1167_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1883_));
 sky130_fd_sc_hd__xor2_1 _5126_ (.A(_1882_),
    .B(_1883_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1884_));
 sky130_fd_sc_hd__o21ai_1 _5127_ (.A1(_1831_),
    .A2(_1855_),
    .B1(_1857_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1885_));
 sky130_fd_sc_hd__xor2_1 _5128_ (.A(_1884_),
    .B(_1885_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1886_));
 sky130_fd_sc_hd__nand2_1 _5129_ (.A(\i_tinyqv.cpu.i_core.multiplier.accum[9] ),
    .B(_1886_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1887_));
 sky130_fd_sc_hd__or2_1 _5130_ (.A(\i_tinyqv.cpu.i_core.multiplier.accum[9] ),
    .B(_1886_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1888_));
 sky130_fd_sc_hd__nand2_1 _5131_ (.A(_1887_),
    .B(_1888_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1889_));
 sky130_fd_sc_hd__a21o_1 _5132_ (.A1(_1877_),
    .A2(_1862_),
    .B1(_1889_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1890_));
 sky130_fd_sc_hd__nand3_1 _5133_ (.A(_1877_),
    .B(_1862_),
    .C(_1889_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1891_));
 sky130_fd_sc_hd__nand2_1 _5134_ (.A(_1890_),
    .B(_1891_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1892_));
 sky130_fd_sc_hd__nand2_1 _5135_ (.A(\i_tinyqv.cpu.i_core.i_shift.a[8] ),
    .B(_1845_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1893_));
 sky130_fd_sc_hd__xor2_1 _5136_ (.A(_1892_),
    .B(_1893_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1894_));
 sky130_fd_sc_hd__or2b_1 _5137_ (.A(_1864_),
    .B_N(_1865_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1895_));
 sky130_fd_sc_hd__o21ai_1 _5138_ (.A1(_1866_),
    .A2(_1867_),
    .B1(_1895_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1896_));
 sky130_fd_sc_hd__nand2_1 _5139_ (.A(_1894_),
    .B(_1896_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1897_));
 sky130_fd_sc_hd__or2_1 _5140_ (.A(_1894_),
    .B(_1896_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1898_));
 sky130_fd_sc_hd__and2_1 _5141_ (.A(_1897_),
    .B(_1898_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1899_));
 sky130_fd_sc_hd__nand2_1 _5142_ (.A(_1871_),
    .B(_1874_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1900_));
 sky130_fd_sc_hd__xor2_1 _5143_ (.A(_1899_),
    .B(_1900_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0023_));
 sky130_fd_sc_hd__nand2_1 _5144_ (.A(_1884_),
    .B(_1885_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1901_));
 sky130_fd_sc_hd__nand2_1 _5145_ (.A(\i_tinyqv.cpu.i_core.i_shift.a[8] ),
    .B(_1880_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1902_));
 sky130_fd_sc_hd__xnor2_1 _5146_ (.A(_1878_),
    .B(_1902_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1903_));
 sky130_fd_sc_hd__nand2_1 _5147_ (.A(\i_tinyqv.cpu.i_core.i_shift.a[10] ),
    .B(_1167_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1904_));
 sky130_fd_sc_hd__xor2_1 _5148_ (.A(_1903_),
    .B(_1904_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1905_));
 sky130_fd_sc_hd__o21ai_1 _5149_ (.A1(_1882_),
    .A2(_1883_),
    .B1(_1879_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1906_));
 sky130_fd_sc_hd__nand2_1 _5150_ (.A(_1905_),
    .B(_1906_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1907_));
 sky130_fd_sc_hd__or2_1 _5151_ (.A(_1905_),
    .B(_1906_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1908_));
 sky130_fd_sc_hd__and2_1 _5152_ (.A(_1907_),
    .B(_1908_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1909_));
 sky130_fd_sc_hd__nand2_1 _5153_ (.A(\i_tinyqv.cpu.i_core.multiplier.accum[10] ),
    .B(_1909_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1910_));
 sky130_fd_sc_hd__or2_1 _5154_ (.A(\i_tinyqv.cpu.i_core.multiplier.accum[10] ),
    .B(_1909_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1911_));
 sky130_fd_sc_hd__nand2_1 _5155_ (.A(_1910_),
    .B(_1911_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1912_));
 sky130_fd_sc_hd__a21o_1 _5156_ (.A1(_1901_),
    .A2(_1887_),
    .B1(_1912_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1913_));
 sky130_fd_sc_hd__nand3_1 _5157_ (.A(_1901_),
    .B(_1887_),
    .C(_1912_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1914_));
 sky130_fd_sc_hd__nand2_1 _5158_ (.A(_1913_),
    .B(_1914_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1915_));
 sky130_fd_sc_hd__nand2_1 _5159_ (.A(\i_tinyqv.cpu.i_core.i_shift.a[9] ),
    .B(_1845_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1916_));
 sky130_fd_sc_hd__xor2_1 _5160_ (.A(_1915_),
    .B(_1916_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1917_));
 sky130_fd_sc_hd__o21ai_1 _5161_ (.A1(_1892_),
    .A2(_1893_),
    .B1(_1890_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1918_));
 sky130_fd_sc_hd__nand2_1 _5162_ (.A(_1917_),
    .B(_1918_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1919_));
 sky130_fd_sc_hd__or2_1 _5163_ (.A(_1917_),
    .B(_1918_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1920_));
 sky130_fd_sc_hd__and2_1 _5164_ (.A(_1919_),
    .B(_1920_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1921_));
 sky130_fd_sc_hd__a21bo_1 _5165_ (.A1(_1871_),
    .A2(_1874_),
    .B1_N(_1899_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1922_));
 sky130_fd_sc_hd__nand2_1 _5166_ (.A(_1897_),
    .B(_1922_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1923_));
 sky130_fd_sc_hd__xor2_1 _5167_ (.A(_1921_),
    .B(_1923_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0024_));
 sky130_fd_sc_hd__nand2_1 _5168_ (.A(\i_tinyqv.cpu.i_core.i_shift.a[8] ),
    .B(_1813_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1924_));
 sky130_fd_sc_hd__nand2_1 _5169_ (.A(\i_tinyqv.cpu.i_core.i_shift.a[9] ),
    .B(_1880_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1925_));
 sky130_fd_sc_hd__xnor2_1 _5170_ (.A(_1924_),
    .B(_1925_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1926_));
 sky130_fd_sc_hd__nand2_1 _5171_ (.A(\i_tinyqv.cpu.i_core.i_shift.a[11] ),
    .B(_1167_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1927_));
 sky130_fd_sc_hd__xor2_1 _5172_ (.A(_1926_),
    .B(_1927_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1928_));
 sky130_fd_sc_hd__nand2_1 _5173_ (.A(_1054_),
    .B(_1880_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1929_));
 sky130_fd_sc_hd__or2_1 _5174_ (.A(_1929_),
    .B(_1924_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1930_));
 sky130_fd_sc_hd__o21ai_1 _5175_ (.A1(_1903_),
    .A2(_1904_),
    .B1(_1930_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1931_));
 sky130_fd_sc_hd__nand2_1 _5176_ (.A(_1928_),
    .B(_1931_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1932_));
 sky130_fd_sc_hd__or2_1 _5177_ (.A(_1928_),
    .B(_1931_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1933_));
 sky130_fd_sc_hd__and2_1 _5178_ (.A(_1932_),
    .B(_1933_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1934_));
 sky130_fd_sc_hd__nand2_1 _5179_ (.A(\i_tinyqv.cpu.i_core.multiplier.accum[11] ),
    .B(_1934_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1935_));
 sky130_fd_sc_hd__or2_1 _5180_ (.A(\i_tinyqv.cpu.i_core.multiplier.accum[11] ),
    .B(_1934_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1936_));
 sky130_fd_sc_hd__nand2_1 _5181_ (.A(_1935_),
    .B(_1936_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1937_));
 sky130_fd_sc_hd__a21o_1 _5182_ (.A1(_1907_),
    .A2(_1910_),
    .B1(_1937_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1938_));
 sky130_fd_sc_hd__nand3_1 _5183_ (.A(_1907_),
    .B(_1910_),
    .C(_1937_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1939_));
 sky130_fd_sc_hd__nand2_1 _5184_ (.A(_1938_),
    .B(_1939_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1940_));
 sky130_fd_sc_hd__nand2_1 _5185_ (.A(\i_tinyqv.cpu.i_core.i_shift.a[10] ),
    .B(_1845_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1941_));
 sky130_fd_sc_hd__xor2_1 _5186_ (.A(_1940_),
    .B(_1941_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1942_));
 sky130_fd_sc_hd__o21ai_1 _5187_ (.A1(_1915_),
    .A2(_1916_),
    .B1(_1913_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1943_));
 sky130_fd_sc_hd__and2_1 _5188_ (.A(_1942_),
    .B(_1943_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1944_));
 sky130_fd_sc_hd__inv_2 _5189_ (.A(_1944_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1945_));
 sky130_fd_sc_hd__or2_1 _5190_ (.A(_1942_),
    .B(_1943_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1946_));
 sky130_fd_sc_hd__and2_1 _5191_ (.A(_1945_),
    .B(_1946_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1947_));
 sky130_fd_sc_hd__a21bo_1 _5192_ (.A1(_1897_),
    .A2(_1922_),
    .B1_N(_1921_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1948_));
 sky130_fd_sc_hd__nand2_1 _5193_ (.A(_1919_),
    .B(_1948_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1949_));
 sky130_fd_sc_hd__xor2_1 _5194_ (.A(_1947_),
    .B(_1949_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0025_));
 sky130_fd_sc_hd__nand2_1 _5195_ (.A(\i_tinyqv.cpu.i_core.i_shift.a[9] ),
    .B(_1813_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1950_));
 sky130_fd_sc_hd__nand2_1 _5196_ (.A(\i_tinyqv.cpu.i_core.i_shift.a[10] ),
    .B(_1880_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1951_));
 sky130_fd_sc_hd__xnor2_1 _5197_ (.A(_1950_),
    .B(_1951_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1952_));
 sky130_fd_sc_hd__nand2_1 _5198_ (.A(\i_tinyqv.cpu.i_core.i_shift.a[12] ),
    .B(_1167_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1953_));
 sky130_fd_sc_hd__xor2_1 _5199_ (.A(_1952_),
    .B(_1953_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1954_));
 sky130_fd_sc_hd__or2_1 _5200_ (.A(_1902_),
    .B(_1950_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1955_));
 sky130_fd_sc_hd__o21ai_1 _5201_ (.A1(_1926_),
    .A2(_1927_),
    .B1(_1955_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1956_));
 sky130_fd_sc_hd__nand2_1 _5202_ (.A(_1954_),
    .B(_1956_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1957_));
 sky130_fd_sc_hd__or2_1 _5203_ (.A(_1954_),
    .B(_1956_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1958_));
 sky130_fd_sc_hd__and2_1 _5204_ (.A(_1957_),
    .B(_1958_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1959_));
 sky130_fd_sc_hd__nand2_1 _5205_ (.A(\i_tinyqv.cpu.i_core.multiplier.accum[12] ),
    .B(_1959_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1960_));
 sky130_fd_sc_hd__or2_1 _5206_ (.A(\i_tinyqv.cpu.i_core.multiplier.accum[12] ),
    .B(_1959_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1961_));
 sky130_fd_sc_hd__nand2_1 _5207_ (.A(_1960_),
    .B(_1961_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1962_));
 sky130_fd_sc_hd__a21o_1 _5208_ (.A1(_1932_),
    .A2(_1935_),
    .B1(_1962_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1963_));
 sky130_fd_sc_hd__nand3_1 _5209_ (.A(_1932_),
    .B(_1935_),
    .C(_1962_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1964_));
 sky130_fd_sc_hd__nand2_1 _5210_ (.A(_1963_),
    .B(_1964_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1965_));
 sky130_fd_sc_hd__nand2_1 _5211_ (.A(\i_tinyqv.cpu.i_core.i_shift.a[11] ),
    .B(_1845_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1966_));
 sky130_fd_sc_hd__xor2_1 _5212_ (.A(_1965_),
    .B(_1966_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1967_));
 sky130_fd_sc_hd__o21ai_1 _5213_ (.A1(_1940_),
    .A2(_1941_),
    .B1(_1938_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1968_));
 sky130_fd_sc_hd__nand2_1 _5214_ (.A(_1967_),
    .B(_1968_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1969_));
 sky130_fd_sc_hd__or2_1 _5215_ (.A(_1967_),
    .B(_1968_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1970_));
 sky130_fd_sc_hd__and2_1 _5216_ (.A(_1969_),
    .B(_1970_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1971_));
 sky130_fd_sc_hd__a21bo_1 _5217_ (.A1(_1919_),
    .A2(_1948_),
    .B1_N(_1947_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1972_));
 sky130_fd_sc_hd__nand2_1 _5218_ (.A(_1945_),
    .B(_1972_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1973_));
 sky130_fd_sc_hd__xor2_1 _5219_ (.A(_1971_),
    .B(_1973_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0026_));
 sky130_fd_sc_hd__nand2_1 _5220_ (.A(\i_tinyqv.cpu.i_core.i_shift.a[10] ),
    .B(_1813_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1974_));
 sky130_fd_sc_hd__nand2_1 _5221_ (.A(\i_tinyqv.cpu.i_core.i_shift.a[11] ),
    .B(_1880_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1975_));
 sky130_fd_sc_hd__xnor2_1 _5222_ (.A(_1974_),
    .B(_1975_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1976_));
 sky130_fd_sc_hd__nand2_1 _5223_ (.A(\i_tinyqv.cpu.i_core.i_shift.a[13] ),
    .B(_1167_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1977_));
 sky130_fd_sc_hd__xor2_1 _5224_ (.A(_1976_),
    .B(_1977_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1978_));
 sky130_fd_sc_hd__or2_1 _5225_ (.A(_1925_),
    .B(_1974_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1979_));
 sky130_fd_sc_hd__o21ai_1 _5226_ (.A1(_1952_),
    .A2(_1953_),
    .B1(_1979_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1980_));
 sky130_fd_sc_hd__nand2_1 _5227_ (.A(_1978_),
    .B(_1980_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1981_));
 sky130_fd_sc_hd__or2_1 _5228_ (.A(_1978_),
    .B(_1980_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1982_));
 sky130_fd_sc_hd__and2_1 _5229_ (.A(_1981_),
    .B(_1982_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1983_));
 sky130_fd_sc_hd__nand2_1 _5230_ (.A(\i_tinyqv.cpu.i_core.multiplier.accum[13] ),
    .B(_1983_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1984_));
 sky130_fd_sc_hd__or2_1 _5231_ (.A(\i_tinyqv.cpu.i_core.multiplier.accum[13] ),
    .B(_1983_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1985_));
 sky130_fd_sc_hd__nand2_1 _5232_ (.A(_1984_),
    .B(_1985_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1986_));
 sky130_fd_sc_hd__a21o_1 _5233_ (.A1(_1957_),
    .A2(_1960_),
    .B1(_1986_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1987_));
 sky130_fd_sc_hd__nand3_1 _5234_ (.A(_1957_),
    .B(_1960_),
    .C(_1986_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1988_));
 sky130_fd_sc_hd__nand2_1 _5235_ (.A(_1987_),
    .B(_1988_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1989_));
 sky130_fd_sc_hd__nand2_1 _5236_ (.A(\i_tinyqv.cpu.i_core.i_shift.a[12] ),
    .B(_1845_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1990_));
 sky130_fd_sc_hd__xor2_1 _5237_ (.A(_1989_),
    .B(_1990_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1991_));
 sky130_fd_sc_hd__o21ai_1 _5238_ (.A1(_1965_),
    .A2(_1966_),
    .B1(_1963_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1992_));
 sky130_fd_sc_hd__nand2_1 _5239_ (.A(_1991_),
    .B(_1992_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1993_));
 sky130_fd_sc_hd__or2_1 _5240_ (.A(_1991_),
    .B(_1992_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1994_));
 sky130_fd_sc_hd__and2_1 _5241_ (.A(_1993_),
    .B(_1994_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1995_));
 sky130_fd_sc_hd__a21bo_1 _5242_ (.A1(_1945_),
    .A2(_1972_),
    .B1_N(_1971_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1996_));
 sky130_fd_sc_hd__nand2_1 _5243_ (.A(_1969_),
    .B(_1996_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1997_));
 sky130_fd_sc_hd__xor2_1 _5244_ (.A(_1995_),
    .B(_1997_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0027_));
 sky130_fd_sc_hd__nand2_1 _5245_ (.A(\i_tinyqv.cpu.i_core.i_shift.a[11] ),
    .B(_1813_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1998_));
 sky130_fd_sc_hd__nand2_1 _5246_ (.A(\i_tinyqv.cpu.i_core.i_shift.a[12] ),
    .B(_1880_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1999_));
 sky130_fd_sc_hd__xnor2_1 _5247_ (.A(_1998_),
    .B(_1999_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2000_));
 sky130_fd_sc_hd__nand2_1 _5248_ (.A(\i_tinyqv.cpu.i_core.i_shift.a[14] ),
    .B(_1167_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2001_));
 sky130_fd_sc_hd__xor2_1 _5249_ (.A(_2000_),
    .B(_2001_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2002_));
 sky130_fd_sc_hd__or2_1 _5250_ (.A(_1951_),
    .B(_1998_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2003_));
 sky130_fd_sc_hd__o21ai_1 _5251_ (.A1(_1976_),
    .A2(_1977_),
    .B1(_2003_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2004_));
 sky130_fd_sc_hd__nand2_1 _5252_ (.A(_2002_),
    .B(_2004_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2005_));
 sky130_fd_sc_hd__or2_1 _5253_ (.A(_2002_),
    .B(_2004_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2006_));
 sky130_fd_sc_hd__and2_1 _5254_ (.A(_2005_),
    .B(_2006_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2007_));
 sky130_fd_sc_hd__nand2_1 _5255_ (.A(\i_tinyqv.cpu.i_core.multiplier.accum[14] ),
    .B(_2007_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2008_));
 sky130_fd_sc_hd__or2_1 _5256_ (.A(\i_tinyqv.cpu.i_core.multiplier.accum[14] ),
    .B(_2007_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2009_));
 sky130_fd_sc_hd__nand2_1 _5257_ (.A(_2008_),
    .B(_2009_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2010_));
 sky130_fd_sc_hd__a21o_1 _5258_ (.A1(_1981_),
    .A2(_1984_),
    .B1(_2010_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2011_));
 sky130_fd_sc_hd__nand3_1 _5259_ (.A(_1981_),
    .B(_1984_),
    .C(_2010_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2012_));
 sky130_fd_sc_hd__nand2_1 _5260_ (.A(_2011_),
    .B(_2012_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2013_));
 sky130_fd_sc_hd__nand2_1 _5261_ (.A(\i_tinyqv.cpu.i_core.i_shift.a[13] ),
    .B(_1845_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2014_));
 sky130_fd_sc_hd__xor2_1 _5262_ (.A(_2013_),
    .B(_2014_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2015_));
 sky130_fd_sc_hd__o21ai_1 _5263_ (.A1(_1989_),
    .A2(_1990_),
    .B1(_1987_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2016_));
 sky130_fd_sc_hd__nand2_1 _5264_ (.A(_2015_),
    .B(_2016_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2017_));
 sky130_fd_sc_hd__or2_1 _5265_ (.A(_2015_),
    .B(_2016_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2018_));
 sky130_fd_sc_hd__and2_1 _5266_ (.A(_2017_),
    .B(_2018_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2019_));
 sky130_fd_sc_hd__a21bo_1 _5267_ (.A1(_1969_),
    .A2(_1996_),
    .B1_N(_1995_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2020_));
 sky130_fd_sc_hd__nand2_1 _5268_ (.A(_1993_),
    .B(_2020_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2021_));
 sky130_fd_sc_hd__xor2_1 _5269_ (.A(_2019_),
    .B(_2021_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0017_));
 sky130_fd_sc_hd__inv_2 _5270_ (.A(\i_tinyqv.cpu.i_core.i_shift.a[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2022_));
 sky130_fd_sc_hd__nand2_1 _5271_ (.A(\i_tinyqv.cpu.i_core.i_shift.a[12] ),
    .B(_1813_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2023_));
 sky130_fd_sc_hd__nand2_1 _5272_ (.A(\i_tinyqv.cpu.i_core.i_shift.a[13] ),
    .B(_1880_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2024_));
 sky130_fd_sc_hd__xnor2_1 _5273_ (.A(_2023_),
    .B(_2024_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2025_));
 sky130_fd_sc_hd__or3_1 _5274_ (.A(_2022_),
    .B(_1313_),
    .C(_2025_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2026_));
 sky130_fd_sc_hd__o21ai_1 _5275_ (.A1(_2022_),
    .A2(_1313_),
    .B1(_2025_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2027_));
 sky130_fd_sc_hd__and2_1 _5276_ (.A(_2026_),
    .B(_2027_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2028_));
 sky130_fd_sc_hd__or2_1 _5277_ (.A(_1975_),
    .B(_2023_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2029_));
 sky130_fd_sc_hd__o21ai_1 _5278_ (.A1(_2000_),
    .A2(_2001_),
    .B1(_2029_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2030_));
 sky130_fd_sc_hd__xor2_1 _5279_ (.A(_2028_),
    .B(_2030_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2031_));
 sky130_fd_sc_hd__nor2_1 _5280_ (.A(\i_tinyqv.cpu.i_core.multiplier.accum[15] ),
    .B(_2031_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2032_));
 sky130_fd_sc_hd__and2_1 _5281_ (.A(\i_tinyqv.cpu.i_core.multiplier.accum[15] ),
    .B(_2031_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2033_));
 sky130_fd_sc_hd__or2_1 _5282_ (.A(_2032_),
    .B(_2033_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2034_));
 sky130_fd_sc_hd__nand3_1 _5283_ (.A(_2005_),
    .B(_2008_),
    .C(_2034_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2035_));
 sky130_fd_sc_hd__a21o_1 _5284_ (.A1(_2005_),
    .A2(_2008_),
    .B1(_2034_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2036_));
 sky130_fd_sc_hd__nand2_1 _5285_ (.A(_2035_),
    .B(_2036_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2037_));
 sky130_fd_sc_hd__nand2_1 _5286_ (.A(\i_tinyqv.cpu.i_core.i_shift.a[14] ),
    .B(_1845_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2038_));
 sky130_fd_sc_hd__xor2_1 _5287_ (.A(_2037_),
    .B(_2038_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2039_));
 sky130_fd_sc_hd__o21ai_1 _5288_ (.A1(_2013_),
    .A2(_2014_),
    .B1(_2011_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2040_));
 sky130_fd_sc_hd__nand2_1 _5289_ (.A(_2039_),
    .B(_2040_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2041_));
 sky130_fd_sc_hd__or2_1 _5290_ (.A(_2039_),
    .B(_2040_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2042_));
 sky130_fd_sc_hd__and2_1 _5291_ (.A(_2041_),
    .B(_2042_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2043_));
 sky130_fd_sc_hd__a21bo_1 _5292_ (.A1(_1993_),
    .A2(_2020_),
    .B1_N(_2019_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2044_));
 sky130_fd_sc_hd__nand2_1 _5293_ (.A(_2017_),
    .B(_2044_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2045_));
 sky130_fd_sc_hd__xor2_1 _5294_ (.A(_2043_),
    .B(_2045_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0018_));
 sky130_fd_sc_hd__and2_1 _5295_ (.A(_0701_),
    .B(_0821_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2046_));
 sky130_fd_sc_hd__clkbuf_1 _5296_ (.A(_2046_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.cy_out ));
 sky130_fd_sc_hd__and3_1 _5297_ (.A(\i_tinyqv.cpu.data_ready_core ),
    .B(\i_tinyqv.cpu.i_core.cycle[1] ),
    .C(_0744_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2047_));
 sky130_fd_sc_hd__a21o_1 _5298_ (.A1(net138),
    .A2(_1026_),
    .B1(_2047_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0084_));
 sky130_fd_sc_hd__and4_1 _5299_ (.A(_1752_),
    .B(_1387_),
    .C(_0861_),
    .D(_1031_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2048_));
 sky130_fd_sc_hd__a31o_1 _5300_ (.A1(_1753_),
    .A2(\i_tinyqv.cpu.i_core.cycle[0] ),
    .A3(_1604_),
    .B1(_2048_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0085_));
 sky130_fd_sc_hd__clkbuf_4 _5301_ (.A(_1752_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2049_));
 sky130_fd_sc_hd__o2111a_1 _5302_ (.A1(\i_tinyqv.cpu.i_core.cycle[1] ),
    .A2(_1387_),
    .B1(_0862_),
    .C1(_1755_),
    .D1(_2049_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0086_));
 sky130_fd_sc_hd__nand2_1 _5303_ (.A(\i_tinyqv.cpu.i_core.mie[16] ),
    .B(\i_tinyqv.cpu.i_core.mip[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2050_));
 sky130_fd_sc_hd__and3_1 _5304_ (.A(\i_tinyqv.cpu.i_core.mie[19] ),
    .B(_0991_),
    .C(_1402_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2051_));
 sky130_fd_sc_hd__a31o_1 _5305_ (.A1(\i_tinyqv.cpu.i_core.mie[17] ),
    .A2(\i_tinyqv.cpu.i_core.mip[17] ),
    .A3(_2050_),
    .B1(_2051_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2052_));
 sky130_fd_sc_hd__and3_1 _5306_ (.A(\i_tinyqv.cpu.i_core.is_interrupt ),
    .B(_0744_),
    .C(_2052_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2053_));
 sky130_fd_sc_hd__or4_2 _5307_ (.A(_1026_),
    .B(_0855_),
    .C(_1173_),
    .D(_0924_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2054_));
 sky130_fd_sc_hd__or2_1 _5308_ (.A(\i_tinyqv.cpu.i_core.is_interrupt ),
    .B(_2054_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2055_));
 sky130_fd_sc_hd__a21o_2 _5309_ (.A1(_1394_),
    .A2(_1392_),
    .B1(\i_tinyqv.cpu.i_core.is_interrupt ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2056_));
 sky130_fd_sc_hd__nand2_2 _5310_ (.A(_0744_),
    .B(_2056_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2057_));
 sky130_fd_sc_hd__a2bb2o_1 _5311_ (.A1_N(_0922_),
    .A2_N(_2055_),
    .B1(_2057_),
    .B2(\i_tinyqv.cpu.i_core.mcause[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2058_));
 sky130_fd_sc_hd__nor2_1 _5312_ (.A(_0777_),
    .B(_2055_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2059_));
 sky130_fd_sc_hd__and4_1 _5313_ (.A(_0697_),
    .B(_0814_),
    .C(_0707_),
    .D(_2059_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2060_));
 sky130_fd_sc_hd__clkbuf_4 _5314_ (.A(_1752_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2061_));
 sky130_fd_sc_hd__o31a_1 _5315_ (.A1(_2053_),
    .A2(_2058_),
    .A3(_2060_),
    .B1(_2061_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0087_));
 sky130_fd_sc_hd__inv_2 _5316_ (.A(_2057_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2062_));
 sky130_fd_sc_hd__nand2_1 _5317_ (.A(\i_tinyqv.cpu.i_core.mie[18] ),
    .B(_1228_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2063_));
 sky130_fd_sc_hd__nand2_1 _5318_ (.A(\i_tinyqv.cpu.i_core.is_interrupt ),
    .B(_0744_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2064_));
 sky130_fd_sc_hd__o21bai_1 _5319_ (.A1(_1401_),
    .A2(_2063_),
    .B1_N(_2064_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2065_));
 sky130_fd_sc_hd__o221a_1 _5320_ (.A1(net159),
    .A2(_2062_),
    .B1(_2065_),
    .B2(_2051_),
    .C1(_1753_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0088_));
 sky130_fd_sc_hd__buf_4 _5321_ (.A(_1400_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2066_));
 sky130_fd_sc_hd__clkbuf_4 _5322_ (.A(_2066_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2067_));
 sky130_fd_sc_hd__a21oi_1 _5323_ (.A1(net123),
    .A2(_2057_),
    .B1(_2060_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2068_));
 sky130_fd_sc_hd__nor2_1 _5324_ (.A(_2067_),
    .B(_2068_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0089_));
 sky130_fd_sc_hd__nand2_1 _5325_ (.A(net158),
    .B(_2054_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2069_));
 sky130_fd_sc_hd__a21oi_1 _5326_ (.A1(_2064_),
    .A2(_2069_),
    .B1(_2067_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0090_));
 sky130_fd_sc_hd__nor2_1 _5327_ (.A(\i_tinyqv.cpu.i_core.mstatus_mte ),
    .B(_2054_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2070_));
 sky130_fd_sc_hd__a21o_1 _5328_ (.A1(net99),
    .A2(_1026_),
    .B1(_2070_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0091_));
 sky130_fd_sc_hd__o21a_1 _5329_ (.A1(\i_tinyqv.cpu.i_core.i_cycles.cy ),
    .A2(_0744_),
    .B1(\i_tinyqv.cpu.i_core.cycle_count[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2071_));
 sky130_fd_sc_hd__and3_1 _5330_ (.A(\i_tinyqv.cpu.i_core.cycle_count[2] ),
    .B(\i_tinyqv.cpu.i_core.cycle_count[1] ),
    .C(_2071_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2072_));
 sky130_fd_sc_hd__nand2_1 _5331_ (.A(net235),
    .B(_2072_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2073_));
 sky130_fd_sc_hd__nor2_1 _5332_ (.A(_1604_),
    .B(_2073_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2074_));
 sky130_fd_sc_hd__and2_1 _5333_ (.A(\i_tinyqv.cpu.i_core.time_hi[0] ),
    .B(_2074_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2075_));
 sky130_fd_sc_hd__o21ai_1 _5334_ (.A1(net246),
    .A2(_2074_),
    .B1(_2049_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2076_));
 sky130_fd_sc_hd__nor2_1 _5335_ (.A(_2075_),
    .B(_2076_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0092_));
 sky130_fd_sc_hd__and3_1 _5336_ (.A(\i_tinyqv.cpu.i_core.time_hi[1] ),
    .B(\i_tinyqv.cpu.i_core.time_hi[0] ),
    .C(_2074_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2077_));
 sky130_fd_sc_hd__o21ai_1 _5337_ (.A1(net218),
    .A2(_2075_),
    .B1(_2049_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2078_));
 sky130_fd_sc_hd__nor2_1 _5338_ (.A(_2077_),
    .B(_2078_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0093_));
 sky130_fd_sc_hd__clkbuf_4 _5339_ (.A(_1752_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2079_));
 sky130_fd_sc_hd__o21ai_1 _5340_ (.A1(net108),
    .A2(_2077_),
    .B1(_2079_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2080_));
 sky130_fd_sc_hd__a21oi_1 _5341_ (.A1(net108),
    .A2(_2077_),
    .B1(_2080_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0094_));
 sky130_fd_sc_hd__nand2_1 _5342_ (.A(_0956_),
    .B(_1619_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2081_));
 sky130_fd_sc_hd__or3_1 _5343_ (.A(_1400_),
    .B(\i_tinyqv.cpu.i_core.is_double_fault_r ),
    .C(_2070_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2082_));
 sky130_fd_sc_hd__clkbuf_4 _5344_ (.A(_2082_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2083_));
 sky130_fd_sc_hd__nor2_1 _5345_ (.A(_2081_),
    .B(_2083_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2084_));
 sky130_fd_sc_hd__mux2_1 _5346_ (.A0(net250),
    .A1(\i_tinyqv.cpu.i_core.interrupt_req[0] ),
    .S(_2084_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2085_));
 sky130_fd_sc_hd__clkbuf_1 _5347_ (.A(net251),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0095_));
 sky130_fd_sc_hd__mux2_1 _5348_ (.A0(\i_tinyqv.cpu.i_core.last_interrupt_req[1] ),
    .A1(\i_tinyqv.cpu.i_core.interrupt_req[1] ),
    .S(_2084_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2086_));
 sky130_fd_sc_hd__clkbuf_1 _5349_ (.A(_2086_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0096_));
 sky130_fd_sc_hd__nor2_2 _5350_ (.A(_2066_),
    .B(_0840_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2087_));
 sky130_fd_sc_hd__or2_2 _5351_ (.A(_1124_),
    .B(_0855_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2088_));
 sky130_fd_sc_hd__nor3_1 _5352_ (.A(_0937_),
    .B(_0922_),
    .C(_2088_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2089_));
 sky130_fd_sc_hd__or2_1 _5353_ (.A(\i_tinyqv.cpu.i_core.mepc[0] ),
    .B(net18),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2090_));
 sky130_fd_sc_hd__a21oi_1 _5354_ (.A1(_1312_),
    .A2(net18),
    .B1(_2056_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2091_));
 sky130_fd_sc_hd__a22o_1 _5355_ (.A1(_0729_),
    .A2(_2056_),
    .B1(_2090_),
    .B2(_2091_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2092_));
 sky130_fd_sc_hd__a22o_1 _5356_ (.A1(net244),
    .A2(_0840_),
    .B1(_2087_),
    .B2(_2092_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0097_));
 sky130_fd_sc_hd__nor2_1 _5357_ (.A(\i_tinyqv.cpu.i_core.mepc[1] ),
    .B(net18),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2093_));
 sky130_fd_sc_hd__a211o_1 _5358_ (.A1(net66),
    .A2(net18),
    .B1(_2093_),
    .C1(_2056_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2094_));
 sky130_fd_sc_hd__o21ai_1 _5359_ (.A1(_0754_),
    .A2(_1395_),
    .B1(_2094_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2095_));
 sky130_fd_sc_hd__a22o_1 _5360_ (.A1(net222),
    .A2(_0840_),
    .B1(_2087_),
    .B2(_2095_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0098_));
 sky130_fd_sc_hd__nor2_1 _5361_ (.A(\i_tinyqv.cpu.i_core.mepc[2] ),
    .B(net18),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2096_));
 sky130_fd_sc_hd__a211o_1 _5362_ (.A1(_0798_),
    .A2(net18),
    .B1(_2096_),
    .C1(_2056_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2097_));
 sky130_fd_sc_hd__o21ai_1 _5363_ (.A1(_0788_),
    .A2(_1395_),
    .B1(_2097_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2098_));
 sky130_fd_sc_hd__a22o_1 _5364_ (.A1(net223),
    .A2(_0840_),
    .B1(_2087_),
    .B2(_2098_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0099_));
 sky130_fd_sc_hd__or2b_1 _5365_ (.A(net43),
    .B_N(_2089_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2099_));
 sky130_fd_sc_hd__o21a_1 _5366_ (.A1(\i_tinyqv.cpu.i_core.mepc[3] ),
    .A2(net18),
    .B1(_1395_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2100_));
 sky130_fd_sc_hd__a22o_1 _5367_ (.A1(_0623_),
    .A2(_2056_),
    .B1(_2099_),
    .B2(_2100_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2101_));
 sky130_fd_sc_hd__a22o_1 _5368_ (.A1(net211),
    .A2(_0840_),
    .B1(_2087_),
    .B2(_2101_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0100_));
 sky130_fd_sc_hd__a21o_1 _5369_ (.A1(_0656_),
    .A2(net69),
    .B1(_1185_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2102_));
 sky130_fd_sc_hd__and2b_1 _5370_ (.A_N(_2102_),
    .B(net41),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2103_));
 sky130_fd_sc_hd__mux2_1 _5371_ (.A0(\i_tinyqv.cpu.i_core.mstatus_mie ),
    .A1(_2103_),
    .S(_2057_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2104_));
 sky130_fd_sc_hd__and3_1 _5372_ (.A(\i_tinyqv.cpu.i_core.imm_lo[8] ),
    .B(\i_tinyqv.cpu.i_core.imm_lo[9] ),
    .C(_1392_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2105_));
 sky130_fd_sc_hd__clkbuf_4 _5373_ (.A(_2105_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2106_));
 sky130_fd_sc_hd__clkbuf_4 _5374_ (.A(_2106_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2107_));
 sky130_fd_sc_hd__o21ai_1 _5375_ (.A1(_0844_),
    .A2(_0652_),
    .B1(_0920_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2108_));
 sky130_fd_sc_hd__o41a_1 _5376_ (.A1(_0939_),
    .A2(_1348_),
    .A3(_2107_),
    .A4(_2108_),
    .B1(_2057_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2109_));
 sky130_fd_sc_hd__mux2_1 _5377_ (.A0(_2104_),
    .A1(\i_tinyqv.cpu.i_core.mstatus_mpie ),
    .S(_2109_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2110_));
 sky130_fd_sc_hd__and2b_1 _5378_ (.A_N(_2083_),
    .B(_2110_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2111_));
 sky130_fd_sc_hd__clkbuf_1 _5379_ (.A(_2111_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0101_));
 sky130_fd_sc_hd__or3_1 _5380_ (.A(_1026_),
    .B(_1348_),
    .C(_2108_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2112_));
 sky130_fd_sc_hd__mux2_1 _5381_ (.A0(_2103_),
    .A1(\i_tinyqv.cpu.i_core.mstatus_mie ),
    .S(_2112_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2113_));
 sky130_fd_sc_hd__or2_1 _5382_ (.A(_2107_),
    .B(_2113_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2114_));
 sky130_fd_sc_hd__or2_1 _5383_ (.A(net262),
    .B(_1393_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2115_));
 sky130_fd_sc_hd__a31o_1 _5384_ (.A1(_2057_),
    .A2(_2114_),
    .A3(_2115_),
    .B1(_2083_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0102_));
 sky130_fd_sc_hd__o21a_1 _5385_ (.A1(\i_tinyqv.cpu.i_core.mstatus_mte ),
    .A2(_2107_),
    .B1(_2057_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2116_));
 sky130_fd_sc_hd__or2_1 _5386_ (.A(_2083_),
    .B(_2116_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2117_));
 sky130_fd_sc_hd__clkbuf_1 _5387_ (.A(_2117_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0103_));
 sky130_fd_sc_hd__inv_2 _5388_ (.A(_1486_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2118_));
 sky130_fd_sc_hd__or2_1 _5389_ (.A(_1469_),
    .B(_2118_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2119_));
 sky130_fd_sc_hd__nor2_1 _5390_ (.A(_1483_),
    .B(_2119_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2120_));
 sky130_fd_sc_hd__buf_2 _5391_ (.A(_2120_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2121_));
 sky130_fd_sc_hd__or2_2 _5392_ (.A(_1469_),
    .B(_1486_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2122_));
 sky130_fd_sc_hd__clkbuf_4 _5393_ (.A(_1481_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2123_));
 sky130_fd_sc_hd__clkbuf_4 _5394_ (.A(_1476_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2124_));
 sky130_fd_sc_hd__nand2_1 _5395_ (.A(_2123_),
    .B(_2124_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2125_));
 sky130_fd_sc_hd__nor2_2 _5396_ (.A(_2122_),
    .B(_2125_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2126_));
 sky130_fd_sc_hd__nand2_1 _5397_ (.A(_1420_),
    .B(_2118_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2127_));
 sky130_fd_sc_hd__or2_2 _5398_ (.A(_1426_),
    .B(_2127_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2128_));
 sky130_fd_sc_hd__nor2_1 _5399_ (.A(_1483_),
    .B(_2128_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2129_));
 sky130_fd_sc_hd__o21bai_2 _5400_ (.A1(_2123_),
    .A2(_2122_),
    .B1_N(_2129_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2130_));
 sky130_fd_sc_hd__nor2_1 _5401_ (.A(_1477_),
    .B(_1488_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2131_));
 sky130_fd_sc_hd__nor2_1 _5402_ (.A(_1426_),
    .B(_2127_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2132_));
 sky130_fd_sc_hd__and2_1 _5403_ (.A(_2124_),
    .B(_2132_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2133_));
 sky130_fd_sc_hd__or4_1 _5404_ (.A(_2126_),
    .B(_2130_),
    .C(_2131_),
    .D(_2133_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2134_));
 sky130_fd_sc_hd__nor2_1 _5405_ (.A(_1452_),
    .B(_1493_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2135_));
 sky130_fd_sc_hd__o21ai_1 _5406_ (.A1(_1490_),
    .A2(_2135_),
    .B1(_1427_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2136_));
 sky130_fd_sc_hd__or3_1 _5407_ (.A(_2121_),
    .B(_2134_),
    .C(_2136_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2137_));
 sky130_fd_sc_hd__nand2_1 _5408_ (.A(_1490_),
    .B(_2128_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2138_));
 sky130_fd_sc_hd__nor2_1 _5409_ (.A(_2134_),
    .B(_2138_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2139_));
 sky130_fd_sc_hd__clkbuf_4 _5410_ (.A(_1427_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2140_));
 sky130_fd_sc_hd__o211a_1 _5411_ (.A1(_1469_),
    .A2(_2124_),
    .B1(_2139_),
    .C1(_2140_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2141_));
 sky130_fd_sc_hd__nor2_1 _5412_ (.A(_1490_),
    .B(_1507_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2142_));
 sky130_fd_sc_hd__nor2_4 _5413_ (.A(_1477_),
    .B(_2128_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2143_));
 sky130_fd_sc_hd__a221o_1 _5414_ (.A1(_1478_),
    .A2(_2118_),
    .B1(_2135_),
    .B2(_2142_),
    .C1(_2143_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2144_));
 sky130_fd_sc_hd__a221o_1 _5415_ (.A1(_1510_),
    .A2(_2137_),
    .B1(_2141_),
    .B2(_1460_),
    .C1(_2144_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2145_));
 sky130_fd_sc_hd__or2b_1 _5416_ (.A(_1439_),
    .B_N(_1440_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2146_));
 sky130_fd_sc_hd__clkbuf_4 _5417_ (.A(_2146_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2147_));
 sky130_fd_sc_hd__mux2_1 _5418_ (.A0(_1640_),
    .A1(_2145_),
    .S(_2147_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2148_));
 sky130_fd_sc_hd__and3_2 _5419_ (.A(_0837_),
    .B(_0863_),
    .C(_1440_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2149_));
 sky130_fd_sc_hd__nor2_1 _5420_ (.A(_1405_),
    .B(_1438_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2150_));
 sky130_fd_sc_hd__o21a_1 _5421_ (.A1(_1399_),
    .A2(_1443_),
    .B1(_2150_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2151_));
 sky130_fd_sc_hd__or2_2 _5422_ (.A(_2149_),
    .B(_2151_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2152_));
 sky130_fd_sc_hd__nand2_4 _5423_ (.A(_1752_),
    .B(_2152_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2153_));
 sky130_fd_sc_hd__mux2_1 _5424_ (.A0(_2148_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.rd[0] ),
    .S(_2153_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2154_));
 sky130_fd_sc_hd__clkbuf_1 _5425_ (.A(_2154_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0104_));
 sky130_fd_sc_hd__buf_2 _5426_ (.A(_1448_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2155_));
 sky130_fd_sc_hd__a221o_1 _5427_ (.A1(_1514_),
    .A2(_2137_),
    .B1(_2141_),
    .B2(_2155_),
    .C1(_2149_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2156_));
 sky130_fd_sc_hd__o31a_1 _5428_ (.A1(_2147_),
    .A2(_1641_),
    .A3(_1647_),
    .B1(_2156_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2157_));
 sky130_fd_sc_hd__mux2_1 _5429_ (.A0(_2157_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.rd[1] ),
    .S(_2153_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2158_));
 sky130_fd_sc_hd__clkbuf_1 _5430_ (.A(_2158_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0105_));
 sky130_fd_sc_hd__a21o_1 _5431_ (.A1(\i_tinyqv.cpu.i_core.i_registers.rd[1] ),
    .A2(\i_tinyqv.cpu.i_core.i_registers.rd[0] ),
    .B1(\i_tinyqv.cpu.i_core.i_registers.rd[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2159_));
 sky130_fd_sc_hd__a21o_1 _5432_ (.A1(_1679_),
    .A2(_2159_),
    .B1(_2147_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2160_));
 sky130_fd_sc_hd__a221o_1 _5433_ (.A1(_1501_),
    .A2(_2137_),
    .B1(_2141_),
    .B2(_1491_),
    .C1(_2149_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2161_));
 sky130_fd_sc_hd__and4_1 _5434_ (.A(_1752_),
    .B(_2152_),
    .C(_2160_),
    .D(_2161_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2162_));
 sky130_fd_sc_hd__a21o_1 _5435_ (.A1(\i_tinyqv.cpu.i_core.i_registers.rd[2] ),
    .A2(_2153_),
    .B1(_2162_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0106_));
 sky130_fd_sc_hd__o21ai_1 _5436_ (.A1(\i_tinyqv.cpu.i_core.i_registers.rd[3] ),
    .A2(_1679_),
    .B1(_2149_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2163_));
 sky130_fd_sc_hd__a21oi_1 _5437_ (.A1(\i_tinyqv.cpu.i_core.i_registers.rd[3] ),
    .A2(_1679_),
    .B1(_2163_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2164_));
 sky130_fd_sc_hd__clkbuf_4 _5438_ (.A(_1498_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2165_));
 sky130_fd_sc_hd__o31a_1 _5439_ (.A1(_2134_),
    .A2(_2136_),
    .A3(_2143_),
    .B1(_2165_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2166_));
 sky130_fd_sc_hd__or4_1 _5440_ (.A(_2149_),
    .B(_2121_),
    .C(_2141_),
    .D(_2166_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2167_));
 sky130_fd_sc_hd__or3b_1 _5441_ (.A(_2164_),
    .B(_2153_),
    .C_N(_2167_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2168_));
 sky130_fd_sc_hd__a21bo_1 _5442_ (.A1(net252),
    .A2(_2153_),
    .B1_N(_2168_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0107_));
 sky130_fd_sc_hd__nand3_4 _5443_ (.A(_0997_),
    .B(_0991_),
    .C(_1725_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2169_));
 sky130_fd_sc_hd__o21ai_1 _5444_ (.A1(\i_uart_tx.fsm_state[2] ),
    .A2(\i_uart_tx.fsm_state[1] ),
    .B1(\i_uart_tx.fsm_state[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2170_));
 sky130_fd_sc_hd__nand2_1 _5445_ (.A(net206),
    .B(\i_uart_tx.cycle_counter[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2171_));
 sky130_fd_sc_hd__or4bb_1 _5446_ (.A(\i_uart_tx.cycle_counter[6] ),
    .B(\i_uart_tx.cycle_counter[4] ),
    .C_N(\i_uart_tx.cycle_counter[3] ),
    .D_N(\i_uart_tx.cycle_counter[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2172_));
 sky130_fd_sc_hd__or4b_1 _5447_ (.A(\i_uart_tx.cycle_counter[10] ),
    .B(\i_uart_tx.cycle_counter[8] ),
    .C(\i_uart_tx.cycle_counter[7] ),
    .D_N(\i_uart_tx.cycle_counter[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2173_));
 sky130_fd_sc_hd__or4_1 _5448_ (.A(\i_uart_tx.cycle_counter[2] ),
    .B(_2171_),
    .C(_2172_),
    .D(_2173_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2174_));
 sky130_fd_sc_hd__inv_2 _5449_ (.A(_2174_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2175_));
 sky130_fd_sc_hd__and3_1 _5450_ (.A(_0990_),
    .B(_2170_),
    .C(_2175_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2176_));
 sky130_fd_sc_hd__clkbuf_4 _5451_ (.A(_2176_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2177_));
 sky130_fd_sc_hd__mux2_1 _5452_ (.A0(\i_uart_tx.data_to_send[0] ),
    .A1(\i_uart_tx.data_to_send[1] ),
    .S(_2177_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2178_));
 sky130_fd_sc_hd__and3_2 _5453_ (.A(_0997_),
    .B(_0991_),
    .C(_1557_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2179_));
 sky130_fd_sc_hd__or2_1 _5454_ (.A(_2178_),
    .B(_2179_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2180_));
 sky130_fd_sc_hd__clkbuf_4 _5455_ (.A(_1728_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2181_));
 sky130_fd_sc_hd__clkbuf_4 _5456_ (.A(_2181_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2182_));
 sky130_fd_sc_hd__o211a_1 _5457_ (.A1(net117),
    .A2(_2169_),
    .B1(_2180_),
    .C1(_2182_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0108_));
 sky130_fd_sc_hd__mux2_1 _5458_ (.A0(\i_uart_tx.data_to_send[1] ),
    .A1(\i_uart_tx.data_to_send[2] ),
    .S(_2177_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2183_));
 sky130_fd_sc_hd__or2_1 _5459_ (.A(_2179_),
    .B(_2183_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2184_));
 sky130_fd_sc_hd__o211a_1 _5460_ (.A1(net97),
    .A2(_2169_),
    .B1(_2184_),
    .C1(_2182_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0109_));
 sky130_fd_sc_hd__mux2_1 _5461_ (.A0(\i_uart_tx.data_to_send[2] ),
    .A1(\i_uart_tx.data_to_send[3] ),
    .S(_2177_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2185_));
 sky130_fd_sc_hd__or2_1 _5462_ (.A(_2179_),
    .B(_2185_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2186_));
 sky130_fd_sc_hd__o211a_1 _5463_ (.A1(net98),
    .A2(_2169_),
    .B1(_2186_),
    .C1(_2182_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0110_));
 sky130_fd_sc_hd__mux2_1 _5464_ (.A0(\i_uart_tx.data_to_send[3] ),
    .A1(\i_uart_tx.data_to_send[4] ),
    .S(_2177_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2187_));
 sky130_fd_sc_hd__or2_1 _5465_ (.A(_2179_),
    .B(_2187_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2188_));
 sky130_fd_sc_hd__o211a_1 _5466_ (.A1(\i_debug_uart_tx.uart_tx_data[3] ),
    .A2(_2169_),
    .B1(_2188_),
    .C1(_2182_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0111_));
 sky130_fd_sc_hd__mux2_1 _5467_ (.A0(\i_uart_tx.data_to_send[4] ),
    .A1(\i_uart_tx.data_to_send[5] ),
    .S(_2177_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2189_));
 sky130_fd_sc_hd__or2_1 _5468_ (.A(_2179_),
    .B(_2189_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2190_));
 sky130_fd_sc_hd__o211a_1 _5469_ (.A1(\i_debug_uart_tx.uart_tx_data[4] ),
    .A2(_2169_),
    .B1(_2190_),
    .C1(_2182_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0112_));
 sky130_fd_sc_hd__mux2_1 _5470_ (.A0(\i_uart_tx.data_to_send[5] ),
    .A1(\i_uart_tx.data_to_send[6] ),
    .S(_2177_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2191_));
 sky130_fd_sc_hd__or2_1 _5471_ (.A(_2179_),
    .B(_2191_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2192_));
 sky130_fd_sc_hd__o211a_1 _5472_ (.A1(\i_debug_uart_tx.uart_tx_data[5] ),
    .A2(_2169_),
    .B1(_2192_),
    .C1(_2182_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0113_));
 sky130_fd_sc_hd__mux2_1 _5473_ (.A0(\i_uart_tx.data_to_send[6] ),
    .A1(\i_uart_tx.data_to_send[7] ),
    .S(_2177_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2193_));
 sky130_fd_sc_hd__or2_1 _5474_ (.A(_2179_),
    .B(_2193_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2194_));
 sky130_fd_sc_hd__o211a_1 _5475_ (.A1(net316),
    .A2(_2169_),
    .B1(_2194_),
    .C1(_2182_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0114_));
 sky130_fd_sc_hd__inv_2 _5476_ (.A(_2177_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2195_));
 sky130_fd_sc_hd__a21o_1 _5477_ (.A1(\i_uart_tx.data_to_send[7] ),
    .A2(_2195_),
    .B1(_2179_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2196_));
 sky130_fd_sc_hd__o211a_1 _5478_ (.A1(\i_debug_uart_tx.uart_tx_data[7] ),
    .A2(_2169_),
    .B1(_2196_),
    .C1(_2182_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0115_));
 sky130_fd_sc_hd__or2_2 _5479_ (.A(\i_uart_tx.fsm_state[0] ),
    .B(_0990_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2197_));
 sky130_fd_sc_hd__inv_2 _5480_ (.A(\i_debug_uart_tx.resetn ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2198_));
 sky130_fd_sc_hd__nor2_1 _5481_ (.A(_2198_),
    .B(_2175_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2199_));
 sky130_fd_sc_hd__buf_2 _5482_ (.A(_2199_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2200_));
 sky130_fd_sc_hd__a21boi_1 _5483_ (.A1(\i_uart_tx.cycle_counter[0] ),
    .A2(_2197_),
    .B1_N(_2200_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2201_));
 sky130_fd_sc_hd__o21a_1 _5484_ (.A1(\i_uart_tx.cycle_counter[0] ),
    .A2(_2197_),
    .B1(_2201_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0116_));
 sky130_fd_sc_hd__a21o_1 _5485_ (.A1(\i_uart_tx.cycle_counter[0] ),
    .A2(_2197_),
    .B1(net206),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2202_));
 sky130_fd_sc_hd__o211a_1 _5486_ (.A1(_0991_),
    .A2(_2171_),
    .B1(_2200_),
    .C1(_2202_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0117_));
 sky130_fd_sc_hd__and4_1 _5487_ (.A(\i_uart_tx.cycle_counter[2] ),
    .B(net206),
    .C(\i_uart_tx.cycle_counter[0] ),
    .D(_2197_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2203_));
 sky130_fd_sc_hd__a31o_1 _5488_ (.A1(net206),
    .A2(\i_uart_tx.cycle_counter[0] ),
    .A3(_2197_),
    .B1(\i_uart_tx.cycle_counter[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2204_));
 sky130_fd_sc_hd__and3b_1 _5489_ (.A_N(_2203_),
    .B(_2200_),
    .C(_2204_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2205_));
 sky130_fd_sc_hd__clkbuf_1 _5490_ (.A(_2205_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0118_));
 sky130_fd_sc_hd__and2_1 _5491_ (.A(\i_uart_tx.cycle_counter[3] ),
    .B(_2203_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2206_));
 sky130_fd_sc_hd__o21ai_1 _5492_ (.A1(net219),
    .A2(_2203_),
    .B1(_2200_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2207_));
 sky130_fd_sc_hd__nor2_1 _5493_ (.A(_2206_),
    .B(_2207_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0119_));
 sky130_fd_sc_hd__o21ai_1 _5494_ (.A1(\i_uart_tx.cycle_counter[4] ),
    .A2(_2206_),
    .B1(_2200_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2208_));
 sky130_fd_sc_hd__a21oi_1 _5495_ (.A1(net174),
    .A2(_2206_),
    .B1(_2208_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0120_));
 sky130_fd_sc_hd__and3_1 _5496_ (.A(\i_uart_tx.cycle_counter[5] ),
    .B(\i_uart_tx.cycle_counter[4] ),
    .C(_2206_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2209_));
 sky130_fd_sc_hd__a31o_1 _5497_ (.A1(\i_uart_tx.cycle_counter[4] ),
    .A2(\i_uart_tx.cycle_counter[3] ),
    .A3(_2203_),
    .B1(\i_uart_tx.cycle_counter[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2210_));
 sky130_fd_sc_hd__and3b_1 _5498_ (.A_N(_2209_),
    .B(_2199_),
    .C(_2210_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2211_));
 sky130_fd_sc_hd__clkbuf_1 _5499_ (.A(_2211_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0121_));
 sky130_fd_sc_hd__and2_1 _5500_ (.A(\i_uart_tx.cycle_counter[6] ),
    .B(_2209_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2212_));
 sky130_fd_sc_hd__o21ai_1 _5501_ (.A1(net214),
    .A2(_2209_),
    .B1(_2200_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2213_));
 sky130_fd_sc_hd__nor2_1 _5502_ (.A(_2212_),
    .B(_2213_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0122_));
 sky130_fd_sc_hd__o21ai_1 _5503_ (.A1(net157),
    .A2(_2212_),
    .B1(_2200_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2214_));
 sky130_fd_sc_hd__a21oi_1 _5504_ (.A1(net157),
    .A2(_2212_),
    .B1(_2214_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0123_));
 sky130_fd_sc_hd__and3_1 _5505_ (.A(net170),
    .B(net157),
    .C(_2212_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2215_));
 sky130_fd_sc_hd__a31o_1 _5506_ (.A1(\i_uart_tx.cycle_counter[7] ),
    .A2(\i_uart_tx.cycle_counter[6] ),
    .A3(_2209_),
    .B1(\i_uart_tx.cycle_counter[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2216_));
 sky130_fd_sc_hd__and3b_1 _5507_ (.A_N(_2215_),
    .B(_2199_),
    .C(_2216_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2217_));
 sky130_fd_sc_hd__clkbuf_1 _5508_ (.A(_2217_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0124_));
 sky130_fd_sc_hd__and2_1 _5509_ (.A(\i_uart_tx.cycle_counter[9] ),
    .B(_2215_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2218_));
 sky130_fd_sc_hd__o21ai_1 _5510_ (.A1(\i_uart_tx.cycle_counter[9] ),
    .A2(_2215_),
    .B1(_2200_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2219_));
 sky130_fd_sc_hd__nor2_1 _5511_ (.A(_2218_),
    .B(net171),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0125_));
 sky130_fd_sc_hd__o21ai_1 _5512_ (.A1(net102),
    .A2(_2218_),
    .B1(_2200_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2220_));
 sky130_fd_sc_hd__a21oi_1 _5513_ (.A1(net102),
    .A2(_2218_),
    .B1(_2220_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0126_));
 sky130_fd_sc_hd__clkbuf_4 _5514_ (.A(_1728_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2221_));
 sky130_fd_sc_hd__inv_2 _5515_ (.A(\i_uart_tx.fsm_state[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2222_));
 sky130_fd_sc_hd__a31oi_1 _5516_ (.A1(\i_uart_tx.fsm_state[3] ),
    .A2(_2222_),
    .A3(\i_uart_tx.fsm_state[1] ),
    .B1(\i_uart_tx.fsm_state[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2223_));
 sky130_fd_sc_hd__a21o_1 _5517_ (.A1(_0990_),
    .A2(_2223_),
    .B1(_2179_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2224_));
 sky130_fd_sc_hd__nand2_1 _5518_ (.A(_2197_),
    .B(_2174_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2225_));
 sky130_fd_sc_hd__a32o_1 _5519_ (.A1(_2221_),
    .A2(_2224_),
    .A3(_2225_),
    .B1(_2200_),
    .B2(net270),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0127_));
 sky130_fd_sc_hd__nand3b_1 _5520_ (.A_N(_2223_),
    .B(_2225_),
    .C(\i_uart_tx.fsm_state[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2226_));
 sky130_fd_sc_hd__a21o_1 _5521_ (.A1(\i_uart_tx.fsm_state[0] ),
    .A2(_2225_),
    .B1(\i_uart_tx.fsm_state[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2227_));
 sky130_fd_sc_hd__and3_1 _5522_ (.A(_2181_),
    .B(_2226_),
    .C(_2227_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2228_));
 sky130_fd_sc_hd__clkbuf_1 _5523_ (.A(_2228_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0128_));
 sky130_fd_sc_hd__clkbuf_4 _5524_ (.A(_2198_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2229_));
 sky130_fd_sc_hd__and3_1 _5525_ (.A(\i_uart_tx.fsm_state[1] ),
    .B(\i_uart_tx.fsm_state[0] ),
    .C(_2175_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2230_));
 sky130_fd_sc_hd__xnor2_1 _5526_ (.A(\i_uart_tx.fsm_state[2] ),
    .B(_2230_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2231_));
 sky130_fd_sc_hd__nor2_1 _5527_ (.A(_2229_),
    .B(_2231_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0129_));
 sky130_fd_sc_hd__a21oi_1 _5528_ (.A1(net164),
    .A2(_2230_),
    .B1(\i_uart_tx.fsm_state[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2232_));
 sky130_fd_sc_hd__xnor2_1 _5529_ (.A(\i_uart_tx.fsm_state[2] ),
    .B(\i_uart_tx.fsm_state[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2233_));
 sky130_fd_sc_hd__a41o_1 _5530_ (.A1(\i_uart_tx.fsm_state[3] ),
    .A2(\i_uart_tx.fsm_state[1] ),
    .A3(_2225_),
    .A4(_2233_),
    .B1(_2198_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2234_));
 sky130_fd_sc_hd__nor2_1 _5531_ (.A(net165),
    .B(_2234_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0130_));
 sky130_fd_sc_hd__and4bb_1 _5532_ (.A_N(\i_uart_rx.cycle_counter[2] ),
    .B_N(\i_uart_rx.cycle_counter[4] ),
    .C(\i_uart_rx.cycle_counter[5] ),
    .D(\i_uart_rx.cycle_counter[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2235_));
 sky130_fd_sc_hd__and2_1 _5533_ (.A(net91),
    .B(\i_uart_rx.cycle_counter[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2236_));
 sky130_fd_sc_hd__and4bb_1 _5534_ (.A_N(\i_uart_rx.cycle_counter[7] ),
    .B_N(\i_uart_rx.cycle_counter[6] ),
    .C(_2235_),
    .D(_2236_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2237_));
 sky130_fd_sc_hd__and4bb_4 _5535_ (.A_N(\i_uart_rx.cycle_counter[8] ),
    .B_N(\i_uart_rx.cycle_counter[10] ),
    .C(_2237_),
    .D(\i_uart_rx.cycle_counter[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2238_));
 sky130_fd_sc_hd__or3_4 _5536_ (.A(\i_uart_rx.fsm_state[3] ),
    .B(\i_uart_rx.fsm_state[2] ),
    .C(\i_uart_rx.fsm_state[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2239_));
 sky130_fd_sc_hd__o21a_2 _5537_ (.A1(\i_uart_rx.fsm_state[0] ),
    .A2(_2239_),
    .B1(_1728_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2240_));
 sky130_fd_sc_hd__nor3b_1 _5538_ (.A(_1228_),
    .B(_2238_),
    .C_N(_2240_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2241_));
 sky130_fd_sc_hd__buf_2 _5539_ (.A(net17),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2242_));
 sky130_fd_sc_hd__and2b_1 _5540_ (.A_N(\i_uart_rx.cycle_counter[0] ),
    .B(_2242_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2243_));
 sky130_fd_sc_hd__clkbuf_1 _5541_ (.A(_2243_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0131_));
 sky130_fd_sc_hd__o21ai_1 _5542_ (.A1(net91),
    .A2(net307),
    .B1(_2242_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2244_));
 sky130_fd_sc_hd__nor2_1 _5543_ (.A(_2236_),
    .B(_2244_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0132_));
 sky130_fd_sc_hd__o21ai_1 _5544_ (.A1(net178),
    .A2(_2236_),
    .B1(_2242_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2245_));
 sky130_fd_sc_hd__a21oi_1 _5545_ (.A1(net178),
    .A2(_2236_),
    .B1(_2245_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0133_));
 sky130_fd_sc_hd__and3_1 _5546_ (.A(\i_uart_rx.cycle_counter[3] ),
    .B(\i_uart_rx.cycle_counter[2] ),
    .C(_2236_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2246_));
 sky130_fd_sc_hd__a31o_1 _5547_ (.A1(net91),
    .A2(\i_uart_rx.cycle_counter[1] ),
    .A3(net224),
    .B1(\i_uart_rx.cycle_counter[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2247_));
 sky130_fd_sc_hd__and3b_1 _5548_ (.A_N(_2246_),
    .B(_2247_),
    .C(net17),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2248_));
 sky130_fd_sc_hd__clkbuf_1 _5549_ (.A(_2248_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0134_));
 sky130_fd_sc_hd__and2_1 _5550_ (.A(net148),
    .B(_2246_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2249_));
 sky130_fd_sc_hd__o21ai_1 _5551_ (.A1(net148),
    .A2(_2246_),
    .B1(_2242_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2250_));
 sky130_fd_sc_hd__nor2_1 _5552_ (.A(_2249_),
    .B(_2250_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0135_));
 sky130_fd_sc_hd__and3_1 _5553_ (.A(\i_uart_rx.cycle_counter[5] ),
    .B(net148),
    .C(_2246_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2251_));
 sky130_fd_sc_hd__o21ai_1 _5554_ (.A1(net306),
    .A2(_2249_),
    .B1(_2242_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2252_));
 sky130_fd_sc_hd__nor2_1 _5555_ (.A(_2251_),
    .B(_2252_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0136_));
 sky130_fd_sc_hd__and2_1 _5556_ (.A(\i_uart_rx.cycle_counter[6] ),
    .B(_2251_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2253_));
 sky130_fd_sc_hd__o21ai_1 _5557_ (.A1(\i_uart_rx.cycle_counter[6] ),
    .A2(_2251_),
    .B1(_2242_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2254_));
 sky130_fd_sc_hd__nor2_1 _5558_ (.A(_2253_),
    .B(_2254_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0137_));
 sky130_fd_sc_hd__o21ai_1 _5559_ (.A1(\i_uart_rx.cycle_counter[7] ),
    .A2(_2253_),
    .B1(_2242_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2255_));
 sky130_fd_sc_hd__a21oi_1 _5560_ (.A1(net199),
    .A2(_2253_),
    .B1(_2255_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0138_));
 sky130_fd_sc_hd__and3_1 _5561_ (.A(\i_uart_rx.cycle_counter[7] ),
    .B(\i_uart_rx.cycle_counter[8] ),
    .C(_2253_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2256_));
 sky130_fd_sc_hd__a31o_1 _5562_ (.A1(\i_uart_rx.cycle_counter[7] ),
    .A2(\i_uart_rx.cycle_counter[6] ),
    .A3(_2251_),
    .B1(\i_uart_rx.cycle_counter[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2257_));
 sky130_fd_sc_hd__and3b_1 _5563_ (.A_N(_2256_),
    .B(_2242_),
    .C(_2257_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2258_));
 sky130_fd_sc_hd__clkbuf_1 _5564_ (.A(_2258_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0139_));
 sky130_fd_sc_hd__and2_1 _5565_ (.A(\i_uart_rx.cycle_counter[9] ),
    .B(_2256_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2259_));
 sky130_fd_sc_hd__o21ai_1 _5566_ (.A1(net247),
    .A2(_2256_),
    .B1(_2242_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2260_));
 sky130_fd_sc_hd__nor2_1 _5567_ (.A(_2259_),
    .B(_2260_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0140_));
 sky130_fd_sc_hd__o21ai_1 _5568_ (.A1(net142),
    .A2(_2259_),
    .B1(_2242_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2261_));
 sky130_fd_sc_hd__a21oi_1 _5569_ (.A1(net142),
    .A2(_2259_),
    .B1(_2261_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0141_));
 sky130_fd_sc_hd__o21ai_2 _5570_ (.A1(\i_uart_rx.fsm_state[2] ),
    .A2(\i_uart_rx.fsm_state[1] ),
    .B1(\i_uart_rx.fsm_state[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2262_));
 sky130_fd_sc_hd__nand3_4 _5571_ (.A(_2239_),
    .B(_2238_),
    .C(_2262_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2263_));
 sky130_fd_sc_hd__and3_2 _5572_ (.A(_2239_),
    .B(_2238_),
    .C(_2262_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2264_));
 sky130_fd_sc_hd__or2_1 _5573_ (.A(\i_uart_rx.recieved_data[0] ),
    .B(_2264_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2265_));
 sky130_fd_sc_hd__o211a_1 _5574_ (.A1(net201),
    .A2(_2263_),
    .B1(_2265_),
    .C1(_2240_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0142_));
 sky130_fd_sc_hd__or2_1 _5575_ (.A(\i_uart_rx.recieved_data[1] ),
    .B(_2264_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2266_));
 sky130_fd_sc_hd__o211a_1 _5576_ (.A1(net225),
    .A2(_2263_),
    .B1(_2266_),
    .C1(_2240_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0143_));
 sky130_fd_sc_hd__or2_1 _5577_ (.A(\i_uart_rx.recieved_data[2] ),
    .B(_2264_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2267_));
 sky130_fd_sc_hd__o211a_1 _5578_ (.A1(net241),
    .A2(_2263_),
    .B1(_2267_),
    .C1(_2240_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0144_));
 sky130_fd_sc_hd__or2_1 _5579_ (.A(\i_uart_rx.recieved_data[3] ),
    .B(_2264_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2268_));
 sky130_fd_sc_hd__o211a_1 _5580_ (.A1(net207),
    .A2(_2263_),
    .B1(_2268_),
    .C1(_2240_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0145_));
 sky130_fd_sc_hd__or2_1 _5581_ (.A(\i_uart_rx.recieved_data[4] ),
    .B(_2264_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2269_));
 sky130_fd_sc_hd__o211a_1 _5582_ (.A1(net160),
    .A2(_2263_),
    .B1(_2269_),
    .C1(_2240_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0146_));
 sky130_fd_sc_hd__or2_1 _5583_ (.A(\i_uart_rx.recieved_data[5] ),
    .B(_2264_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2270_));
 sky130_fd_sc_hd__o211a_1 _5584_ (.A1(net240),
    .A2(_2263_),
    .B1(_2270_),
    .C1(_2240_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0147_));
 sky130_fd_sc_hd__or2_1 _5585_ (.A(\i_uart_rx.recieved_data[6] ),
    .B(_2264_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2271_));
 sky130_fd_sc_hd__o211a_1 _5586_ (.A1(net172),
    .A2(_2263_),
    .B1(_2271_),
    .C1(_2240_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0148_));
 sky130_fd_sc_hd__or2_1 _5587_ (.A(\i_uart_rx.recieved_data[7] ),
    .B(_2264_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2272_));
 sky130_fd_sc_hd__o211a_1 _5588_ (.A1(net191),
    .A2(_2263_),
    .B1(_2272_),
    .C1(_2240_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0149_));
 sky130_fd_sc_hd__or3b_1 _5589_ (.A(\i_uart_rx.cycle_counter[9] ),
    .B(\i_uart_rx.cycle_counter[10] ),
    .C_N(\i_uart_rx.cycle_counter[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2273_));
 sky130_fd_sc_hd__or4b_1 _5590_ (.A(\i_uart_rx.cycle_counter[1] ),
    .B(\i_uart_rx.cycle_counter[7] ),
    .C(\i_uart_rx.cycle_counter[6] ),
    .D_N(\i_uart_rx.cycle_counter[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2274_));
 sky130_fd_sc_hd__or4bb_1 _5591_ (.A(\i_uart_rx.cycle_counter[3] ),
    .B(\i_uart_rx.cycle_counter[5] ),
    .C_N(\i_uart_rx.cycle_counter[4] ),
    .D_N(\i_uart_rx.cycle_counter[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2275_));
 sky130_fd_sc_hd__or3_2 _5592_ (.A(_2273_),
    .B(_2274_),
    .C(_2275_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2276_));
 sky130_fd_sc_hd__inv_2 _5593_ (.A(_2276_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2277_));
 sky130_fd_sc_hd__or2_1 _5594_ (.A(\i_uart_rx.rxd_reg[0] ),
    .B(_2276_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2278_));
 sky130_fd_sc_hd__o211a_1 _5595_ (.A1(net191),
    .A2(_2277_),
    .B1(_2278_),
    .C1(_2182_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0150_));
 sky130_fd_sc_hd__or2_1 _5596_ (.A(_2229_),
    .B(_2239_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2279_));
 sky130_fd_sc_hd__clkbuf_1 _5597_ (.A(_2279_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0151_));
 sky130_fd_sc_hd__o21ai_2 _5598_ (.A1(\i_uart_rx.fsm_state[0] ),
    .A2(_2239_),
    .B1(_1227_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2280_));
 sky130_fd_sc_hd__or2_2 _5599_ (.A(_2238_),
    .B(_2280_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2281_));
 sky130_fd_sc_hd__nand2_1 _5600_ (.A(_0997_),
    .B(_1558_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2282_));
 sky130_fd_sc_hd__nand2_1 _5601_ (.A(_1228_),
    .B(_2282_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2283_));
 sky130_fd_sc_hd__o31a_1 _5602_ (.A1(\i_uart_rx.fsm_state[0] ),
    .A2(\i_uart_rx.rxd_reg[0] ),
    .A3(_2239_),
    .B1(_2280_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2284_));
 sky130_fd_sc_hd__nor2_1 _5603_ (.A(\i_uart_rx.fsm_state[0] ),
    .B(_1227_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2285_));
 sky130_fd_sc_hd__nand3_1 _5604_ (.A(\i_uart_rx.rxd_reg[0] ),
    .B(_2277_),
    .C(_2285_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2286_));
 sky130_fd_sc_hd__a32o_1 _5605_ (.A1(_2283_),
    .A2(_2284_),
    .A3(_2286_),
    .B1(_1227_),
    .B2(\i_uart_rx.fsm_state[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2287_));
 sky130_fd_sc_hd__a21oi_1 _5606_ (.A1(_2281_),
    .A2(_2287_),
    .B1(_2229_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2288_));
 sky130_fd_sc_hd__o21a_1 _5607_ (.A1(_2281_),
    .A2(_2287_),
    .B1(_2288_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0152_));
 sky130_fd_sc_hd__nand2_1 _5608_ (.A(\i_uart_rx.fsm_state[1] ),
    .B(\i_uart_rx.fsm_state[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2289_));
 sky130_fd_sc_hd__or2_1 _5609_ (.A(\i_uart_rx.fsm_state[1] ),
    .B(\i_uart_rx.fsm_state[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2290_));
 sky130_fd_sc_hd__a22o_1 _5610_ (.A1(_1228_),
    .A2(_2282_),
    .B1(_2285_),
    .B2(_2278_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2291_));
 sky130_fd_sc_hd__inv_2 _5611_ (.A(_2281_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2292_));
 sky130_fd_sc_hd__a311o_1 _5612_ (.A1(_2289_),
    .A2(_1227_),
    .A3(_2290_),
    .B1(_2291_),
    .C1(_2292_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2293_));
 sky130_fd_sc_hd__o211a_1 _5613_ (.A1(\i_uart_rx.fsm_state[1] ),
    .A2(_2281_),
    .B1(_2293_),
    .C1(_2182_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0153_));
 sky130_fd_sc_hd__and3_1 _5614_ (.A(\i_uart_rx.fsm_state[2] ),
    .B(\i_uart_rx.fsm_state[1] ),
    .C(\i_uart_rx.fsm_state[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2294_));
 sky130_fd_sc_hd__o21ba_1 _5615_ (.A1(_2289_),
    .A2(_2292_),
    .B1_N(\i_uart_rx.fsm_state[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2295_));
 sky130_fd_sc_hd__a2111oi_1 _5616_ (.A1(_2238_),
    .A2(_2294_),
    .B1(_2280_),
    .C1(_2229_),
    .D1(_2295_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0154_));
 sky130_fd_sc_hd__xnor2_1 _5617_ (.A(\i_uart_rx.fsm_state[3] ),
    .B(_2294_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2296_));
 sky130_fd_sc_hd__a21oi_1 _5618_ (.A1(_2238_),
    .A2(_2296_),
    .B1(_2280_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2297_));
 sky130_fd_sc_hd__or2_1 _5619_ (.A(\i_uart_rx.fsm_state[3] ),
    .B(_2281_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2298_));
 sky130_fd_sc_hd__buf_2 _5620_ (.A(_1729_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2299_));
 sky130_fd_sc_hd__o211a_1 _5621_ (.A1(_2291_),
    .A2(_2297_),
    .B1(_2298_),
    .C1(_2299_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0155_));
 sky130_fd_sc_hd__or2_1 _5622_ (.A(_2229_),
    .B(net193),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2300_));
 sky130_fd_sc_hd__clkbuf_1 _5623_ (.A(_2300_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0156_));
 sky130_fd_sc_hd__or2_1 _5624_ (.A(_2229_),
    .B(net9),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2301_));
 sky130_fd_sc_hd__clkbuf_1 _5625_ (.A(_2301_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0157_));
 sky130_fd_sc_hd__inv_2 _5626_ (.A(\i_tinyqv.mem.q_ctrl.spi_clk_out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2302_));
 sky130_fd_sc_hd__a21o_1 _5627_ (.A1(_2302_),
    .A2(\i_tinyqv.mem.q_ctrl.is_writing ),
    .B1(_1543_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2303_));
 sky130_fd_sc_hd__and3b_1 _5628_ (.A_N(\i_tinyqv.mem.q_ctrl.stop_txn_reg ),
    .B(_2303_),
    .C(\i_debug_uart_tx.resetn ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2304_));
 sky130_fd_sc_hd__inv_2 _5629_ (.A(_2304_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2305_));
 sky130_fd_sc_hd__nor2_1 _5630_ (.A(_1543_),
    .B(_2305_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0158_));
 sky130_fd_sc_hd__nor2_4 _5631_ (.A(_1399_),
    .B(_1546_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2306_));
 sky130_fd_sc_hd__and4_1 _5632_ (.A(\i_tinyqv.cpu.instr_fetch_running ),
    .B(\i_tinyqv.mem.instr_active ),
    .C(_1552_),
    .D(_2306_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2307_));
 sky130_fd_sc_hd__and4_4 _5633_ (.A(\i_tinyqv.cpu.i_core.i_cycles.rstn ),
    .B(\i_tinyqv.cpu.instr_write_offset[2] ),
    .C(_1406_),
    .D(_2307_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2308_));
 sky130_fd_sc_hd__buf_4 _5634_ (.A(_2308_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2309_));
 sky130_fd_sc_hd__mux2_1 _5635_ (.A0(net263),
    .A1(\i_tinyqv.cpu.instr_data_in[2] ),
    .S(_2309_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2310_));
 sky130_fd_sc_hd__clkbuf_1 _5636_ (.A(_2310_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0159_));
 sky130_fd_sc_hd__mux2_1 _5637_ (.A0(net260),
    .A1(\i_tinyqv.cpu.instr_data_in[3] ),
    .S(_2309_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2311_));
 sky130_fd_sc_hd__clkbuf_1 _5638_ (.A(_2311_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0160_));
 sky130_fd_sc_hd__mux2_1 _5639_ (.A0(\i_tinyqv.cpu.instr_data[3][4] ),
    .A1(\i_tinyqv.cpu.instr_data_in[4] ),
    .S(_2309_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2312_));
 sky130_fd_sc_hd__clkbuf_1 _5640_ (.A(_2312_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0161_));
 sky130_fd_sc_hd__mux2_1 _5641_ (.A0(\i_tinyqv.cpu.instr_data[3][5] ),
    .A1(\i_tinyqv.cpu.instr_data_in[5] ),
    .S(_2309_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2313_));
 sky130_fd_sc_hd__clkbuf_1 _5642_ (.A(_2313_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0162_));
 sky130_fd_sc_hd__mux2_1 _5643_ (.A0(\i_tinyqv.cpu.instr_data[3][6] ),
    .A1(\i_tinyqv.cpu.instr_data_in[6] ),
    .S(_2309_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2314_));
 sky130_fd_sc_hd__clkbuf_1 _5644_ (.A(_2314_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0163_));
 sky130_fd_sc_hd__mux2_1 _5645_ (.A0(\i_tinyqv.cpu.instr_data[3][7] ),
    .A1(\i_tinyqv.cpu.instr_data_in[7] ),
    .S(_2309_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2315_));
 sky130_fd_sc_hd__clkbuf_1 _5646_ (.A(_2315_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0164_));
 sky130_fd_sc_hd__buf_2 _5647_ (.A(\i_tinyqv.cpu.instr_data_in[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2316_));
 sky130_fd_sc_hd__mux2_1 _5648_ (.A0(\i_tinyqv.cpu.instr_data[3][8] ),
    .A1(_2316_),
    .S(_2309_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2317_));
 sky130_fd_sc_hd__clkbuf_1 _5649_ (.A(_2317_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0165_));
 sky130_fd_sc_hd__clkbuf_4 _5650_ (.A(\i_tinyqv.cpu.instr_data_in[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2318_));
 sky130_fd_sc_hd__mux2_1 _5651_ (.A0(\i_tinyqv.cpu.instr_data[3][9] ),
    .A1(_2318_),
    .S(_2309_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2319_));
 sky130_fd_sc_hd__clkbuf_1 _5652_ (.A(_2319_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0166_));
 sky130_fd_sc_hd__clkbuf_4 _5653_ (.A(\i_tinyqv.cpu.instr_data_in[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2320_));
 sky130_fd_sc_hd__mux2_1 _5654_ (.A0(\i_tinyqv.cpu.instr_data[3][10] ),
    .A1(_2320_),
    .S(_2309_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2321_));
 sky130_fd_sc_hd__clkbuf_1 _5655_ (.A(_2321_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0167_));
 sky130_fd_sc_hd__clkbuf_4 _5656_ (.A(\i_tinyqv.cpu.instr_data_in[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2322_));
 sky130_fd_sc_hd__mux2_1 _5657_ (.A0(\i_tinyqv.cpu.instr_data[3][11] ),
    .A1(_2322_),
    .S(_2308_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2323_));
 sky130_fd_sc_hd__clkbuf_1 _5658_ (.A(_2323_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0168_));
 sky130_fd_sc_hd__mux2_1 _5659_ (.A0(\i_tinyqv.cpu.instr_data[3][12] ),
    .A1(_1712_),
    .S(_2308_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2324_));
 sky130_fd_sc_hd__clkbuf_1 _5660_ (.A(_2324_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0169_));
 sky130_fd_sc_hd__mux2_1 _5661_ (.A0(net272),
    .A1(_1717_),
    .S(_2308_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2325_));
 sky130_fd_sc_hd__clkbuf_1 _5662_ (.A(_2325_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0170_));
 sky130_fd_sc_hd__mux2_1 _5663_ (.A0(\i_tinyqv.cpu.instr_data[3][14] ),
    .A1(_1720_),
    .S(_2308_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2326_));
 sky130_fd_sc_hd__clkbuf_1 _5664_ (.A(_2326_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0171_));
 sky130_fd_sc_hd__mux2_1 _5665_ (.A0(net281),
    .A1(_1721_),
    .S(_2308_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2327_));
 sky130_fd_sc_hd__clkbuf_1 _5666_ (.A(_2327_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0172_));
 sky130_fd_sc_hd__nand3_1 _5667_ (.A(_0984_),
    .B(_0987_),
    .C(_1557_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2328_));
 sky130_fd_sc_hd__or3_1 _5668_ (.A(_0995_),
    .B(_0989_),
    .C(_2328_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2329_));
 sky130_fd_sc_hd__buf_2 _5669_ (.A(_2329_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2330_));
 sky130_fd_sc_hd__and3b_1 _5670_ (.A_N(\i_debug_uart_tx.cycle_counter[4] ),
    .B(\i_debug_uart_tx.cycle_counter[3] ),
    .C(\i_debug_uart_tx.cycle_counter[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2331_));
 sky130_fd_sc_hd__and3_1 _5671_ (.A(\i_debug_uart_tx.cycle_counter[2] ),
    .B(\i_debug_uart_tx.cycle_counter[0] ),
    .C(_2331_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2332_));
 sky130_fd_sc_hd__buf_2 _5672_ (.A(_2332_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2333_));
 sky130_fd_sc_hd__o21a_1 _5673_ (.A1(\i_debug_uart_tx.fsm_state[2] ),
    .A2(\i_debug_uart_tx.fsm_state[1] ),
    .B1(\i_debug_uart_tx.fsm_state[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2334_));
 sky130_fd_sc_hd__inv_2 _5674_ (.A(_2334_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2335_));
 sky130_fd_sc_hd__nand3_4 _5675_ (.A(_0988_),
    .B(_2333_),
    .C(_2335_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2336_));
 sky130_fd_sc_hd__and3_1 _5676_ (.A(_0988_),
    .B(_2333_),
    .C(_2335_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2337_));
 sky130_fd_sc_hd__and2_1 _5677_ (.A(\i_debug_uart_tx.data_to_send[1] ),
    .B(_2337_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2338_));
 sky130_fd_sc_hd__inv_2 _5678_ (.A(_0989_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2339_));
 sky130_fd_sc_hd__and3b_1 _5679_ (.A_N(_2328_),
    .B(_0969_),
    .C(_2339_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2340_));
 sky130_fd_sc_hd__buf_2 _5680_ (.A(_2340_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2341_));
 sky130_fd_sc_hd__a211o_1 _5681_ (.A1(\i_debug_uart_tx.data_to_send[0] ),
    .A2(_2336_),
    .B1(_2338_),
    .C1(_2341_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2342_));
 sky130_fd_sc_hd__o211a_1 _5682_ (.A1(net117),
    .A2(_2330_),
    .B1(_2342_),
    .C1(_2299_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0173_));
 sky130_fd_sc_hd__and2_1 _5683_ (.A(\i_debug_uart_tx.data_to_send[2] ),
    .B(_2337_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2343_));
 sky130_fd_sc_hd__a211o_1 _5684_ (.A1(net233),
    .A2(_2336_),
    .B1(_2341_),
    .C1(_2343_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2344_));
 sky130_fd_sc_hd__o211a_1 _5685_ (.A1(net97),
    .A2(_2330_),
    .B1(_2344_),
    .C1(_2299_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0174_));
 sky130_fd_sc_hd__and2_1 _5686_ (.A(\i_debug_uart_tx.data_to_send[3] ),
    .B(_2337_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2345_));
 sky130_fd_sc_hd__a211o_1 _5687_ (.A1(net255),
    .A2(_2336_),
    .B1(_2341_),
    .C1(_2345_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2346_));
 sky130_fd_sc_hd__o211a_1 _5688_ (.A1(net98),
    .A2(_2330_),
    .B1(_2346_),
    .C1(_2299_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0175_));
 sky130_fd_sc_hd__and2_1 _5689_ (.A(\i_debug_uart_tx.data_to_send[4] ),
    .B(_2337_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2347_));
 sky130_fd_sc_hd__a211o_1 _5690_ (.A1(\i_debug_uart_tx.data_to_send[3] ),
    .A2(_2336_),
    .B1(_2341_),
    .C1(_2347_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2348_));
 sky130_fd_sc_hd__o211a_1 _5691_ (.A1(\i_debug_uart_tx.uart_tx_data[3] ),
    .A2(_2330_),
    .B1(_2348_),
    .C1(_2299_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0176_));
 sky130_fd_sc_hd__and2_1 _5692_ (.A(\i_debug_uart_tx.data_to_send[5] ),
    .B(_2337_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2349_));
 sky130_fd_sc_hd__a211o_1 _5693_ (.A1(\i_debug_uart_tx.data_to_send[4] ),
    .A2(_2336_),
    .B1(_2341_),
    .C1(_2349_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2350_));
 sky130_fd_sc_hd__o211a_1 _5694_ (.A1(\i_debug_uart_tx.uart_tx_data[4] ),
    .A2(_2330_),
    .B1(_2350_),
    .C1(_2299_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0177_));
 sky130_fd_sc_hd__and2_1 _5695_ (.A(\i_debug_uart_tx.data_to_send[6] ),
    .B(_2337_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2351_));
 sky130_fd_sc_hd__a211o_1 _5696_ (.A1(\i_debug_uart_tx.data_to_send[5] ),
    .A2(_2336_),
    .B1(_2341_),
    .C1(_2351_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2352_));
 sky130_fd_sc_hd__o211a_1 _5697_ (.A1(\i_debug_uart_tx.uart_tx_data[5] ),
    .A2(_2330_),
    .B1(_2352_),
    .C1(_2299_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0178_));
 sky130_fd_sc_hd__and2_1 _5698_ (.A(\i_debug_uart_tx.data_to_send[7] ),
    .B(_2337_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2353_));
 sky130_fd_sc_hd__a211o_1 _5699_ (.A1(\i_debug_uart_tx.data_to_send[6] ),
    .A2(_2336_),
    .B1(_2341_),
    .C1(_2353_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2354_));
 sky130_fd_sc_hd__o211a_1 _5700_ (.A1(net319),
    .A2(_2330_),
    .B1(_2354_),
    .C1(_2299_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0179_));
 sky130_fd_sc_hd__a21o_1 _5701_ (.A1(net278),
    .A2(_2336_),
    .B1(_2341_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2355_));
 sky130_fd_sc_hd__o211a_1 _5702_ (.A1(\i_debug_uart_tx.uart_tx_data[7] ),
    .A2(_2330_),
    .B1(_2355_),
    .C1(_2299_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0180_));
 sky130_fd_sc_hd__nand2_1 _5703_ (.A(\i_debug_uart_tx.cycle_counter[0] ),
    .B(_0989_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2356_));
 sky130_fd_sc_hd__nor2_1 _5704_ (.A(_2198_),
    .B(_2333_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2357_));
 sky130_fd_sc_hd__o211a_1 _5705_ (.A1(\i_debug_uart_tx.cycle_counter[0] ),
    .A2(_0989_),
    .B1(_2356_),
    .C1(_2357_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0181_));
 sky130_fd_sc_hd__inv_2 _5706_ (.A(net188),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2358_));
 sky130_fd_sc_hd__o21ai_1 _5707_ (.A1(_2358_),
    .A2(_2356_),
    .B1(_2357_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2359_));
 sky130_fd_sc_hd__a21oi_1 _5708_ (.A1(_2358_),
    .A2(_2356_),
    .B1(_2359_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0182_));
 sky130_fd_sc_hd__and4_1 _5709_ (.A(\i_debug_uart_tx.cycle_counter[2] ),
    .B(\i_debug_uart_tx.cycle_counter[1] ),
    .C(\i_debug_uart_tx.cycle_counter[0] ),
    .D(_0989_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2360_));
 sky130_fd_sc_hd__a31o_1 _5710_ (.A1(\i_debug_uart_tx.cycle_counter[1] ),
    .A2(\i_debug_uart_tx.cycle_counter[0] ),
    .A3(_0989_),
    .B1(\i_debug_uart_tx.cycle_counter[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2361_));
 sky130_fd_sc_hd__and3b_1 _5711_ (.A_N(_2360_),
    .B(_2357_),
    .C(_2361_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2362_));
 sky130_fd_sc_hd__clkbuf_1 _5712_ (.A(_2362_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0183_));
 sky130_fd_sc_hd__or2_1 _5713_ (.A(\i_debug_uart_tx.cycle_counter[3] ),
    .B(_2360_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2363_));
 sky130_fd_sc_hd__nand2_1 _5714_ (.A(\i_debug_uart_tx.cycle_counter[3] ),
    .B(_2360_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2364_));
 sky130_fd_sc_hd__and3_1 _5715_ (.A(_2357_),
    .B(_2363_),
    .C(_2364_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2365_));
 sky130_fd_sc_hd__clkbuf_1 _5716_ (.A(_2365_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0184_));
 sky130_fd_sc_hd__and3_1 _5717_ (.A(\i_debug_uart_tx.cycle_counter[4] ),
    .B(_1729_),
    .C(_2364_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2366_));
 sky130_fd_sc_hd__clkbuf_1 _5718_ (.A(_2366_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0185_));
 sky130_fd_sc_hd__nand2_1 _5719_ (.A(\i_debug_uart_tx.fsm_state[3] ),
    .B(\i_debug_uart_tx.fsm_state[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2367_));
 sky130_fd_sc_hd__o21ba_1 _5720_ (.A1(\i_debug_uart_tx.fsm_state[2] ),
    .A2(_2367_),
    .B1_N(\i_debug_uart_tx.fsm_state[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2368_));
 sky130_fd_sc_hd__a21o_1 _5721_ (.A1(_0988_),
    .A2(_2368_),
    .B1(_2341_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2369_));
 sky130_fd_sc_hd__or2_1 _5722_ (.A(_2339_),
    .B(_2333_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2370_));
 sky130_fd_sc_hd__a32o_1 _5723_ (.A1(_2221_),
    .A2(_2369_),
    .A3(_2370_),
    .B1(_2357_),
    .B2(\i_debug_uart_tx.fsm_state[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0186_));
 sky130_fd_sc_hd__nor2_1 _5724_ (.A(_2339_),
    .B(_2333_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2371_));
 sky130_fd_sc_hd__or3b_1 _5725_ (.A(_2368_),
    .B(_2371_),
    .C_N(\i_debug_uart_tx.fsm_state[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2372_));
 sky130_fd_sc_hd__a21o_1 _5726_ (.A1(\i_debug_uart_tx.fsm_state[0] ),
    .A2(_2333_),
    .B1(\i_debug_uart_tx.fsm_state[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2373_));
 sky130_fd_sc_hd__and3_1 _5727_ (.A(_2181_),
    .B(_2372_),
    .C(_2373_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2374_));
 sky130_fd_sc_hd__clkbuf_1 _5728_ (.A(_2374_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0187_));
 sky130_fd_sc_hd__and4_1 _5729_ (.A(\i_debug_uart_tx.fsm_state[2] ),
    .B(\i_debug_uart_tx.fsm_state[1] ),
    .C(\i_debug_uart_tx.fsm_state[0] ),
    .D(_2333_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2375_));
 sky130_fd_sc_hd__a31o_1 _5730_ (.A1(\i_debug_uart_tx.fsm_state[1] ),
    .A2(\i_debug_uart_tx.fsm_state[0] ),
    .A3(_2333_),
    .B1(\i_debug_uart_tx.fsm_state[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2376_));
 sky130_fd_sc_hd__and3b_1 _5731_ (.A_N(_2375_),
    .B(_2376_),
    .C(_1729_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2377_));
 sky130_fd_sc_hd__clkbuf_1 _5732_ (.A(_2377_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0188_));
 sky130_fd_sc_hd__xor2_1 _5733_ (.A(\i_debug_uart_tx.fsm_state[2] ),
    .B(\i_debug_uart_tx.fsm_state[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2378_));
 sky130_fd_sc_hd__or2_1 _5734_ (.A(\i_debug_uart_tx.fsm_state[3] ),
    .B(_2375_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2379_));
 sky130_fd_sc_hd__o311a_1 _5735_ (.A1(_2367_),
    .A2(_2371_),
    .A3(_2378_),
    .B1(_2379_),
    .C1(_2221_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0189_));
 sky130_fd_sc_hd__nand2_1 _5736_ (.A(\i_spi.clock_divider[1] ),
    .B(\i_spi.clock_count[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2380_));
 sky130_fd_sc_hd__or2_1 _5737_ (.A(\i_spi.clock_divider[1] ),
    .B(\i_spi.clock_count[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2381_));
 sky130_fd_sc_hd__xor2_1 _5738_ (.A(\i_spi.clock_divider[0] ),
    .B(\i_spi.clock_count[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2382_));
 sky130_fd_sc_hd__a21oi_1 _5739_ (.A1(_2380_),
    .A2(_2381_),
    .B1(_2382_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2383_));
 sky130_fd_sc_hd__nand2_1 _5740_ (.A(\i_spi.busy ),
    .B(_2383_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2384_));
 sky130_fd_sc_hd__nand2_1 _5741_ (.A(\i_spi.busy ),
    .B(\i_spi.clock_count[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2385_));
 sky130_fd_sc_hd__clkbuf_4 _5742_ (.A(\i_spi.busy ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2386_));
 sky130_fd_sc_hd__or2_1 _5743_ (.A(_2386_),
    .B(\i_spi.clock_count[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2387_));
 sky130_fd_sc_hd__and4_1 _5744_ (.A(_1729_),
    .B(_2384_),
    .C(_2385_),
    .D(_2387_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2388_));
 sky130_fd_sc_hd__clkbuf_1 _5745_ (.A(_2388_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0190_));
 sky130_fd_sc_hd__xnor2_1 _5746_ (.A(\i_spi.clock_count[1] ),
    .B(_2385_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2389_));
 sky130_fd_sc_hd__and3_1 _5747_ (.A(_2181_),
    .B(_2384_),
    .C(_2389_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2390_));
 sky130_fd_sc_hd__clkbuf_1 _5748_ (.A(_2390_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0191_));
 sky130_fd_sc_hd__mux2_1 _5749_ (.A0(\i_debug_uart_tx.uart_tx_data[0] ),
    .A1(net4),
    .S(_2386_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2391_));
 sky130_fd_sc_hd__and2_1 _5750_ (.A(\i_spi.busy ),
    .B(_2383_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2392_));
 sky130_fd_sc_hd__and3b_1 _5751_ (.A_N(\i_spi.busy ),
    .B(_1000_),
    .C(_1557_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2393_));
 sky130_fd_sc_hd__clkbuf_2 _5752_ (.A(_2393_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2394_));
 sky130_fd_sc_hd__nor2_1 _5753_ (.A(_2392_),
    .B(_2394_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2395_));
 sky130_fd_sc_hd__or2_1 _5754_ (.A(_2198_),
    .B(_2395_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2396_));
 sky130_fd_sc_hd__nor2_1 _5755_ (.A(\i_spi.bits_remaining[3] ),
    .B(_2396_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2397_));
 sky130_fd_sc_hd__nor2_1 _5756_ (.A(\i_spi.spi_clk_out ),
    .B(_2384_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2398_));
 sky130_fd_sc_hd__nor2_4 _5757_ (.A(_2396_),
    .B(_2398_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2399_));
 sky130_fd_sc_hd__a21oi_1 _5758_ (.A1(\i_spi.read_latency ),
    .A2(_2397_),
    .B1(_2399_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2400_));
 sky130_fd_sc_hd__mux2_1 _5759_ (.A0(_2391_),
    .A1(\i_spi.data[0] ),
    .S(_2400_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2401_));
 sky130_fd_sc_hd__clkbuf_1 _5760_ (.A(_2401_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0192_));
 sky130_fd_sc_hd__or2_1 _5761_ (.A(\i_spi.bits_remaining[1] ),
    .B(\i_spi.bits_remaining[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2402_));
 sky130_fd_sc_hd__or3_1 _5762_ (.A(\i_spi.bits_remaining[3] ),
    .B(\i_spi.bits_remaining[2] ),
    .C(_2402_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2403_));
 sky130_fd_sc_hd__and3_2 _5763_ (.A(\i_spi.spi_clk_out ),
    .B(_2392_),
    .C(_2403_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2404_));
 sky130_fd_sc_hd__o21ai_1 _5764_ (.A1(_2394_),
    .A2(_2404_),
    .B1(net239),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2405_));
 sky130_fd_sc_hd__o211a_1 _5765_ (.A1(net239),
    .A2(_2404_),
    .B1(_2405_),
    .C1(_2299_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0193_));
 sky130_fd_sc_hd__nor2_1 _5766_ (.A(_2394_),
    .B(_2404_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2406_));
 sky130_fd_sc_hd__nand2_1 _5767_ (.A(\i_spi.bits_remaining[1] ),
    .B(\i_spi.bits_remaining[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2407_));
 sky130_fd_sc_hd__nand2_1 _5768_ (.A(_2402_),
    .B(_2407_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2408_));
 sky130_fd_sc_hd__a22o_1 _5769_ (.A1(\i_spi.bits_remaining[1] ),
    .A2(_2406_),
    .B1(_2408_),
    .B2(_2404_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2409_));
 sky130_fd_sc_hd__and2_1 _5770_ (.A(_2221_),
    .B(_2409_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2410_));
 sky130_fd_sc_hd__clkbuf_1 _5771_ (.A(_2410_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0194_));
 sky130_fd_sc_hd__xnor2_1 _5772_ (.A(\i_spi.bits_remaining[2] ),
    .B(_2402_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2411_));
 sky130_fd_sc_hd__a22o_1 _5773_ (.A1(\i_spi.bits_remaining[2] ),
    .A2(_2406_),
    .B1(_2411_),
    .B2(_2404_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2412_));
 sky130_fd_sc_hd__and2_1 _5774_ (.A(_2181_),
    .B(_2412_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2413_));
 sky130_fd_sc_hd__clkbuf_1 _5775_ (.A(_2413_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0195_));
 sky130_fd_sc_hd__or3b_1 _5776_ (.A(\i_spi.bits_remaining[2] ),
    .B(_2402_),
    .C_N(_2404_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2414_));
 sky130_fd_sc_hd__nand2_2 _5777_ (.A(_1728_),
    .B(_2394_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2415_));
 sky130_fd_sc_hd__inv_2 _5778_ (.A(_2415_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2416_));
 sky130_fd_sc_hd__a31o_1 _5779_ (.A1(net194),
    .A2(_2221_),
    .A3(_2414_),
    .B1(_2416_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0196_));
 sky130_fd_sc_hd__a21o_1 _5780_ (.A1(_1000_),
    .A2(_1725_),
    .B1(_2386_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2417_));
 sky130_fd_sc_hd__or3_1 _5781_ (.A(\i_spi.spi_clk_out ),
    .B(_2384_),
    .C(_2403_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2418_));
 sky130_fd_sc_hd__and3_1 _5782_ (.A(_2181_),
    .B(_2417_),
    .C(_2418_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2419_));
 sky130_fd_sc_hd__clkbuf_1 _5783_ (.A(_2419_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0197_));
 sky130_fd_sc_hd__mux2_1 _5784_ (.A0(\i_spi.dc_in ),
    .A1(net282),
    .S(_2415_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2420_));
 sky130_fd_sc_hd__clkbuf_1 _5785_ (.A(_2420_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0198_));
 sky130_fd_sc_hd__inv_2 _5786_ (.A(net184),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2421_));
 sky130_fd_sc_hd__nand2_1 _5787_ (.A(\i_spi.spi_select ),
    .B(_2418_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2422_));
 sky130_fd_sc_hd__o221ai_1 _5788_ (.A1(_2421_),
    .A2(_2418_),
    .B1(_2422_),
    .B2(_2394_),
    .C1(_2221_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0199_));
 sky130_fd_sc_hd__a22o_1 _5789_ (.A1(\i_spi.spi_clk_out ),
    .A2(_2395_),
    .B1(_2398_),
    .B2(_2403_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2423_));
 sky130_fd_sc_hd__and2_1 _5790_ (.A(_2181_),
    .B(_2423_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2424_));
 sky130_fd_sc_hd__clkbuf_1 _5791_ (.A(_2424_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0200_));
 sky130_fd_sc_hd__o21a_1 _5792_ (.A1(net205),
    .A2(_2334_),
    .B1(_0988_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2425_));
 sky130_fd_sc_hd__or3_1 _5793_ (.A(_2198_),
    .B(_2339_),
    .C(_2425_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2426_));
 sky130_fd_sc_hd__clkbuf_1 _5794_ (.A(_2426_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0201_));
 sky130_fd_sc_hd__nand2_1 _5795_ (.A(_1004_),
    .B(_1725_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2427_));
 sky130_fd_sc_hd__a21o_1 _5796_ (.A1(_1004_),
    .A2(_1725_),
    .B1(net220),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2428_));
 sky130_fd_sc_hd__o211a_1 _5797_ (.A1(net98),
    .A2(_2427_),
    .B1(_2428_),
    .C1(_2221_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0202_));
 sky130_fd_sc_hd__a31o_1 _5798_ (.A1(\i_debug_uart_tx.uart_tx_data[0] ),
    .A2(_1004_),
    .A3(_1725_),
    .B1(_2229_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2429_));
 sky130_fd_sc_hd__a21o_1 _5799_ (.A1(net162),
    .A2(_2427_),
    .B1(_2429_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0203_));
 sky130_fd_sc_hd__a21o_1 _5800_ (.A1(_1004_),
    .A2(_1725_),
    .B1(net204),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2430_));
 sky130_fd_sc_hd__o211a_1 _5801_ (.A1(net97),
    .A2(_2427_),
    .B1(_2430_),
    .C1(_2221_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0204_));
 sky130_fd_sc_hd__inv_2 _5802_ (.A(net192),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2431_));
 sky130_fd_sc_hd__inv_2 _5803_ (.A(_0942_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2432_));
 sky130_fd_sc_hd__a41o_1 _5804_ (.A1(_0920_),
    .A2(_0936_),
    .A3(_0932_),
    .A4(_2432_),
    .B1(_0974_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2433_));
 sky130_fd_sc_hd__nand2_2 _5805_ (.A(_0920_),
    .B(_0944_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2434_));
 sky130_fd_sc_hd__or4bb_1 _5806_ (.A(_0752_),
    .B(_0907_),
    .C_N(_2433_),
    .D_N(_2434_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2435_));
 sky130_fd_sc_hd__a31o_1 _5807_ (.A1(_0613_),
    .A2(net66),
    .A3(_2088_),
    .B1(_2435_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2436_));
 sky130_fd_sc_hd__o21ai_1 _5808_ (.A1(net66),
    .A2(_2102_),
    .B1(_0613_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2437_));
 sky130_fd_sc_hd__inv_2 _5809_ (.A(\i_tinyqv.cpu.i_core.last_interrupt_req[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2438_));
 sky130_fd_sc_hd__a211o_1 _5810_ (.A1(\i_tinyqv.cpu.i_core.interrupt_req[1] ),
    .A2(_2438_),
    .B1(_0613_),
    .C1(\i_tinyqv.cpu.i_core.mip[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2439_));
 sky130_fd_sc_hd__a21oi_1 _5811_ (.A1(_2437_),
    .A2(_2439_),
    .B1(_2436_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2440_));
 sky130_fd_sc_hd__a211oi_1 _5812_ (.A1(_2431_),
    .A2(_2436_),
    .B1(_2440_),
    .C1(_2083_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0205_));
 sky130_fd_sc_hd__a31o_1 _5813_ (.A1(_0613_),
    .A2(_1312_),
    .A3(_2088_),
    .B1(_2435_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2441_));
 sky130_fd_sc_hd__nor2_1 _5814_ (.A(_1312_),
    .B(_2102_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2442_));
 sky130_fd_sc_hd__or2b_1 _5815_ (.A(\i_tinyqv.cpu.i_core.last_interrupt_req[0] ),
    .B_N(\i_tinyqv.cpu.i_core.interrupt_req[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2443_));
 sky130_fd_sc_hd__a21oi_1 _5816_ (.A1(_0916_),
    .A2(_2443_),
    .B1(_2441_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2444_));
 sky130_fd_sc_hd__o32a_1 _5817_ (.A1(_0916_),
    .A2(_2441_),
    .A3(_2442_),
    .B1(_2444_),
    .B2(\i_tinyqv.cpu.i_core.mip[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2445_));
 sky130_fd_sc_hd__and2b_1 _5818_ (.A_N(_2083_),
    .B(_2445_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2446_));
 sky130_fd_sc_hd__clkbuf_1 _5819_ (.A(_2446_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0206_));
 sky130_fd_sc_hd__and2b_1 _5820_ (.A_N(net42),
    .B(_2088_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2447_));
 sky130_fd_sc_hd__o21ai_1 _5821_ (.A1(_2434_),
    .A2(_2447_),
    .B1(net200),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2448_));
 sky130_fd_sc_hd__nand2_1 _5822_ (.A(_0944_),
    .B(_2103_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2449_));
 sky130_fd_sc_hd__a21oi_1 _5823_ (.A1(_2448_),
    .A2(_2449_),
    .B1(_2083_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0207_));
 sky130_fd_sc_hd__a21o_1 _5824_ (.A1(net81),
    .A2(_2088_),
    .B1(_2434_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2450_));
 sky130_fd_sc_hd__nand2_1 _5825_ (.A(net179),
    .B(_2450_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2451_));
 sky130_fd_sc_hd__a211o_1 _5826_ (.A1(net69),
    .A2(_2088_),
    .B1(_2434_),
    .C1(net81),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2452_));
 sky130_fd_sc_hd__a21oi_1 _5827_ (.A1(_2451_),
    .A2(_2452_),
    .B1(_2083_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0208_));
 sky130_fd_sc_hd__a21o_1 _5828_ (.A1(net66),
    .A2(_2088_),
    .B1(_2434_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2453_));
 sky130_fd_sc_hd__nand2_1 _5829_ (.A(net182),
    .B(_2453_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2454_));
 sky130_fd_sc_hd__or3b_1 _5830_ (.A(_2102_),
    .B(net67),
    .C_N(_0944_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2455_));
 sky130_fd_sc_hd__a21oi_1 _5831_ (.A1(_2454_),
    .A2(_2455_),
    .B1(_2083_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0209_));
 sky130_fd_sc_hd__a21o_1 _5832_ (.A1(_1312_),
    .A2(_2088_),
    .B1(_2434_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2456_));
 sky130_fd_sc_hd__a22oi_1 _5833_ (.A1(_0944_),
    .A2(_2442_),
    .B1(_2456_),
    .B2(net230),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2457_));
 sky130_fd_sc_hd__nor2_1 _5834_ (.A(_2083_),
    .B(_2457_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0210_));
 sky130_fd_sc_hd__nand2_1 _5835_ (.A(_2221_),
    .B(_2170_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2458_));
 sky130_fd_sc_hd__a211o_1 _5836_ (.A1(net116),
    .A2(_0990_),
    .B1(_0991_),
    .C1(_2458_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0211_));
 sky130_fd_sc_hd__inv_2 _5837__1 (.A(clknet_leaf_18_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net29));
 sky130_fd_sc_hd__or2_1 _5838_ (.A(_2066_),
    .B(\i_tinyqv.cpu.instr_data[1][0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2459_));
 sky130_fd_sc_hd__nand2_1 _5839_ (.A(\i_tinyqv.cpu.i_core.i_cycles.rstn ),
    .B(_2307_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2460_));
 sky130_fd_sc_hd__or3b_1 _5840_ (.A(_2460_),
    .B(\i_tinyqv.cpu.instr_write_offset[2] ),
    .C_N(_1406_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2461_));
 sky130_fd_sc_hd__clkbuf_4 _5841_ (.A(_2461_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2462_));
 sky130_fd_sc_hd__buf_4 _5842_ (.A(_2462_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2463_));
 sky130_fd_sc_hd__mux2_1 _5843_ (.A0(\i_tinyqv.cpu.instr_data_in[0] ),
    .A1(_2459_),
    .S(_2463_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2464_));
 sky130_fd_sc_hd__clkbuf_1 _5844_ (.A(_2464_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0212_));
 sky130_fd_sc_hd__or2_1 _5845_ (.A(_1400_),
    .B(\i_tinyqv.cpu.instr_data[1][1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2465_));
 sky130_fd_sc_hd__mux2_1 _5846_ (.A0(\i_tinyqv.cpu.instr_data_in[1] ),
    .A1(_2465_),
    .S(_2463_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2466_));
 sky130_fd_sc_hd__clkbuf_1 _5847_ (.A(_2466_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0213_));
 sky130_fd_sc_hd__or3_1 _5848_ (.A(\i_tinyqv.cpu.instr_write_offset[2] ),
    .B(_1406_),
    .C(_2460_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2467_));
 sky130_fd_sc_hd__clkbuf_4 _5849_ (.A(_2467_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2468_));
 sky130_fd_sc_hd__buf_4 _5850_ (.A(_2468_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2469_));
 sky130_fd_sc_hd__mux2_1 _5851_ (.A0(\i_tinyqv.cpu.instr_data_in[2] ),
    .A1(\i_tinyqv.cpu.instr_data[0][2] ),
    .S(_2469_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2470_));
 sky130_fd_sc_hd__clkbuf_1 _5852_ (.A(_2470_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0214_));
 sky130_fd_sc_hd__mux2_1 _5853_ (.A0(\i_tinyqv.cpu.instr_data_in[3] ),
    .A1(net291),
    .S(_2469_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2471_));
 sky130_fd_sc_hd__clkbuf_1 _5854_ (.A(_2471_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0215_));
 sky130_fd_sc_hd__mux2_1 _5855_ (.A0(\i_tinyqv.cpu.instr_data_in[4] ),
    .A1(\i_tinyqv.cpu.instr_data[0][4] ),
    .S(_2469_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2472_));
 sky130_fd_sc_hd__clkbuf_1 _5856_ (.A(_2472_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0216_));
 sky130_fd_sc_hd__mux2_1 _5857_ (.A0(\i_tinyqv.cpu.instr_data_in[5] ),
    .A1(\i_tinyqv.cpu.instr_data[0][5] ),
    .S(_2469_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2473_));
 sky130_fd_sc_hd__clkbuf_1 _5858_ (.A(_2473_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0217_));
 sky130_fd_sc_hd__mux2_1 _5859_ (.A0(\i_tinyqv.cpu.instr_data_in[6] ),
    .A1(\i_tinyqv.cpu.instr_data[0][6] ),
    .S(_2469_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2474_));
 sky130_fd_sc_hd__clkbuf_1 _5860_ (.A(_2474_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0218_));
 sky130_fd_sc_hd__mux2_1 _5861_ (.A0(\i_tinyqv.cpu.instr_data_in[7] ),
    .A1(\i_tinyqv.cpu.instr_data[0][7] ),
    .S(_2469_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2475_));
 sky130_fd_sc_hd__clkbuf_1 _5862_ (.A(_2475_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0219_));
 sky130_fd_sc_hd__mux2_1 _5863_ (.A0(_2316_),
    .A1(\i_tinyqv.cpu.instr_data[0][8] ),
    .S(_2469_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2476_));
 sky130_fd_sc_hd__clkbuf_1 _5864_ (.A(_2476_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0220_));
 sky130_fd_sc_hd__mux2_1 _5865_ (.A0(_2318_),
    .A1(\i_tinyqv.cpu.instr_data[0][9] ),
    .S(_2469_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2477_));
 sky130_fd_sc_hd__clkbuf_1 _5866_ (.A(_2477_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0221_));
 sky130_fd_sc_hd__mux2_1 _5867_ (.A0(_2320_),
    .A1(\i_tinyqv.cpu.instr_data[0][10] ),
    .S(_2469_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2478_));
 sky130_fd_sc_hd__clkbuf_1 _5868_ (.A(_2478_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0222_));
 sky130_fd_sc_hd__mux2_1 _5869_ (.A0(_2322_),
    .A1(\i_tinyqv.cpu.instr_data[0][11] ),
    .S(_2469_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2479_));
 sky130_fd_sc_hd__clkbuf_1 _5870_ (.A(_2479_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0223_));
 sky130_fd_sc_hd__mux2_1 _5871_ (.A0(_1712_),
    .A1(\i_tinyqv.cpu.instr_data[0][12] ),
    .S(_2468_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2480_));
 sky130_fd_sc_hd__clkbuf_1 _5872_ (.A(_2480_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0224_));
 sky130_fd_sc_hd__mux2_1 _5873_ (.A0(_1717_),
    .A1(\i_tinyqv.cpu.instr_data[0][13] ),
    .S(_2468_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2481_));
 sky130_fd_sc_hd__clkbuf_1 _5874_ (.A(_2481_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0225_));
 sky130_fd_sc_hd__mux2_1 _5875_ (.A0(_1720_),
    .A1(net266),
    .S(_2468_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2482_));
 sky130_fd_sc_hd__clkbuf_1 _5876_ (.A(_2482_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0226_));
 sky130_fd_sc_hd__mux2_1 _5877_ (.A0(_1721_),
    .A1(net283),
    .S(_2468_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2483_));
 sky130_fd_sc_hd__clkbuf_1 _5878_ (.A(_2483_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0227_));
 sky130_fd_sc_hd__inv_2 _5879_ (.A(_2309_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2484_));
 sky130_fd_sc_hd__a31o_1 _5880_ (.A1(\i_tinyqv.cpu.instr_write_offset[2] ),
    .A2(_1406_),
    .A3(_2307_),
    .B1(_2066_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2485_));
 sky130_fd_sc_hd__o22a_1 _5881_ (.A1(\i_tinyqv.cpu.instr_data_in[0] ),
    .A2(_2484_),
    .B1(_2485_),
    .B2(net100),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0228_));
 sky130_fd_sc_hd__o22a_1 _5882_ (.A1(\i_tinyqv.cpu.instr_data_in[1] ),
    .A2(_2484_),
    .B1(_2485_),
    .B2(net106),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0229_));
 sky130_fd_sc_hd__mux2_1 _5883_ (.A0(\i_debug_uart_tx.uart_tx_data[1] ),
    .A1(\i_spi.data[0] ),
    .S(_2386_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2486_));
 sky130_fd_sc_hd__mux2_1 _5884_ (.A0(\i_spi.data[1] ),
    .A1(_2486_),
    .S(_2399_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2487_));
 sky130_fd_sc_hd__clkbuf_1 _5885_ (.A(_2487_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0230_));
 sky130_fd_sc_hd__mux2_1 _5886_ (.A0(\i_debug_uart_tx.uart_tx_data[2] ),
    .A1(\i_spi.data[1] ),
    .S(_2386_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2488_));
 sky130_fd_sc_hd__mux2_1 _5887_ (.A0(\i_spi.data[2] ),
    .A1(_2488_),
    .S(_2399_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2489_));
 sky130_fd_sc_hd__clkbuf_1 _5888_ (.A(_2489_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0231_));
 sky130_fd_sc_hd__mux2_1 _5889_ (.A0(\i_debug_uart_tx.uart_tx_data[3] ),
    .A1(\i_spi.data[2] ),
    .S(_2386_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2490_));
 sky130_fd_sc_hd__mux2_1 _5890_ (.A0(\i_spi.data[3] ),
    .A1(_2490_),
    .S(_2399_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2491_));
 sky130_fd_sc_hd__clkbuf_1 _5891_ (.A(_2491_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0232_));
 sky130_fd_sc_hd__mux2_1 _5892_ (.A0(\i_debug_uart_tx.uart_tx_data[4] ),
    .A1(\i_spi.data[3] ),
    .S(_2386_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2492_));
 sky130_fd_sc_hd__mux2_1 _5893_ (.A0(\i_spi.data[4] ),
    .A1(_2492_),
    .S(_2399_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2493_));
 sky130_fd_sc_hd__clkbuf_1 _5894_ (.A(_2493_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0233_));
 sky130_fd_sc_hd__mux2_1 _5895_ (.A0(\i_debug_uart_tx.uart_tx_data[5] ),
    .A1(\i_spi.data[4] ),
    .S(_2386_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2494_));
 sky130_fd_sc_hd__mux2_1 _5896_ (.A0(\i_spi.data[5] ),
    .A1(_2494_),
    .S(_2399_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2495_));
 sky130_fd_sc_hd__clkbuf_1 _5897_ (.A(_2495_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0234_));
 sky130_fd_sc_hd__mux2_1 _5898_ (.A0(\i_debug_uart_tx.uart_tx_data[6] ),
    .A1(\i_spi.data[5] ),
    .S(_2386_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2496_));
 sky130_fd_sc_hd__mux2_1 _5899_ (.A0(\i_spi.data[6] ),
    .A1(_2496_),
    .S(_2399_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2497_));
 sky130_fd_sc_hd__clkbuf_1 _5900_ (.A(_2497_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0235_));
 sky130_fd_sc_hd__mux2_1 _5901_ (.A0(\i_debug_uart_tx.uart_tx_data[7] ),
    .A1(\i_spi.data[6] ),
    .S(_2386_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2498_));
 sky130_fd_sc_hd__mux2_1 _5902_ (.A0(\i_spi.data[7] ),
    .A1(_2498_),
    .S(_2399_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2499_));
 sky130_fd_sc_hd__clkbuf_1 _5903_ (.A(_2499_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0236_));
 sky130_fd_sc_hd__mux2_1 _5904_ (.A0(\i_tinyqv.cpu.i_core.mepc[0] ),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[4] ),
    .S(_1393_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2500_));
 sky130_fd_sc_hd__nor2_4 _5905_ (.A(_1400_),
    .B(_1758_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2501_));
 sky130_fd_sc_hd__buf_4 _5906_ (.A(_2501_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2502_));
 sky130_fd_sc_hd__mux2_1 _5907_ (.A0(\i_tinyqv.cpu.data_addr[0] ),
    .A1(_2500_),
    .S(_2502_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2503_));
 sky130_fd_sc_hd__clkbuf_1 _5908_ (.A(_2503_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0237_));
 sky130_fd_sc_hd__clkbuf_4 _5909_ (.A(_2106_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2504_));
 sky130_fd_sc_hd__mux2_2 _5910_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[5] ),
    .A1(\i_tinyqv.cpu.i_core.mepc[1] ),
    .S(_2504_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2505_));
 sky130_fd_sc_hd__mux2_1 _5911_ (.A0(net137),
    .A1(_2505_),
    .S(_2502_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2506_));
 sky130_fd_sc_hd__clkbuf_1 _5912_ (.A(_2506_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0238_));
 sky130_fd_sc_hd__mux2_2 _5913_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[6] ),
    .A1(\i_tinyqv.cpu.i_core.mepc[2] ),
    .S(_2504_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2507_));
 sky130_fd_sc_hd__mux2_1 _5914_ (.A0(\i_tinyqv.cpu.data_addr[2] ),
    .A1(_2507_),
    .S(_2502_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2508_));
 sky130_fd_sc_hd__clkbuf_1 _5915_ (.A(_2508_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0239_));
 sky130_fd_sc_hd__mux2_1 _5916_ (.A0(_1054_),
    .A1(\i_tinyqv.cpu.i_core.mepc[3] ),
    .S(_2106_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2509_));
 sky130_fd_sc_hd__mux2_1 _5917_ (.A0(\i_tinyqv.cpu.data_addr[3] ),
    .A1(_2509_),
    .S(_2502_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2510_));
 sky130_fd_sc_hd__clkbuf_1 _5918_ (.A(_2510_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0240_));
 sky130_fd_sc_hd__mux2_1 _5919_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[8] ),
    .A1(\i_tinyqv.cpu.i_core.mepc[4] ),
    .S(_2504_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2511_));
 sky130_fd_sc_hd__mux2_1 _5920_ (.A0(\i_tinyqv.cpu.data_addr[4] ),
    .A1(_2511_),
    .S(_2502_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2512_));
 sky130_fd_sc_hd__clkbuf_1 _5921_ (.A(_2512_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0241_));
 sky130_fd_sc_hd__mux2_2 _5922_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[9] ),
    .A1(\i_tinyqv.cpu.i_core.mepc[5] ),
    .S(_2107_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2513_));
 sky130_fd_sc_hd__mux2_1 _5923_ (.A0(\i_tinyqv.cpu.data_addr[5] ),
    .A1(_2513_),
    .S(_2502_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2514_));
 sky130_fd_sc_hd__clkbuf_1 _5924_ (.A(_2514_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0242_));
 sky130_fd_sc_hd__mux2_1 _5925_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[10] ),
    .A1(\i_tinyqv.cpu.i_core.mepc[6] ),
    .S(_2504_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2515_));
 sky130_fd_sc_hd__mux2_1 _5926_ (.A0(\i_tinyqv.cpu.data_addr[6] ),
    .A1(_2515_),
    .S(_2502_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2516_));
 sky130_fd_sc_hd__clkbuf_1 _5927_ (.A(_2516_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0243_));
 sky130_fd_sc_hd__mux2_1 _5928_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[11] ),
    .A1(\i_tinyqv.cpu.i_core.mepc[7] ),
    .S(_2107_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2517_));
 sky130_fd_sc_hd__mux2_1 _5929_ (.A0(\i_tinyqv.cpu.data_addr[7] ),
    .A1(_2517_),
    .S(_2502_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2518_));
 sky130_fd_sc_hd__clkbuf_1 _5930_ (.A(_2518_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0244_));
 sky130_fd_sc_hd__mux2_1 _5931_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[12] ),
    .A1(\i_tinyqv.cpu.i_core.mepc[8] ),
    .S(_2106_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2519_));
 sky130_fd_sc_hd__mux2_1 _5932_ (.A0(\i_tinyqv.cpu.data_addr[8] ),
    .A1(_2519_),
    .S(_2502_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2520_));
 sky130_fd_sc_hd__clkbuf_1 _5933_ (.A(_2520_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0245_));
 sky130_fd_sc_hd__mux2_1 _5934_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[13] ),
    .A1(\i_tinyqv.cpu.i_core.mepc[9] ),
    .S(_2106_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2521_));
 sky130_fd_sc_hd__mux2_1 _5935_ (.A0(\i_tinyqv.cpu.data_addr[9] ),
    .A1(_2521_),
    .S(_2502_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2522_));
 sky130_fd_sc_hd__clkbuf_1 _5936_ (.A(_2522_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0246_));
 sky130_fd_sc_hd__mux2_1 _5937_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[14] ),
    .A1(\i_tinyqv.cpu.i_core.mepc[10] ),
    .S(_2504_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2523_));
 sky130_fd_sc_hd__clkbuf_4 _5938_ (.A(_2501_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2524_));
 sky130_fd_sc_hd__mux2_1 _5939_ (.A0(\i_tinyqv.cpu.data_addr[10] ),
    .A1(_2523_),
    .S(_2524_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2525_));
 sky130_fd_sc_hd__clkbuf_1 _5940_ (.A(_2525_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0247_));
 sky130_fd_sc_hd__mux2_1 _5941_ (.A0(_1060_),
    .A1(\i_tinyqv.cpu.i_core.mepc[11] ),
    .S(_2106_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2526_));
 sky130_fd_sc_hd__mux2_1 _5942_ (.A0(net314),
    .A1(_2526_),
    .S(_2524_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2527_));
 sky130_fd_sc_hd__clkbuf_1 _5943_ (.A(_2527_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0248_));
 sky130_fd_sc_hd__mux2_1 _5944_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[16] ),
    .A1(\i_tinyqv.cpu.i_core.mepc[12] ),
    .S(_2504_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2528_));
 sky130_fd_sc_hd__mux2_1 _5945_ (.A0(\i_tinyqv.cpu.data_addr[12] ),
    .A1(_2528_),
    .S(_2524_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2529_));
 sky130_fd_sc_hd__clkbuf_1 _5946_ (.A(_2529_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0249_));
 sky130_fd_sc_hd__mux2_1 _5947_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[17] ),
    .A1(\i_tinyqv.cpu.i_core.mepc[13] ),
    .S(_2106_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2530_));
 sky130_fd_sc_hd__mux2_1 _5948_ (.A0(\i_tinyqv.cpu.data_addr[13] ),
    .A1(_2530_),
    .S(_2524_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2531_));
 sky130_fd_sc_hd__clkbuf_1 _5949_ (.A(_2531_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0250_));
 sky130_fd_sc_hd__mux2_1 _5950_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[18] ),
    .A1(\i_tinyqv.cpu.i_core.mepc[14] ),
    .S(_2107_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2532_));
 sky130_fd_sc_hd__mux2_1 _5951_ (.A0(net111),
    .A1(_2532_),
    .S(_2524_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2533_));
 sky130_fd_sc_hd__clkbuf_1 _5952_ (.A(_2533_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0251_));
 sky130_fd_sc_hd__mux2_1 _5953_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[19] ),
    .A1(\i_tinyqv.cpu.i_core.mepc[15] ),
    .S(_2107_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2534_));
 sky130_fd_sc_hd__mux2_1 _5954_ (.A0(\i_tinyqv.cpu.data_addr[15] ),
    .A1(_2534_),
    .S(_2524_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2535_));
 sky130_fd_sc_hd__clkbuf_1 _5955_ (.A(_2535_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0252_));
 sky130_fd_sc_hd__mux2_1 _5956_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[20] ),
    .A1(\i_tinyqv.cpu.i_core.mepc[16] ),
    .S(_2504_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2536_));
 sky130_fd_sc_hd__mux2_1 _5957_ (.A0(\i_tinyqv.cpu.data_addr[16] ),
    .A1(_2536_),
    .S(_2524_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2537_));
 sky130_fd_sc_hd__clkbuf_1 _5958_ (.A(_2537_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0253_));
 sky130_fd_sc_hd__mux2_1 _5959_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[21] ),
    .A1(\i_tinyqv.cpu.i_core.mepc[17] ),
    .S(_2504_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2538_));
 sky130_fd_sc_hd__mux2_1 _5960_ (.A0(\i_tinyqv.cpu.data_addr[17] ),
    .A1(_2538_),
    .S(_2524_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2539_));
 sky130_fd_sc_hd__clkbuf_1 _5961_ (.A(_2539_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0254_));
 sky130_fd_sc_hd__mux2_1 _5962_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[22] ),
    .A1(\i_tinyqv.cpu.i_core.mepc[18] ),
    .S(_2504_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2540_));
 sky130_fd_sc_hd__mux2_1 _5963_ (.A0(\i_tinyqv.cpu.data_addr[18] ),
    .A1(_2540_),
    .S(_2524_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2541_));
 sky130_fd_sc_hd__clkbuf_1 _5964_ (.A(_2541_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0255_));
 sky130_fd_sc_hd__mux2_1 _5965_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[23] ),
    .A1(\i_tinyqv.cpu.i_core.mepc[19] ),
    .S(_2107_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2542_));
 sky130_fd_sc_hd__mux2_1 _5966_ (.A0(\i_tinyqv.cpu.data_addr[19] ),
    .A1(_2542_),
    .S(_2524_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2543_));
 sky130_fd_sc_hd__clkbuf_1 _5967_ (.A(_2543_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0256_));
 sky130_fd_sc_hd__mux2_1 _5968_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[24] ),
    .A1(\i_tinyqv.cpu.i_core.mepc[20] ),
    .S(_2106_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2544_));
 sky130_fd_sc_hd__mux2_1 _5969_ (.A0(\i_tinyqv.cpu.data_addr[20] ),
    .A1(_2544_),
    .S(_2501_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2545_));
 sky130_fd_sc_hd__clkbuf_1 _5970_ (.A(_2545_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0257_));
 sky130_fd_sc_hd__mux2_1 _5971_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[25] ),
    .A1(\i_tinyqv.cpu.i_core.mepc[21] ),
    .S(_2107_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2546_));
 sky130_fd_sc_hd__mux2_1 _5972_ (.A0(\i_tinyqv.cpu.data_addr[21] ),
    .A1(_2546_),
    .S(_2501_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2547_));
 sky130_fd_sc_hd__clkbuf_1 _5973_ (.A(_2547_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0258_));
 sky130_fd_sc_hd__mux2_1 _5974_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[26] ),
    .A1(\i_tinyqv.cpu.i_core.mepc[22] ),
    .S(_2106_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2548_));
 sky130_fd_sc_hd__mux2_1 _5975_ (.A0(\i_tinyqv.cpu.data_addr[22] ),
    .A1(_2548_),
    .S(_2501_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2549_));
 sky130_fd_sc_hd__clkbuf_1 _5976_ (.A(_2549_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0259_));
 sky130_fd_sc_hd__mux2_1 _5977_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[27] ),
    .A1(\i_tinyqv.cpu.i_core.mepc[23] ),
    .S(_2504_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2550_));
 sky130_fd_sc_hd__mux2_1 _5978_ (.A0(\i_tinyqv.cpu.data_addr[23] ),
    .A1(_2550_),
    .S(_2501_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2551_));
 sky130_fd_sc_hd__clkbuf_1 _5979_ (.A(_2551_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0260_));
 sky130_fd_sc_hd__nor2_1 _5980_ (.A(_2107_),
    .B(_1758_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2552_));
 sky130_fd_sc_hd__a22o_1 _5981_ (.A1(\i_tinyqv.cpu.data_addr[24] ),
    .A2(_1758_),
    .B1(_2552_),
    .B2(\i_tinyqv.cpu.i_core.i_shift.a[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2553_));
 sky130_fd_sc_hd__and2_1 _5982_ (.A(_2079_),
    .B(_2553_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2554_));
 sky130_fd_sc_hd__clkbuf_1 _5983_ (.A(_2554_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0261_));
 sky130_fd_sc_hd__a22o_1 _5984_ (.A1(\i_tinyqv.cpu.data_addr[25] ),
    .A2(_1758_),
    .B1(_2552_),
    .B2(\i_tinyqv.cpu.i_core.i_shift.a[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2555_));
 sky130_fd_sc_hd__and2_1 _5985_ (.A(_2079_),
    .B(_2555_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2556_));
 sky130_fd_sc_hd__clkbuf_1 _5986_ (.A(_2556_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0262_));
 sky130_fd_sc_hd__a22o_1 _5987_ (.A1(\i_tinyqv.cpu.data_addr[26] ),
    .A2(_1758_),
    .B1(_2552_),
    .B2(\i_tinyqv.cpu.i_core.i_shift.a[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2557_));
 sky130_fd_sc_hd__and2_1 _5988_ (.A(_2079_),
    .B(_2557_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2558_));
 sky130_fd_sc_hd__clkbuf_1 _5989_ (.A(_2558_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0263_));
 sky130_fd_sc_hd__a22o_1 _5990_ (.A1(\i_tinyqv.cpu.data_addr[27] ),
    .A2(_1758_),
    .B1(_2552_),
    .B2(\i_tinyqv.cpu.i_core.i_shift.a[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2559_));
 sky130_fd_sc_hd__and2_1 _5991_ (.A(_2079_),
    .B(_2559_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2560_));
 sky130_fd_sc_hd__clkbuf_1 _5992_ (.A(_2560_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0264_));
 sky130_fd_sc_hd__or3b_1 _5993_ (.A(_1406_),
    .B(_2460_),
    .C_N(\i_tinyqv.cpu.instr_write_offset[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2561_));
 sky130_fd_sc_hd__clkbuf_4 _5994_ (.A(_2561_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2562_));
 sky130_fd_sc_hd__buf_4 _5995_ (.A(_2562_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2563_));
 sky130_fd_sc_hd__mux2_1 _5996_ (.A0(\i_tinyqv.cpu.instr_data_in[2] ),
    .A1(\i_tinyqv.cpu.instr_data[2][2] ),
    .S(_2563_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2564_));
 sky130_fd_sc_hd__clkbuf_1 _5997_ (.A(_2564_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0265_));
 sky130_fd_sc_hd__mux2_1 _5998_ (.A0(\i_tinyqv.cpu.instr_data_in[3] ),
    .A1(\i_tinyqv.cpu.instr_data[2][3] ),
    .S(_2563_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2565_));
 sky130_fd_sc_hd__clkbuf_1 _5999_ (.A(_2565_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0266_));
 sky130_fd_sc_hd__mux2_1 _6000_ (.A0(\i_tinyqv.cpu.instr_data_in[4] ),
    .A1(\i_tinyqv.cpu.instr_data[2][4] ),
    .S(_2563_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2566_));
 sky130_fd_sc_hd__clkbuf_1 _6001_ (.A(_2566_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0267_));
 sky130_fd_sc_hd__mux2_1 _6002_ (.A0(\i_tinyqv.cpu.instr_data_in[5] ),
    .A1(\i_tinyqv.cpu.instr_data[2][5] ),
    .S(_2563_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2567_));
 sky130_fd_sc_hd__clkbuf_1 _6003_ (.A(_2567_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0268_));
 sky130_fd_sc_hd__mux2_1 _6004_ (.A0(\i_tinyqv.cpu.instr_data_in[6] ),
    .A1(\i_tinyqv.cpu.instr_data[2][6] ),
    .S(_2563_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2568_));
 sky130_fd_sc_hd__clkbuf_1 _6005_ (.A(_2568_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0269_));
 sky130_fd_sc_hd__mux2_1 _6006_ (.A0(\i_tinyqv.cpu.instr_data_in[7] ),
    .A1(\i_tinyqv.cpu.instr_data[2][7] ),
    .S(_2563_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2569_));
 sky130_fd_sc_hd__clkbuf_1 _6007_ (.A(_2569_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0270_));
 sky130_fd_sc_hd__mux2_1 _6008_ (.A0(_2316_),
    .A1(\i_tinyqv.cpu.instr_data[2][8] ),
    .S(_2563_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2570_));
 sky130_fd_sc_hd__clkbuf_1 _6009_ (.A(_2570_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0271_));
 sky130_fd_sc_hd__mux2_1 _6010_ (.A0(_2318_),
    .A1(\i_tinyqv.cpu.instr_data[2][9] ),
    .S(_2563_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2571_));
 sky130_fd_sc_hd__clkbuf_1 _6011_ (.A(_2571_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0272_));
 sky130_fd_sc_hd__mux2_1 _6012_ (.A0(_2320_),
    .A1(\i_tinyqv.cpu.instr_data[2][10] ),
    .S(_2563_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2572_));
 sky130_fd_sc_hd__clkbuf_1 _6013_ (.A(_2572_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0273_));
 sky130_fd_sc_hd__mux2_1 _6014_ (.A0(_2322_),
    .A1(\i_tinyqv.cpu.instr_data[2][11] ),
    .S(_2563_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2573_));
 sky130_fd_sc_hd__clkbuf_1 _6015_ (.A(_2573_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0274_));
 sky130_fd_sc_hd__mux2_1 _6016_ (.A0(_1712_),
    .A1(\i_tinyqv.cpu.instr_data[2][12] ),
    .S(_2562_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2574_));
 sky130_fd_sc_hd__clkbuf_1 _6017_ (.A(_2574_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0275_));
 sky130_fd_sc_hd__mux2_1 _6018_ (.A0(_1717_),
    .A1(\i_tinyqv.cpu.instr_data[2][13] ),
    .S(_2562_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2575_));
 sky130_fd_sc_hd__clkbuf_1 _6019_ (.A(_2575_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0276_));
 sky130_fd_sc_hd__mux2_1 _6020_ (.A0(_1720_),
    .A1(\i_tinyqv.cpu.instr_data[2][14] ),
    .S(_2562_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2576_));
 sky130_fd_sc_hd__clkbuf_1 _6021_ (.A(_2576_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0277_));
 sky130_fd_sc_hd__mux2_1 _6022_ (.A0(_1721_),
    .A1(\i_tinyqv.cpu.instr_data[2][15] ),
    .S(_2562_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2577_));
 sky130_fd_sc_hd__clkbuf_1 _6023_ (.A(_2577_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0278_));
 sky130_fd_sc_hd__mux2_1 _6024_ (.A0(\i_tinyqv.cpu.instr_data_in[2] ),
    .A1(\i_tinyqv.cpu.instr_data[1][2] ),
    .S(_2463_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2578_));
 sky130_fd_sc_hd__clkbuf_1 _6025_ (.A(_2578_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0279_));
 sky130_fd_sc_hd__mux2_1 _6026_ (.A0(\i_tinyqv.cpu.instr_data_in[3] ),
    .A1(\i_tinyqv.cpu.instr_data[1][3] ),
    .S(_2463_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2579_));
 sky130_fd_sc_hd__clkbuf_1 _6027_ (.A(_2579_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0280_));
 sky130_fd_sc_hd__mux2_1 _6028_ (.A0(\i_tinyqv.cpu.instr_data_in[4] ),
    .A1(\i_tinyqv.cpu.instr_data[1][4] ),
    .S(_2463_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2580_));
 sky130_fd_sc_hd__clkbuf_1 _6029_ (.A(_2580_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0281_));
 sky130_fd_sc_hd__mux2_1 _6030_ (.A0(\i_tinyqv.cpu.instr_data_in[5] ),
    .A1(\i_tinyqv.cpu.instr_data[1][5] ),
    .S(_2463_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2581_));
 sky130_fd_sc_hd__clkbuf_1 _6031_ (.A(_2581_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0282_));
 sky130_fd_sc_hd__mux2_1 _6032_ (.A0(\i_tinyqv.cpu.instr_data_in[6] ),
    .A1(\i_tinyqv.cpu.instr_data[1][6] ),
    .S(_2463_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2582_));
 sky130_fd_sc_hd__clkbuf_1 _6033_ (.A(_2582_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0283_));
 sky130_fd_sc_hd__mux2_1 _6034_ (.A0(\i_tinyqv.cpu.instr_data_in[7] ),
    .A1(\i_tinyqv.cpu.instr_data[1][7] ),
    .S(_2463_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2583_));
 sky130_fd_sc_hd__clkbuf_1 _6035_ (.A(_2583_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0284_));
 sky130_fd_sc_hd__mux2_1 _6036_ (.A0(_2316_),
    .A1(\i_tinyqv.cpu.instr_data[1][8] ),
    .S(_2463_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2584_));
 sky130_fd_sc_hd__clkbuf_1 _6037_ (.A(_2584_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0285_));
 sky130_fd_sc_hd__mux2_1 _6038_ (.A0(_2318_),
    .A1(\i_tinyqv.cpu.instr_data[1][9] ),
    .S(_2463_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2585_));
 sky130_fd_sc_hd__clkbuf_1 _6039_ (.A(_2585_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0286_));
 sky130_fd_sc_hd__mux2_1 _6040_ (.A0(_2320_),
    .A1(\i_tinyqv.cpu.instr_data[1][10] ),
    .S(_2462_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2586_));
 sky130_fd_sc_hd__clkbuf_1 _6041_ (.A(_2586_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0287_));
 sky130_fd_sc_hd__mux2_1 _6042_ (.A0(_2322_),
    .A1(\i_tinyqv.cpu.instr_data[1][11] ),
    .S(_2462_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2587_));
 sky130_fd_sc_hd__clkbuf_1 _6043_ (.A(_2587_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0288_));
 sky130_fd_sc_hd__mux2_1 _6044_ (.A0(_1712_),
    .A1(\i_tinyqv.cpu.instr_data[1][12] ),
    .S(_2462_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2588_));
 sky130_fd_sc_hd__clkbuf_1 _6045_ (.A(_2588_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0289_));
 sky130_fd_sc_hd__mux2_1 _6046_ (.A0(_1717_),
    .A1(\i_tinyqv.cpu.instr_data[1][13] ),
    .S(_2462_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2589_));
 sky130_fd_sc_hd__clkbuf_1 _6047_ (.A(_2589_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0290_));
 sky130_fd_sc_hd__mux2_1 _6048_ (.A0(_1720_),
    .A1(\i_tinyqv.cpu.instr_data[1][14] ),
    .S(_2462_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2590_));
 sky130_fd_sc_hd__clkbuf_1 _6049_ (.A(_2590_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0291_));
 sky130_fd_sc_hd__mux2_1 _6050_ (.A0(_1721_),
    .A1(\i_tinyqv.cpu.instr_data[1][15] ),
    .S(_2462_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2591_));
 sky130_fd_sc_hd__clkbuf_1 _6051_ (.A(_2591_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0292_));
 sky130_fd_sc_hd__a21o_2 _6052_ (.A1(_1124_),
    .A2(_1563_),
    .B1(_1031_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2592_));
 sky130_fd_sc_hd__clkbuf_4 _6053_ (.A(_2592_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2593_));
 sky130_fd_sc_hd__mux2_1 _6054_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[0] ),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[4] ),
    .S(_2593_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2594_));
 sky130_fd_sc_hd__clkbuf_1 _6055_ (.A(_2594_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0293_));
 sky130_fd_sc_hd__a21oi_4 _6056_ (.A1(_1124_),
    .A2(_1563_),
    .B1(_1031_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2595_));
 sky130_fd_sc_hd__clkbuf_4 _6057_ (.A(_2595_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2596_));
 sky130_fd_sc_hd__mux2_1 _6058_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[5] ),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[1] ),
    .S(_2596_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2597_));
 sky130_fd_sc_hd__clkbuf_1 _6059_ (.A(_2597_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0294_));
 sky130_fd_sc_hd__mux2_1 _6060_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[6] ),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[2] ),
    .S(_2596_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2598_));
 sky130_fd_sc_hd__clkbuf_1 _6061_ (.A(_2598_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0295_));
 sky130_fd_sc_hd__mux2_1 _6062_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[3] ),
    .A1(_1054_),
    .S(_2593_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2599_));
 sky130_fd_sc_hd__clkbuf_1 _6063_ (.A(_2599_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0296_));
 sky130_fd_sc_hd__mux2_1 _6064_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[4] ),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[8] ),
    .S(_2593_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2600_));
 sky130_fd_sc_hd__clkbuf_1 _6065_ (.A(_2600_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0297_));
 sky130_fd_sc_hd__mux2_1 _6066_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[5] ),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[9] ),
    .S(_2593_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2601_));
 sky130_fd_sc_hd__clkbuf_1 _6067_ (.A(_2601_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0298_));
 sky130_fd_sc_hd__mux2_1 _6068_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[6] ),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[10] ),
    .S(_2593_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2602_));
 sky130_fd_sc_hd__clkbuf_1 _6069_ (.A(_2602_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0299_));
 sky130_fd_sc_hd__mux2_1 _6070_ (.A0(_1054_),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[11] ),
    .S(_2593_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2603_));
 sky130_fd_sc_hd__clkbuf_1 _6071_ (.A(_2603_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0300_));
 sky130_fd_sc_hd__mux2_1 _6072_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[8] ),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[12] ),
    .S(_2593_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2604_));
 sky130_fd_sc_hd__clkbuf_1 _6073_ (.A(_2604_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0301_));
 sky130_fd_sc_hd__mux2_1 _6074_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[9] ),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[13] ),
    .S(_2593_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2605_));
 sky130_fd_sc_hd__clkbuf_1 _6075_ (.A(_2605_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0302_));
 sky130_fd_sc_hd__mux2_1 _6076_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[10] ),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[14] ),
    .S(_2593_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2606_));
 sky130_fd_sc_hd__clkbuf_1 _6077_ (.A(_2606_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0303_));
 sky130_fd_sc_hd__mux2_1 _6078_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[11] ),
    .A1(_1060_),
    .S(_2593_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2607_));
 sky130_fd_sc_hd__clkbuf_1 _6079_ (.A(_2607_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0304_));
 sky130_fd_sc_hd__mux2_1 _6080_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[12] ),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[16] ),
    .S(_2592_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2608_));
 sky130_fd_sc_hd__clkbuf_1 _6081_ (.A(_2608_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0305_));
 sky130_fd_sc_hd__mux2_1 _6082_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[13] ),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[17] ),
    .S(_2592_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2609_));
 sky130_fd_sc_hd__clkbuf_1 _6083_ (.A(_2609_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0306_));
 sky130_fd_sc_hd__mux2_1 _6084_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[18] ),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[14] ),
    .S(_2596_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2610_));
 sky130_fd_sc_hd__clkbuf_1 _6085_ (.A(_2610_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0307_));
 sky130_fd_sc_hd__mux2_1 _6086_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[19] ),
    .A1(_1060_),
    .S(_2596_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2611_));
 sky130_fd_sc_hd__clkbuf_1 _6087_ (.A(_2611_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0308_));
 sky130_fd_sc_hd__mux2_1 _6088_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[20] ),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[16] ),
    .S(_2596_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2612_));
 sky130_fd_sc_hd__clkbuf_1 _6089_ (.A(_2612_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0309_));
 sky130_fd_sc_hd__mux2_1 _6090_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[21] ),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[17] ),
    .S(_2596_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2613_));
 sky130_fd_sc_hd__clkbuf_1 _6091_ (.A(_2613_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0310_));
 sky130_fd_sc_hd__mux2_1 _6092_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[22] ),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[18] ),
    .S(_2595_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2614_));
 sky130_fd_sc_hd__clkbuf_1 _6093_ (.A(_2614_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0311_));
 sky130_fd_sc_hd__mux2_1 _6094_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[23] ),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[19] ),
    .S(_2595_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2615_));
 sky130_fd_sc_hd__clkbuf_1 _6095_ (.A(_2615_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0312_));
 sky130_fd_sc_hd__mux2_1 _6096_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[24] ),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[20] ),
    .S(_2595_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2616_));
 sky130_fd_sc_hd__clkbuf_1 _6097_ (.A(_2616_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0313_));
 sky130_fd_sc_hd__mux2_1 _6098_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[25] ),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[21] ),
    .S(_2595_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2617_));
 sky130_fd_sc_hd__clkbuf_1 _6099_ (.A(_2617_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0314_));
 sky130_fd_sc_hd__mux2_1 _6100_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[26] ),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[22] ),
    .S(_2595_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2618_));
 sky130_fd_sc_hd__clkbuf_1 _6101_ (.A(_2618_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0315_));
 sky130_fd_sc_hd__mux2_1 _6102_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[27] ),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[23] ),
    .S(_2595_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2619_));
 sky130_fd_sc_hd__clkbuf_1 _6103_ (.A(_2619_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0316_));
 sky130_fd_sc_hd__mux2_1 _6104_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[28] ),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[24] ),
    .S(_2595_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2620_));
 sky130_fd_sc_hd__clkbuf_1 _6105_ (.A(_2620_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0317_));
 sky130_fd_sc_hd__mux2_1 _6106_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[25] ),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[29] ),
    .S(_2592_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2621_));
 sky130_fd_sc_hd__clkbuf_1 _6107_ (.A(_2621_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0318_));
 sky130_fd_sc_hd__mux2_1 _6108_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[26] ),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[30] ),
    .S(_2592_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2622_));
 sky130_fd_sc_hd__clkbuf_1 _6109_ (.A(_2622_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0319_));
 sky130_fd_sc_hd__mux2_1 _6110_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[31] ),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[27] ),
    .S(_2595_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2623_));
 sky130_fd_sc_hd__clkbuf_1 _6111_ (.A(_2623_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0320_));
 sky130_fd_sc_hd__or2_1 _6112_ (.A(_0846_),
    .B(_1755_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2624_));
 sky130_fd_sc_hd__clkbuf_2 _6113_ (.A(_2624_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2625_));
 sky130_fd_sc_hd__nand3b_1 _6114_ (.A_N(_2625_),
    .B(_1326_),
    .C(_1328_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2626_));
 sky130_fd_sc_hd__a21oi_1 _6115_ (.A1(net16),
    .A2(_2625_),
    .B1(_0845_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2627_));
 sky130_fd_sc_hd__a2bb2o_1 _6116_ (.A1_N(_0798_),
    .A2_N(_1124_),
    .B1(_2626_),
    .B2(_2627_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2628_));
 sky130_fd_sc_hd__nor2_1 _6117_ (.A(_2056_),
    .B(_2596_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2629_));
 sky130_fd_sc_hd__and4_1 _6118_ (.A(\i_tinyqv.cpu.i_core.mstatus_mte ),
    .B(_0744_),
    .C(_1394_),
    .D(_1392_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2630_));
 sky130_fd_sc_hd__a221o_1 _6119_ (.A1(\i_tinyqv.cpu.i_core.i_shift.a[30] ),
    .A2(_2596_),
    .B1(_2628_),
    .B2(_2629_),
    .C1(_2630_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0321_));
 sky130_fd_sc_hd__inv_2 _6120_ (.A(net49),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2631_));
 sky130_fd_sc_hd__mux2_1 _6121_ (.A0(_1569_),
    .A1(_2631_),
    .S(_2625_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2632_));
 sky130_fd_sc_hd__mux2_1 _6122_ (.A0(_0652_),
    .A1(_2632_),
    .S(_1124_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2633_));
 sky130_fd_sc_hd__a21bo_1 _6123_ (.A1(_1395_),
    .A2(_2633_),
    .B1_N(_2064_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2634_));
 sky130_fd_sc_hd__mux2_1 _6124_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[31] ),
    .A1(_2634_),
    .S(_2592_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2635_));
 sky130_fd_sc_hd__clkbuf_1 _6125_ (.A(_2635_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0322_));
 sky130_fd_sc_hd__or2_1 _6126_ (.A(_1400_),
    .B(\i_tinyqv.cpu.instr_data[0][0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2636_));
 sky130_fd_sc_hd__mux2_1 _6127_ (.A0(\i_tinyqv.cpu.instr_data_in[0] ),
    .A1(_2636_),
    .S(_2468_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2637_));
 sky130_fd_sc_hd__clkbuf_1 _6128_ (.A(_2637_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0323_));
 sky130_fd_sc_hd__or2_1 _6129_ (.A(_1400_),
    .B(\i_tinyqv.cpu.instr_data[0][1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2638_));
 sky130_fd_sc_hd__mux2_1 _6130_ (.A0(\i_tinyqv.cpu.instr_data_in[1] ),
    .A1(_2638_),
    .S(_2468_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2639_));
 sky130_fd_sc_hd__clkbuf_1 _6131_ (.A(_2639_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0324_));
 sky130_fd_sc_hd__and2_2 _6132_ (.A(_0714_),
    .B(net59),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2640_));
 sky130_fd_sc_hd__inv_2 _6133_ (.A(_2640_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2641_));
 sky130_fd_sc_hd__nand2_2 _6134_ (.A(_0653_),
    .B(\i_tinyqv.cpu.is_alu_imm ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2642_));
 sky130_fd_sc_hd__nor2_1 _6135_ (.A(_0707_),
    .B(_2642_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2643_));
 sky130_fd_sc_hd__a21o_1 _6136_ (.A1(_2641_),
    .A2(_2642_),
    .B1(_2643_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2644_));
 sky130_fd_sc_hd__nor2_2 _6137_ (.A(_1026_),
    .B(_1755_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2645_));
 sky130_fd_sc_hd__mux2_1 _6138_ (.A0(_1083_),
    .A1(_2644_),
    .S(_2645_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2646_));
 sky130_fd_sc_hd__clkbuf_1 _6139_ (.A(_2646_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0325_));
 sky130_fd_sc_hd__inv_2 _6140_ (.A(_0772_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2647_));
 sky130_fd_sc_hd__mux2_1 _6141_ (.A0(_0777_),
    .A1(_2647_),
    .S(_2642_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2648_));
 sky130_fd_sc_hd__mux2_1 _6142_ (.A0(_1149_),
    .A1(_2648_),
    .S(_2645_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2649_));
 sky130_fd_sc_hd__clkbuf_1 _6143_ (.A(_2649_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0326_));
 sky130_fd_sc_hd__mux2_1 _6144_ (.A0(_0814_),
    .A1(net16),
    .S(_2642_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2650_));
 sky130_fd_sc_hd__inv_2 _6145_ (.A(_2650_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2651_));
 sky130_fd_sc_hd__mux2_1 _6146_ (.A0(\i_tinyqv.cpu.i_core.i_shift.b[2] ),
    .A1(_2651_),
    .S(_2645_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2652_));
 sky130_fd_sc_hd__clkbuf_1 _6147_ (.A(_2652_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0327_));
 sky130_fd_sc_hd__o21a_1 _6148_ (.A1(_0956_),
    .A2(_0693_),
    .B1(_0696_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2653_));
 sky130_fd_sc_hd__mux2_1 _6149_ (.A0(_2653_),
    .A1(_2631_),
    .S(_2642_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2654_));
 sky130_fd_sc_hd__mux2_1 _6150_ (.A0(\i_tinyqv.cpu.i_core.i_shift.b[3] ),
    .A1(_2654_),
    .S(_2645_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2655_));
 sky130_fd_sc_hd__clkbuf_1 _6151_ (.A(_2655_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0328_));
 sky130_fd_sc_hd__buf_4 _6152_ (.A(_1386_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2656_));
 sky130_fd_sc_hd__mux2_1 _6153_ (.A0(\i_tinyqv.cpu.i_core.mepc[0] ),
    .A1(\i_tinyqv.cpu.i_core.mepc[4] ),
    .S(_2656_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2657_));
 sky130_fd_sc_hd__clkbuf_1 _6154_ (.A(_2657_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0329_));
 sky130_fd_sc_hd__mux2_1 _6155_ (.A0(\i_tinyqv.cpu.i_core.mepc[1] ),
    .A1(net264),
    .S(_2656_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2658_));
 sky130_fd_sc_hd__clkbuf_1 _6156_ (.A(_2658_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0330_));
 sky130_fd_sc_hd__mux2_1 _6157_ (.A0(\i_tinyqv.cpu.i_core.mepc[2] ),
    .A1(\i_tinyqv.cpu.i_core.mepc[6] ),
    .S(_2656_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2659_));
 sky130_fd_sc_hd__clkbuf_1 _6158_ (.A(_2659_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0331_));
 sky130_fd_sc_hd__mux2_1 _6159_ (.A0(\i_tinyqv.cpu.i_core.mepc[3] ),
    .A1(\i_tinyqv.cpu.i_core.mepc[7] ),
    .S(_2656_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2660_));
 sky130_fd_sc_hd__clkbuf_1 _6160_ (.A(_2660_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0332_));
 sky130_fd_sc_hd__mux2_1 _6161_ (.A0(\i_tinyqv.cpu.i_core.mepc[4] ),
    .A1(net232),
    .S(_2656_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2661_));
 sky130_fd_sc_hd__clkbuf_1 _6162_ (.A(_2661_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0333_));
 sky130_fd_sc_hd__mux2_1 _6163_ (.A0(\i_tinyqv.cpu.i_core.mepc[5] ),
    .A1(\i_tinyqv.cpu.i_core.mepc[9] ),
    .S(_2656_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2662_));
 sky130_fd_sc_hd__clkbuf_1 _6164_ (.A(_2662_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0334_));
 sky130_fd_sc_hd__mux2_1 _6165_ (.A0(\i_tinyqv.cpu.i_core.mepc[6] ),
    .A1(\i_tinyqv.cpu.i_core.mepc[10] ),
    .S(_2656_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2663_));
 sky130_fd_sc_hd__clkbuf_1 _6166_ (.A(_2663_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0335_));
 sky130_fd_sc_hd__mux2_1 _6167_ (.A0(\i_tinyqv.cpu.i_core.mepc[7] ),
    .A1(\i_tinyqv.cpu.i_core.mepc[11] ),
    .S(_2656_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2664_));
 sky130_fd_sc_hd__clkbuf_1 _6168_ (.A(_2664_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0336_));
 sky130_fd_sc_hd__mux2_1 _6169_ (.A0(\i_tinyqv.cpu.i_core.mepc[8] ),
    .A1(net228),
    .S(_2656_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2665_));
 sky130_fd_sc_hd__clkbuf_1 _6170_ (.A(_2665_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0337_));
 sky130_fd_sc_hd__mux2_1 _6171_ (.A0(\i_tinyqv.cpu.i_core.mepc[9] ),
    .A1(net226),
    .S(_2656_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2666_));
 sky130_fd_sc_hd__clkbuf_1 _6172_ (.A(_2666_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0338_));
 sky130_fd_sc_hd__clkbuf_4 _6173_ (.A(_1386_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2667_));
 sky130_fd_sc_hd__mux2_1 _6174_ (.A0(\i_tinyqv.cpu.i_core.mepc[10] ),
    .A1(\i_tinyqv.cpu.i_core.mepc[14] ),
    .S(_2667_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2668_));
 sky130_fd_sc_hd__clkbuf_1 _6175_ (.A(_2668_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0339_));
 sky130_fd_sc_hd__mux2_1 _6176_ (.A0(\i_tinyqv.cpu.i_core.mepc[11] ),
    .A1(\i_tinyqv.cpu.i_core.mepc[15] ),
    .S(_2667_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2669_));
 sky130_fd_sc_hd__clkbuf_1 _6177_ (.A(_2669_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0340_));
 sky130_fd_sc_hd__mux2_1 _6178_ (.A0(\i_tinyqv.cpu.i_core.mepc[12] ),
    .A1(\i_tinyqv.cpu.i_core.mepc[16] ),
    .S(_2667_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2670_));
 sky130_fd_sc_hd__clkbuf_1 _6179_ (.A(_2670_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0341_));
 sky130_fd_sc_hd__mux2_1 _6180_ (.A0(\i_tinyqv.cpu.i_core.mepc[13] ),
    .A1(\i_tinyqv.cpu.i_core.mepc[17] ),
    .S(_2667_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2671_));
 sky130_fd_sc_hd__clkbuf_1 _6181_ (.A(_2671_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0342_));
 sky130_fd_sc_hd__mux2_1 _6182_ (.A0(\i_tinyqv.cpu.i_core.mepc[14] ),
    .A1(\i_tinyqv.cpu.i_core.mepc[18] ),
    .S(_2667_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2672_));
 sky130_fd_sc_hd__clkbuf_1 _6183_ (.A(_2672_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0343_));
 sky130_fd_sc_hd__mux2_1 _6184_ (.A0(\i_tinyqv.cpu.i_core.mepc[15] ),
    .A1(\i_tinyqv.cpu.i_core.mepc[19] ),
    .S(_2667_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2673_));
 sky130_fd_sc_hd__clkbuf_1 _6185_ (.A(_2673_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0344_));
 sky130_fd_sc_hd__mux2_1 _6186_ (.A0(\i_tinyqv.cpu.i_core.mepc[16] ),
    .A1(\i_tinyqv.cpu.i_core.mepc[20] ),
    .S(_2667_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2674_));
 sky130_fd_sc_hd__clkbuf_1 _6187_ (.A(_2674_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0345_));
 sky130_fd_sc_hd__mux2_1 _6188_ (.A0(\i_tinyqv.cpu.i_core.mepc[17] ),
    .A1(\i_tinyqv.cpu.i_core.mepc[21] ),
    .S(_2667_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2675_));
 sky130_fd_sc_hd__clkbuf_1 _6189_ (.A(_2675_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0346_));
 sky130_fd_sc_hd__mux2_1 _6190_ (.A0(\i_tinyqv.cpu.i_core.mepc[18] ),
    .A1(\i_tinyqv.cpu.i_core.mepc[22] ),
    .S(_2667_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2676_));
 sky130_fd_sc_hd__clkbuf_1 _6191_ (.A(_2676_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0347_));
 sky130_fd_sc_hd__mux2_1 _6192_ (.A0(\i_tinyqv.cpu.i_core.mepc[19] ),
    .A1(\i_tinyqv.cpu.i_core.mepc[23] ),
    .S(_2667_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2677_));
 sky130_fd_sc_hd__clkbuf_1 _6193_ (.A(_2677_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0348_));
 sky130_fd_sc_hd__nor2_1 _6194_ (.A(_1551_),
    .B(_1541_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2678_));
 sky130_fd_sc_hd__and2_1 _6195_ (.A(_1536_),
    .B(_2678_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2679_));
 sky130_fd_sc_hd__or2_1 _6196_ (.A(\i_tinyqv.mem.instr_active ),
    .B(_2679_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2680_));
 sky130_fd_sc_hd__buf_4 _6197_ (.A(_2680_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2681_));
 sky130_fd_sc_hd__buf_4 _6198_ (.A(_2681_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2682_));
 sky130_fd_sc_hd__o2111a_1 _6199_ (.A1(_1540_),
    .A2(_2679_),
    .B1(_2682_),
    .C1(_1543_),
    .D1(_2221_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0349_));
 sky130_fd_sc_hd__and2_1 _6200_ (.A(\i_tinyqv.cpu.i_core.load_top_bit ),
    .B(_1026_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2683_));
 sky130_fd_sc_hd__nor2_1 _6201_ (.A(\i_tinyqv.cpu.i_core.mem_op[0] ),
    .B(_0939_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2684_));
 sky130_fd_sc_hd__a21oi_1 _6202_ (.A1(\i_tinyqv.cpu.i_core.mem_op[0] ),
    .A2(_0725_),
    .B1(_2684_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2685_));
 sky130_fd_sc_hd__or4_1 _6203_ (.A(\i_tinyqv.cpu.i_core.mem_op[1] ),
    .B(\i_tinyqv.cpu.i_core.mem_op[2] ),
    .C(_0878_),
    .D(_2685_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2686_));
 sky130_fd_sc_hd__mux2_1 _6204_ (.A0(_1635_),
    .A1(_2683_),
    .S(_2686_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2687_));
 sky130_fd_sc_hd__clkbuf_1 _6205_ (.A(_2687_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0350_));
 sky130_fd_sc_hd__mux2_1 _6206_ (.A0(net5),
    .A1(\i_debug_uart_tx.uart_tx_data[0] ),
    .S(_1728_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2688_));
 sky130_fd_sc_hd__a31o_1 _6207_ (.A1(_0984_),
    .A2(_0970_),
    .A3(_0995_),
    .B1(_2198_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2689_));
 sky130_fd_sc_hd__mux2_1 _6208_ (.A0(debug_register_data),
    .A1(_2688_),
    .S(_2689_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2690_));
 sky130_fd_sc_hd__clkbuf_1 _6209_ (.A(_2690_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0351_));
 sky130_fd_sc_hd__or4_1 _6210_ (.A(\i_tinyqv.mem.qspi_data_byte_idx[1] ),
    .B(_0868_),
    .C(_0979_),
    .D(_1536_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2691_));
 sky130_fd_sc_hd__mux2_1 _6211_ (.A0(_0871_),
    .A1(_0870_),
    .S(_0867_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2692_));
 sky130_fd_sc_hd__a22o_1 _6212_ (.A1(\i_tinyqv.mem.data_stall ),
    .A2(_2691_),
    .B1(_2692_),
    .B2(\i_tinyqv.mem.q_ctrl.data_req ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2693_));
 sky130_fd_sc_hd__o21a_1 _6213_ (.A1(_0977_),
    .A2(_2693_),
    .B1(net94),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0352_));
 sky130_fd_sc_hd__nand2_1 _6214_ (.A(\i_tinyqv.cpu.i_core.i_shift.a[13] ),
    .B(_1813_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2694_));
 sky130_fd_sc_hd__or2_1 _6215_ (.A(_1999_),
    .B(_2694_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2695_));
 sky130_fd_sc_hd__nand2_1 _6216_ (.A(\i_tinyqv.cpu.i_core.i_shift.a[14] ),
    .B(_1880_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2696_));
 sky130_fd_sc_hd__xnor2_1 _6217_ (.A(_2694_),
    .B(_2696_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2697_));
 sky130_fd_sc_hd__a21o_1 _6218_ (.A1(_2695_),
    .A2(_2026_),
    .B1(_2697_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2698_));
 sky130_fd_sc_hd__nand3_1 _6219_ (.A(_2695_),
    .B(_2026_),
    .C(_2697_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2699_));
 sky130_fd_sc_hd__nand2_1 _6220_ (.A(_2698_),
    .B(_2699_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2700_));
 sky130_fd_sc_hd__nand2_1 _6221_ (.A(_1060_),
    .B(_1845_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2701_));
 sky130_fd_sc_hd__xor2_1 _6222_ (.A(_2700_),
    .B(_2701_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2702_));
 sky130_fd_sc_hd__a21o_1 _6223_ (.A1(_2028_),
    .A2(_2030_),
    .B1(_2033_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2703_));
 sky130_fd_sc_hd__nand2_1 _6224_ (.A(_2702_),
    .B(_2703_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2704_));
 sky130_fd_sc_hd__or2_1 _6225_ (.A(_2702_),
    .B(_2703_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2705_));
 sky130_fd_sc_hd__and2_1 _6226_ (.A(_2704_),
    .B(_2705_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2706_));
 sky130_fd_sc_hd__o21ai_1 _6227_ (.A1(_2037_),
    .A2(_2038_),
    .B1(_2036_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2707_));
 sky130_fd_sc_hd__and2_1 _6228_ (.A(_2706_),
    .B(_2707_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2708_));
 sky130_fd_sc_hd__or2_1 _6229_ (.A(_2706_),
    .B(_2707_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2709_));
 sky130_fd_sc_hd__and2b_1 _6230_ (.A_N(_2708_),
    .B(_2709_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2710_));
 sky130_fd_sc_hd__a21bo_1 _6231_ (.A1(_2017_),
    .A2(_2044_),
    .B1_N(_2043_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2711_));
 sky130_fd_sc_hd__nand2_1 _6232_ (.A(_2041_),
    .B(_2711_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2712_));
 sky130_fd_sc_hd__xor2_1 _6233_ (.A(_2710_),
    .B(_2712_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0353_));
 sky130_fd_sc_hd__a21boi_2 _6234_ (.A1(_2041_),
    .A2(_2711_),
    .B1_N(_2710_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2713_));
 sky130_fd_sc_hd__nor2_1 _6235_ (.A(_2708_),
    .B(_2713_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2714_));
 sky130_fd_sc_hd__or2_1 _6236_ (.A(_2700_),
    .B(_2701_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2715_));
 sky130_fd_sc_hd__nand2_1 _6237_ (.A(_1060_),
    .B(_1880_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2716_));
 sky130_fd_sc_hd__and3_1 _6238_ (.A(\i_tinyqv.cpu.i_core.i_shift.a[14] ),
    .B(_1813_),
    .C(_2024_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2717_));
 sky130_fd_sc_hd__xor2_1 _6239_ (.A(_2716_),
    .B(_2717_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2718_));
 sky130_fd_sc_hd__a21oi_1 _6240_ (.A1(_2698_),
    .A2(_2715_),
    .B1(_2718_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2719_));
 sky130_fd_sc_hd__and3_1 _6241_ (.A(_2698_),
    .B(_2715_),
    .C(_2718_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2720_));
 sky130_fd_sc_hd__or2_1 _6242_ (.A(_2719_),
    .B(_2720_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2721_));
 sky130_fd_sc_hd__nor2_1 _6243_ (.A(_2704_),
    .B(_2721_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2722_));
 sky130_fd_sc_hd__nand2_1 _6244_ (.A(_2704_),
    .B(_2721_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2723_));
 sky130_fd_sc_hd__and2b_1 _6245_ (.A_N(_2722_),
    .B(_2723_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2724_));
 sky130_fd_sc_hd__xnor2_1 _6246_ (.A(_2714_),
    .B(_2724_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0354_));
 sky130_fd_sc_hd__and3_1 _6247_ (.A(_1060_),
    .B(_1813_),
    .C(_2696_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2725_));
 sky130_fd_sc_hd__inv_2 _6248_ (.A(_2719_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2726_));
 sky130_fd_sc_hd__o31a_1 _6249_ (.A1(_1060_),
    .A2(_2694_),
    .A3(_2696_),
    .B1(_2726_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2727_));
 sky130_fd_sc_hd__xnor2_1 _6250_ (.A(_2725_),
    .B(_2727_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2728_));
 sky130_fd_sc_hd__o31a_1 _6251_ (.A1(_2708_),
    .A2(_2713_),
    .A3(_2722_),
    .B1(_2723_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2729_));
 sky130_fd_sc_hd__xor2_1 _6252_ (.A(_2728_),
    .B(_2729_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0355_));
 sky130_fd_sc_hd__nand2_1 _6253_ (.A(_2696_),
    .B(_2726_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2730_));
 sky130_fd_sc_hd__o311a_1 _6254_ (.A1(_2708_),
    .A2(_2713_),
    .A3(_2722_),
    .B1(_2723_),
    .C1(_2728_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2731_));
 sky130_fd_sc_hd__a31o_1 _6255_ (.A1(_1060_),
    .A2(_1813_),
    .A3(_2730_),
    .B1(_2731_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0356_));
 sky130_fd_sc_hd__a21o_4 _6256_ (.A1(_1551_),
    .A2(_1536_),
    .B1(_1541_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2732_));
 sky130_fd_sc_hd__clkbuf_4 _6257_ (.A(_2732_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2733_));
 sky130_fd_sc_hd__nor2_2 _6258_ (.A(\i_tinyqv.mem.instr_active ),
    .B(_2679_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2734_));
 sky130_fd_sc_hd__nor2_1 _6259_ (.A(\i_tinyqv.mem.q_ctrl.data_ready ),
    .B(\i_tinyqv.mem.q_ctrl.data_req ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2735_));
 sky130_fd_sc_hd__a21oi_1 _6260_ (.A1(_0872_),
    .A2(_2734_),
    .B1(_2735_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2736_));
 sky130_fd_sc_hd__mux2_1 _6261_ (.A0(_2736_),
    .A1(_2735_),
    .S(_0868_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2737_));
 sky130_fd_sc_hd__and3_1 _6262_ (.A(_2181_),
    .B(_2733_),
    .C(_2737_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2738_));
 sky130_fd_sc_hd__clkbuf_1 _6263_ (.A(_2738_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0357_));
 sky130_fd_sc_hd__or3b_1 _6264_ (.A(_2681_),
    .B(_1016_),
    .C_N(_1531_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2739_));
 sky130_fd_sc_hd__o21ai_1 _6265_ (.A1(_0864_),
    .A2(_0868_),
    .B1(_2739_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2740_));
 sky130_fd_sc_hd__a22o_1 _6266_ (.A1(\i_tinyqv.mem.qspi_data_byte_idx[1] ),
    .A2(_2735_),
    .B1(_2736_),
    .B2(_2740_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2741_));
 sky130_fd_sc_hd__and3_1 _6267_ (.A(_2181_),
    .B(_2733_),
    .C(_2741_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2742_));
 sky130_fd_sc_hd__clkbuf_1 _6268_ (.A(_2742_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0358_));
 sky130_fd_sc_hd__or3b_1 _6269_ (.A(\i_tinyqv.mem.qspi_data_byte_idx[1] ),
    .B(_0868_),
    .C_N(\i_tinyqv.mem.q_ctrl.data_ready ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2743_));
 sky130_fd_sc_hd__clkbuf_4 _6270_ (.A(_2743_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2744_));
 sky130_fd_sc_hd__mux2_1 _6271_ (.A0(_2316_),
    .A1(\i_tinyqv.cpu.instr_data_in[0] ),
    .S(_2744_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2745_));
 sky130_fd_sc_hd__clkbuf_1 _6272_ (.A(_2745_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0359_));
 sky130_fd_sc_hd__mux2_1 _6273_ (.A0(_2318_),
    .A1(\i_tinyqv.cpu.instr_data_in[1] ),
    .S(_2744_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2746_));
 sky130_fd_sc_hd__clkbuf_1 _6274_ (.A(_2746_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0360_));
 sky130_fd_sc_hd__mux2_1 _6275_ (.A0(_2320_),
    .A1(\i_tinyqv.cpu.instr_data_in[2] ),
    .S(_2744_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2747_));
 sky130_fd_sc_hd__clkbuf_1 _6276_ (.A(_2747_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0361_));
 sky130_fd_sc_hd__mux2_1 _6277_ (.A0(_2322_),
    .A1(\i_tinyqv.cpu.instr_data_in[3] ),
    .S(_2744_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2748_));
 sky130_fd_sc_hd__clkbuf_1 _6278_ (.A(_2748_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0362_));
 sky130_fd_sc_hd__mux2_1 _6279_ (.A0(_1712_),
    .A1(\i_tinyqv.cpu.instr_data_in[4] ),
    .S(_2744_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2749_));
 sky130_fd_sc_hd__clkbuf_1 _6280_ (.A(_2749_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0363_));
 sky130_fd_sc_hd__mux2_1 _6281_ (.A0(_1717_),
    .A1(\i_tinyqv.cpu.instr_data_in[5] ),
    .S(_2744_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2750_));
 sky130_fd_sc_hd__clkbuf_1 _6282_ (.A(_2750_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0364_));
 sky130_fd_sc_hd__mux2_1 _6283_ (.A0(_1720_),
    .A1(\i_tinyqv.cpu.instr_data_in[6] ),
    .S(_2744_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2751_));
 sky130_fd_sc_hd__clkbuf_1 _6284_ (.A(_2751_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0365_));
 sky130_fd_sc_hd__mux2_1 _6285_ (.A0(_1721_),
    .A1(\i_tinyqv.cpu.instr_data_in[7] ),
    .S(_2744_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2752_));
 sky130_fd_sc_hd__clkbuf_1 _6286_ (.A(_2752_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0366_));
 sky130_fd_sc_hd__mux2_1 _6287_ (.A0(net275),
    .A1(_2316_),
    .S(_1552_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2753_));
 sky130_fd_sc_hd__clkbuf_1 _6288_ (.A(_2753_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0367_));
 sky130_fd_sc_hd__mux2_1 _6289_ (.A0(\i_tinyqv.mem.qspi_data_buf[9] ),
    .A1(_2318_),
    .S(_1552_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2754_));
 sky130_fd_sc_hd__clkbuf_1 _6290_ (.A(_2754_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0368_));
 sky130_fd_sc_hd__mux2_1 _6291_ (.A0(\i_tinyqv.mem.qspi_data_buf[10] ),
    .A1(_2320_),
    .S(_1552_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2755_));
 sky130_fd_sc_hd__clkbuf_1 _6292_ (.A(_2755_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0369_));
 sky130_fd_sc_hd__mux2_1 _6293_ (.A0(net229),
    .A1(_2322_),
    .S(_1552_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2756_));
 sky130_fd_sc_hd__clkbuf_1 _6294_ (.A(_2756_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0370_));
 sky130_fd_sc_hd__mux2_1 _6295_ (.A0(net293),
    .A1(_1712_),
    .S(_1552_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2757_));
 sky130_fd_sc_hd__clkbuf_1 _6296_ (.A(_2757_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0371_));
 sky130_fd_sc_hd__mux2_1 _6297_ (.A0(\i_tinyqv.mem.qspi_data_buf[13] ),
    .A1(_1717_),
    .S(_1552_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2758_));
 sky130_fd_sc_hd__clkbuf_1 _6298_ (.A(_2758_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0372_));
 sky130_fd_sc_hd__mux2_1 _6299_ (.A0(\i_tinyqv.mem.qspi_data_buf[14] ),
    .A1(_1720_),
    .S(_1552_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2759_));
 sky130_fd_sc_hd__clkbuf_1 _6300_ (.A(_2759_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0373_));
 sky130_fd_sc_hd__mux2_1 _6301_ (.A0(net256),
    .A1(_1721_),
    .S(_1552_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2760_));
 sky130_fd_sc_hd__clkbuf_1 _6302_ (.A(_2760_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0374_));
 sky130_fd_sc_hd__and3b_1 _6303_ (.A_N(_0868_),
    .B(\i_tinyqv.mem.q_ctrl.data_ready ),
    .C(\i_tinyqv.mem.qspi_data_byte_idx[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2761_));
 sky130_fd_sc_hd__clkbuf_4 _6304_ (.A(_2761_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2762_));
 sky130_fd_sc_hd__mux2_1 _6305_ (.A0(net280),
    .A1(_2316_),
    .S(_2762_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2763_));
 sky130_fd_sc_hd__clkbuf_1 _6306_ (.A(_2763_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0375_));
 sky130_fd_sc_hd__mux2_1 _6307_ (.A0(net277),
    .A1(_2318_),
    .S(_2762_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2764_));
 sky130_fd_sc_hd__clkbuf_1 _6308_ (.A(_2764_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0376_));
 sky130_fd_sc_hd__mux2_1 _6309_ (.A0(net269),
    .A1(_2320_),
    .S(_2762_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2765_));
 sky130_fd_sc_hd__clkbuf_1 _6310_ (.A(_2765_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0377_));
 sky130_fd_sc_hd__mux2_1 _6311_ (.A0(net245),
    .A1(_2322_),
    .S(_2762_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2766_));
 sky130_fd_sc_hd__clkbuf_1 _6312_ (.A(_2766_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0378_));
 sky130_fd_sc_hd__mux2_1 _6313_ (.A0(net292),
    .A1(_1712_),
    .S(_2762_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2767_));
 sky130_fd_sc_hd__clkbuf_1 _6314_ (.A(_2767_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0379_));
 sky130_fd_sc_hd__mux2_1 _6315_ (.A0(\i_tinyqv.mem.data_from_read[21] ),
    .A1(_1717_),
    .S(_2762_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2768_));
 sky130_fd_sc_hd__clkbuf_1 _6316_ (.A(_2768_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0380_));
 sky130_fd_sc_hd__mux2_1 _6317_ (.A0(\i_tinyqv.mem.data_from_read[22] ),
    .A1(_1720_),
    .S(_2762_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2769_));
 sky130_fd_sc_hd__clkbuf_1 _6318_ (.A(_2769_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0381_));
 sky130_fd_sc_hd__mux2_1 _6319_ (.A0(net285),
    .A1(_1721_),
    .S(_2762_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2770_));
 sky130_fd_sc_hd__clkbuf_1 _6320_ (.A(_2770_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0382_));
 sky130_fd_sc_hd__and3_1 _6321_ (.A(\i_tinyqv.mem.qspi_data_byte_idx[1] ),
    .B(_0868_),
    .C(\i_tinyqv.mem.q_ctrl.data_ready ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2771_));
 sky130_fd_sc_hd__clkbuf_4 _6322_ (.A(_2771_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2772_));
 sky130_fd_sc_hd__mux2_1 _6323_ (.A0(net279),
    .A1(_2316_),
    .S(_2772_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2773_));
 sky130_fd_sc_hd__clkbuf_1 _6324_ (.A(_2773_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0383_));
 sky130_fd_sc_hd__mux2_1 _6325_ (.A0(net286),
    .A1(_2318_),
    .S(_2772_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2774_));
 sky130_fd_sc_hd__clkbuf_1 _6326_ (.A(_2774_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0384_));
 sky130_fd_sc_hd__mux2_1 _6327_ (.A0(net267),
    .A1(_2320_),
    .S(_2772_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2775_));
 sky130_fd_sc_hd__clkbuf_1 _6328_ (.A(_2775_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0385_));
 sky130_fd_sc_hd__mux2_1 _6329_ (.A0(net253),
    .A1(_2322_),
    .S(_2772_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2776_));
 sky130_fd_sc_hd__clkbuf_1 _6330_ (.A(_2776_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0386_));
 sky130_fd_sc_hd__mux2_1 _6331_ (.A0(net276),
    .A1(_1712_),
    .S(_2772_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2777_));
 sky130_fd_sc_hd__clkbuf_1 _6332_ (.A(_2777_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0387_));
 sky130_fd_sc_hd__mux2_1 _6333_ (.A0(net287),
    .A1(_1717_),
    .S(_2772_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2778_));
 sky130_fd_sc_hd__clkbuf_1 _6334_ (.A(_2778_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0388_));
 sky130_fd_sc_hd__mux2_1 _6335_ (.A0(net290),
    .A1(_1720_),
    .S(_2772_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2779_));
 sky130_fd_sc_hd__clkbuf_1 _6336_ (.A(_2779_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0389_));
 sky130_fd_sc_hd__mux2_1 _6337_ (.A0(net261),
    .A1(_1721_),
    .S(_2772_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2780_));
 sky130_fd_sc_hd__clkbuf_1 _6338_ (.A(_2780_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0390_));
 sky130_fd_sc_hd__and3_1 _6339_ (.A(_2181_),
    .B(_1536_),
    .C(_2678_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2781_));
 sky130_fd_sc_hd__clkbuf_1 _6340_ (.A(_2781_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0391_));
 sky130_fd_sc_hd__or2_1 _6341_ (.A(\i_tinyqv.mem.q_ctrl.read_cycles_count[1] ),
    .B(\i_tinyqv.mem.q_ctrl.read_cycles_count[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2782_));
 sky130_fd_sc_hd__or2b_2 _6342_ (.A(\i_tinyqv.mem.data_stall ),
    .B_N(_1532_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2783_));
 sky130_fd_sc_hd__nor2_1 _6343_ (.A(_2782_),
    .B(_2783_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2784_));
 sky130_fd_sc_hd__nand2_1 _6344_ (.A(_1706_),
    .B(\i_tinyqv.mem.q_ctrl.fsm_state[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2785_));
 sky130_fd_sc_hd__or2_1 _6345_ (.A(_1707_),
    .B(_2785_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2786_));
 sky130_fd_sc_hd__buf_2 _6346_ (.A(_2786_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2787_));
 sky130_fd_sc_hd__nor2_1 _6347_ (.A(_1713_),
    .B(_2787_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2788_));
 sky130_fd_sc_hd__and3_1 _6348_ (.A(\i_tinyqv.mem.q_ctrl.fsm_state[2] ),
    .B(\i_tinyqv.mem.q_ctrl.fsm_state[1] ),
    .C(_1707_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2789_));
 sky130_fd_sc_hd__or2_1 _6349_ (.A(_1711_),
    .B(_2789_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2790_));
 sky130_fd_sc_hd__or2_1 _6350_ (.A(\i_tinyqv.mem.q_ctrl.read_cycles_count[0] ),
    .B(_2782_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2791_));
 sky130_fd_sc_hd__inv_2 _6351_ (.A(\i_tinyqv.mem.q_ctrl.is_writing ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2792_));
 sky130_fd_sc_hd__a21o_1 _6352_ (.A1(_2792_),
    .A2(_1711_),
    .B1(_2789_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2793_));
 sky130_fd_sc_hd__mux2_2 _6353_ (.A0(_2302_),
    .A1(_2791_),
    .S(_2793_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2794_));
 sky130_fd_sc_hd__or3_4 _6354_ (.A(\i_tinyqv.mem.q_ctrl.nibbles_remaining[2] ),
    .B(\i_tinyqv.mem.q_ctrl.nibbles_remaining[1] ),
    .C(\i_tinyqv.mem.q_ctrl.nibbles_remaining[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2795_));
 sky130_fd_sc_hd__inv_2 _6355_ (.A(\i_tinyqv.mem.q_ctrl.read_cycles_count[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2796_));
 sky130_fd_sc_hd__or3b_2 _6356_ (.A(\i_tinyqv.mem.q_ctrl.fsm_state[1] ),
    .B(_1707_),
    .C_N(_1706_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2797_));
 sky130_fd_sc_hd__mux2_1 _6357_ (.A0(\i_tinyqv.mem.q_ctrl.delay_cycles_cfg[0] ),
    .A1(_2796_),
    .S(_2797_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2798_));
 sky130_fd_sc_hd__or4_1 _6358_ (.A(_2790_),
    .B(_2794_),
    .C(_2795_),
    .D(_2798_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2799_));
 sky130_fd_sc_hd__nand2_2 _6359_ (.A(_1706_),
    .B(_1707_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2800_));
 sky130_fd_sc_hd__or2_2 _6360_ (.A(_2800_),
    .B(_2783_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2801_));
 sky130_fd_sc_hd__nand2_1 _6361_ (.A(\i_tinyqv.mem.q_ctrl.delay_cycles_cfg[2] ),
    .B(_2789_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2802_));
 sky130_fd_sc_hd__and2_2 _6362_ (.A(_2795_),
    .B(_2802_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2803_));
 sky130_fd_sc_hd__nor2_1 _6363_ (.A(_2794_),
    .B(_2803_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2804_));
 sky130_fd_sc_hd__nand2_1 _6364_ (.A(_2787_),
    .B(_2799_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2805_));
 sky130_fd_sc_hd__or2_1 _6365_ (.A(_2786_),
    .B(_2784_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2806_));
 sky130_fd_sc_hd__a21oi_1 _6366_ (.A1(_2805_),
    .A2(_2806_),
    .B1(\i_tinyqv.mem.q_ctrl.read_cycles_count[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2807_));
 sky130_fd_sc_hd__a41o_1 _6367_ (.A1(_2787_),
    .A2(_2799_),
    .A3(_2801_),
    .A4(_2804_),
    .B1(_2807_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2808_));
 sky130_fd_sc_hd__a31o_1 _6368_ (.A1(\i_tinyqv.mem.q_ctrl.delay_cycles_cfg[0] ),
    .A2(_2784_),
    .A3(_2788_),
    .B1(_2808_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2809_));
 sky130_fd_sc_hd__inv_2 _6369_ (.A(_1540_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2810_));
 sky130_fd_sc_hd__nor2_2 _6370_ (.A(_2810_),
    .B(_2305_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2811_));
 sky130_fd_sc_hd__mux2_1 _6371_ (.A0(\i_tinyqv.mem.q_ctrl.read_cycles_count[0] ),
    .A1(_2809_),
    .S(_2811_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2812_));
 sky130_fd_sc_hd__clkbuf_1 _6372_ (.A(_2812_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0392_));
 sky130_fd_sc_hd__nor2_1 _6373_ (.A(_1707_),
    .B(_2785_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2813_));
 sky130_fd_sc_hd__a21oi_1 _6374_ (.A1(_2796_),
    .A2(\i_tinyqv.mem.q_ctrl.read_cycles_count[2] ),
    .B1(\i_tinyqv.mem.q_ctrl.read_cycles_count[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2814_));
 sky130_fd_sc_hd__a21oi_2 _6375_ (.A1(_2796_),
    .A2(\i_tinyqv.mem.q_ctrl.read_cycles_count[1] ),
    .B1(_2814_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2815_));
 sky130_fd_sc_hd__mux2_1 _6376_ (.A0(_2815_),
    .A1(\i_tinyqv.mem.q_ctrl.delay_cycles_cfg[1] ),
    .S(_2783_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2816_));
 sky130_fd_sc_hd__mux2_1 _6377_ (.A0(\i_tinyqv.mem.q_ctrl.delay_cycles_cfg[1] ),
    .A1(_2815_),
    .S(_2797_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2817_));
 sky130_fd_sc_hd__mux2_1 _6378_ (.A0(_2816_),
    .A1(_2817_),
    .S(_2800_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2818_));
 sky130_fd_sc_hd__mux2_1 _6379_ (.A0(_2815_),
    .A1(_2818_),
    .S(_2804_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2819_));
 sky130_fd_sc_hd__a31o_1 _6380_ (.A1(_2792_),
    .A2(\i_tinyqv.mem.q_ctrl.delay_cycles_cfg[2] ),
    .A3(_2784_),
    .B1(_2787_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2820_));
 sky130_fd_sc_hd__o22a_1 _6381_ (.A1(_2813_),
    .A2(_2819_),
    .B1(_2820_),
    .B2(_2815_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2821_));
 sky130_fd_sc_hd__mux2_1 _6382_ (.A0(\i_tinyqv.mem.q_ctrl.read_cycles_count[1] ),
    .A1(_2821_),
    .S(_2811_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2822_));
 sky130_fd_sc_hd__clkbuf_1 _6383_ (.A(_2822_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0393_));
 sky130_fd_sc_hd__o21a_1 _6384_ (.A1(\i_tinyqv.mem.q_ctrl.read_cycles_count[0] ),
    .A2(\i_tinyqv.mem.q_ctrl.read_cycles_count[1] ),
    .B1(\i_tinyqv.mem.q_ctrl.read_cycles_count[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2823_));
 sky130_fd_sc_hd__mux2_1 _6385_ (.A0(\i_tinyqv.mem.q_ctrl.delay_cycles_cfg[2] ),
    .A1(_2823_),
    .S(_2797_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2824_));
 sky130_fd_sc_hd__inv_2 _6386_ (.A(_2804_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2825_));
 sky130_fd_sc_hd__a31o_1 _6387_ (.A1(\i_tinyqv.mem.q_ctrl.delay_cycles_cfg[2] ),
    .A2(_2790_),
    .A3(_2783_),
    .B1(_2825_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2826_));
 sky130_fd_sc_hd__a21oi_1 _6388_ (.A1(_2800_),
    .A2(_2824_),
    .B1(_2826_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2827_));
 sky130_fd_sc_hd__o21ai_1 _6389_ (.A1(_2804_),
    .A2(_2823_),
    .B1(_2787_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2828_));
 sky130_fd_sc_hd__o21ai_1 _6390_ (.A1(_2801_),
    .A2(_2828_),
    .B1(_2806_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2829_));
 sky130_fd_sc_hd__a2bb2o_1 _6391_ (.A1_N(_2827_),
    .A2_N(_2828_),
    .B1(_2823_),
    .B2(_2829_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2830_));
 sky130_fd_sc_hd__mux2_1 _6392_ (.A0(\i_tinyqv.mem.q_ctrl.read_cycles_count[2] ),
    .A1(_2830_),
    .S(_2811_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2831_));
 sky130_fd_sc_hd__clkbuf_1 _6393_ (.A(_2831_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0394_));
 sky130_fd_sc_hd__buf_2 _6394_ (.A(_2304_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2832_));
 sky130_fd_sc_hd__inv_2 _6395_ (.A(_2795_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2833_));
 sky130_fd_sc_hd__and3_1 _6396_ (.A(_1713_),
    .B(_1711_),
    .C(_2794_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2834_));
 sky130_fd_sc_hd__and3_1 _6397_ (.A(_2832_),
    .B(_2833_),
    .C(_2834_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2835_));
 sky130_fd_sc_hd__clkbuf_1 _6398_ (.A(_2835_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0395_));
 sky130_fd_sc_hd__nand2_1 _6399_ (.A(_1540_),
    .B(_2787_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2836_));
 sky130_fd_sc_hd__nor2_1 _6400_ (.A(_2794_),
    .B(_2836_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2837_));
 sky130_fd_sc_hd__or3b_2 _6401_ (.A(\i_tinyqv.cpu.data_addr[23] ),
    .B(_2681_),
    .C_N(\i_tinyqv.cpu.data_addr[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2838_));
 sky130_fd_sc_hd__and4b_1 _6402_ (.A_N(\i_tinyqv.mem.q_ctrl.last_ram_b_sel ),
    .B(_2734_),
    .C(\i_tinyqv.cpu.data_addr[24] ),
    .D(\i_tinyqv.cpu.data_addr[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2839_));
 sky130_fd_sc_hd__nor2_2 _6403_ (.A(_2732_),
    .B(_2839_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2840_));
 sky130_fd_sc_hd__o21a_1 _6404_ (.A1(\i_tinyqv.mem.q_ctrl.last_ram_a_sel ),
    .A2(_2838_),
    .B1(_2840_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2841_));
 sky130_fd_sc_hd__or2_1 _6405_ (.A(_2837_),
    .B(_2841_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2842_));
 sky130_fd_sc_hd__a31o_1 _6406_ (.A1(\i_tinyqv.mem.q_ctrl.nibbles_remaining[0] ),
    .A2(_2802_),
    .A3(_2837_),
    .B1(_2305_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2843_));
 sky130_fd_sc_hd__o21ba_1 _6407_ (.A1(\i_tinyqv.mem.q_ctrl.nibbles_remaining[0] ),
    .A2(_2842_),
    .B1_N(_2843_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0396_));
 sky130_fd_sc_hd__nor2_1 _6408_ (.A(_2837_),
    .B(_2841_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2844_));
 sky130_fd_sc_hd__and3_1 _6409_ (.A(\i_tinyqv.mem.q_ctrl.spi_flash_select ),
    .B(_2792_),
    .C(_1709_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2845_));
 sky130_fd_sc_hd__and2_1 _6410_ (.A(\i_tinyqv.mem.q_ctrl.fsm_state[1] ),
    .B(_1707_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2846_));
 sky130_fd_sc_hd__and2b_1 _6411_ (.A_N(_1706_),
    .B(_2846_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2847_));
 sky130_fd_sc_hd__o21ai_1 _6412_ (.A1(\i_tinyqv.mem.q_ctrl.nibbles_remaining[1] ),
    .A2(\i_tinyqv.mem.q_ctrl.nibbles_remaining[0] ),
    .B1(_2802_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2848_));
 sky130_fd_sc_hd__a21o_1 _6413_ (.A1(\i_tinyqv.mem.q_ctrl.nibbles_remaining[1] ),
    .A2(\i_tinyqv.mem.q_ctrl.nibbles_remaining[0] ),
    .B1(_2848_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2849_));
 sky130_fd_sc_hd__o311a_1 _6414_ (.A1(_2803_),
    .A2(_2845_),
    .A3(_2847_),
    .B1(_2849_),
    .C1(_2837_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2850_));
 sky130_fd_sc_hd__a32o_1 _6415_ (.A1(net265),
    .A2(_2832_),
    .A3(_2844_),
    .B1(_2850_),
    .B2(_2811_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0397_));
 sky130_fd_sc_hd__inv_2 _6416_ (.A(\i_tinyqv.mem.q_ctrl.nibbles_remaining[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2851_));
 sky130_fd_sc_hd__o22ai_1 _6417_ (.A1(_1715_),
    .A2(_2803_),
    .B1(_2848_),
    .B2(_2851_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2852_));
 sky130_fd_sc_hd__a21oi_2 _6418_ (.A1(\i_tinyqv.cpu.data_addr[24] ),
    .A2(_2734_),
    .B1(_1540_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2853_));
 sky130_fd_sc_hd__a211o_1 _6419_ (.A1(_1540_),
    .A2(_2852_),
    .B1(_2853_),
    .C1(_2844_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2854_));
 sky130_fd_sc_hd__o211a_1 _6420_ (.A1(\i_tinyqv.mem.q_ctrl.nibbles_remaining[2] ),
    .A2(_2842_),
    .B1(_2854_),
    .C1(_2832_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0398_));
 sky130_fd_sc_hd__o21ai_4 _6421_ (.A1(\i_tinyqv.mem.q_ctrl.last_ram_a_sel ),
    .A2(_2838_),
    .B1(_2840_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2855_));
 sky130_fd_sc_hd__a211o_1 _6422_ (.A1(\i_tinyqv.cpu.data_read_n[1] ),
    .A2(\i_tinyqv.cpu.data_read_n[0] ),
    .B1(_0957_),
    .C1(_1541_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2856_));
 sky130_fd_sc_hd__and3_1 _6423_ (.A(\i_tinyqv.cpu.data_addr[24] ),
    .B(_2734_),
    .C(_2841_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2857_));
 sky130_fd_sc_hd__a22o_1 _6424_ (.A1(_1713_),
    .A2(_2855_),
    .B1(_2856_),
    .B2(_2857_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2858_));
 sky130_fd_sc_hd__and2_1 _6425_ (.A(_2832_),
    .B(_2858_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2859_));
 sky130_fd_sc_hd__clkbuf_1 _6426_ (.A(_2859_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0399_));
 sky130_fd_sc_hd__inv_2 _6427_ (.A(_2794_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2860_));
 sky130_fd_sc_hd__and3_1 _6428_ (.A(_2785_),
    .B(_2860_),
    .C(_2803_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2861_));
 sky130_fd_sc_hd__o21ai_1 _6429_ (.A1(_2810_),
    .A2(_2861_),
    .B1(_2855_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2862_));
 sky130_fd_sc_hd__o211a_1 _6430_ (.A1(_2860_),
    .A2(_2836_),
    .B1(_2862_),
    .C1(_2806_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2863_));
 sky130_fd_sc_hd__nand2_1 _6431_ (.A(_2795_),
    .B(_2802_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2864_));
 sky130_fd_sc_hd__o211a_1 _6432_ (.A1(_1707_),
    .A2(_2845_),
    .B1(_2864_),
    .C1(_2801_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2865_));
 sky130_fd_sc_hd__o21ai_1 _6433_ (.A1(_2853_),
    .A2(_2865_),
    .B1(_2863_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2866_));
 sky130_fd_sc_hd__o211a_1 _6434_ (.A1(_1707_),
    .A2(_2863_),
    .B1(_2866_),
    .C1(_2832_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0400_));
 sky130_fd_sc_hd__o21a_1 _6435_ (.A1(\i_tinyqv.mem.q_ctrl.spi_flash_select ),
    .A2(_1713_),
    .B1(_1709_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2867_));
 sky130_fd_sc_hd__a21oi_1 _6436_ (.A1(_1714_),
    .A2(_1708_),
    .B1(_2867_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2868_));
 sky130_fd_sc_hd__o2111a_1 _6437_ (.A1(_2790_),
    .A2(_2868_),
    .B1(_2801_),
    .C1(_2787_),
    .D1(_2864_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2869_));
 sky130_fd_sc_hd__o21a_1 _6438_ (.A1(\i_tinyqv.mem.q_ctrl.delay_cycles_cfg[2] ),
    .A2(\i_tinyqv.mem.q_ctrl.delay_cycles_cfg[1] ),
    .B1(_2788_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2870_));
 sky130_fd_sc_hd__or4b_1 _6439_ (.A(_2853_),
    .B(_2869_),
    .C(_2870_),
    .D_N(_2863_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2871_));
 sky130_fd_sc_hd__o211a_1 _6440_ (.A1(\i_tinyqv.mem.q_ctrl.fsm_state[1] ),
    .A2(_2863_),
    .B1(_2871_),
    .C1(_2832_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0401_));
 sky130_fd_sc_hd__o41a_1 _6441_ (.A1(_1706_),
    .A2(_2846_),
    .A3(_2795_),
    .A4(_2867_),
    .B1(_1540_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2872_));
 sky130_fd_sc_hd__mux2_1 _6442_ (.A0(_1706_),
    .A1(_2872_),
    .S(_2863_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2873_));
 sky130_fd_sc_hd__and2_1 _6443_ (.A(_2832_),
    .B(_2873_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2874_));
 sky130_fd_sc_hd__clkbuf_1 _6444_ (.A(_2874_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0402_));
 sky130_fd_sc_hd__o21ai_1 _6445_ (.A1(_2801_),
    .A2(_2825_),
    .B1(_2787_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2875_));
 sky130_fd_sc_hd__and4_1 _6446_ (.A(_2792_),
    .B(_2811_),
    .C(_2806_),
    .D(_2875_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2876_));
 sky130_fd_sc_hd__clkbuf_1 _6447_ (.A(_2876_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0403_));
 sky130_fd_sc_hd__clkbuf_4 _6448_ (.A(_2734_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2877_));
 sky130_fd_sc_hd__buf_4 _6449_ (.A(_2877_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2878_));
 sky130_fd_sc_hd__a31o_1 _6450_ (.A1(\i_tinyqv.cpu.data_addr[24] ),
    .A2(\i_tinyqv.cpu.data_addr[23] ),
    .A3(_2878_),
    .B1(_2855_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2879_));
 sky130_fd_sc_hd__nand2_1 _6451_ (.A(_2832_),
    .B(_2879_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2880_));
 sky130_fd_sc_hd__a21o_1 _6452_ (.A1(net210),
    .A2(_2855_),
    .B1(_2880_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0404_));
 sky130_fd_sc_hd__a221o_1 _6453_ (.A1(_2838_),
    .A2(_2840_),
    .B1(_2855_),
    .B2(net208),
    .C1(_2305_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0405_));
 sky130_fd_sc_hd__a211o_1 _6454_ (.A1(net289),
    .A2(_2855_),
    .B1(_2857_),
    .C1(_2305_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0406_));
 sky130_fd_sc_hd__nor2_1 _6455_ (.A(\i_tinyqv.mem.q_ctrl.spi_clk_out ),
    .B(_2836_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2881_));
 sky130_fd_sc_hd__a31o_1 _6456_ (.A1(\i_tinyqv.mem.q_ctrl.spi_clk_out ),
    .A2(_2810_),
    .A3(_2855_),
    .B1(_2881_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2882_));
 sky130_fd_sc_hd__and2_1 _6457_ (.A(_2832_),
    .B(_2882_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2883_));
 sky130_fd_sc_hd__clkbuf_1 _6458_ (.A(_2883_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0407_));
 sky130_fd_sc_hd__a21o_1 _6459_ (.A1(\i_tinyqv.mem.q_ctrl.spi_flash_select ),
    .A2(_2792_),
    .B1(_1708_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2884_));
 sky130_fd_sc_hd__a211o_1 _6460_ (.A1(_2800_),
    .A2(_2884_),
    .B1(_2803_),
    .C1(_2813_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2885_));
 sky130_fd_sc_hd__mux2_1 _6461_ (.A0(_1715_),
    .A1(_2836_),
    .S(_2803_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2886_));
 sky130_fd_sc_hd__a21o_1 _6462_ (.A1(_2885_),
    .A2(_2886_),
    .B1(_2794_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2887_));
 sky130_fd_sc_hd__o211a_1 _6463_ (.A1(_2797_),
    .A2(_2803_),
    .B1(_2842_),
    .C1(_2887_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2888_));
 sky130_fd_sc_hd__o21ai_1 _6464_ (.A1(net145),
    .A2(_2888_),
    .B1(_2832_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2889_));
 sky130_fd_sc_hd__a21oi_1 _6465_ (.A1(_1540_),
    .A2(_2888_),
    .B1(_2889_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0408_));
 sky130_fd_sc_hd__nor2_1 _6466_ (.A(_1181_),
    .B(_2625_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2890_));
 sky130_fd_sc_hd__a211o_1 _6467_ (.A1(_2640_),
    .A2(_2625_),
    .B1(_2890_),
    .C1(_0845_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2891_));
 sky130_fd_sc_hd__o21ai_1 _6468_ (.A1(_1312_),
    .A2(_1124_),
    .B1(_2891_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2892_));
 sky130_fd_sc_hd__a22o_1 _6469_ (.A1(\i_tinyqv.cpu.i_core.i_shift.a[28] ),
    .A2(_2596_),
    .B1(_2629_),
    .B2(_2892_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0409_));
 sky130_fd_sc_hd__nor2_1 _6470_ (.A(_1260_),
    .B(_2625_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2893_));
 sky130_fd_sc_hd__a211o_1 _6471_ (.A1(_2647_),
    .A2(_2625_),
    .B1(_2893_),
    .C1(_0845_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2894_));
 sky130_fd_sc_hd__nand2_1 _6472_ (.A(net66),
    .B(_0845_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2895_));
 sky130_fd_sc_hd__a32o_1 _6473_ (.A1(_2629_),
    .A2(_2894_),
    .A3(_2895_),
    .B1(_2596_),
    .B2(\i_tinyqv.cpu.i_core.i_shift.a[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0410_));
 sky130_fd_sc_hd__or4b_1 _6474_ (.A(_1713_),
    .B(\i_tinyqv.mem.q_ctrl.read_cycles_count[0] ),
    .C(_2787_),
    .D_N(_2782_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2896_));
 sky130_fd_sc_hd__buf_2 _6475_ (.A(_2896_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2897_));
 sky130_fd_sc_hd__mux2_1 _6476_ (.A0(net10),
    .A1(\i_tinyqv.mem.q_ctrl.spi_in_buffer[0] ),
    .S(_2897_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2898_));
 sky130_fd_sc_hd__clkbuf_1 _6477_ (.A(_2898_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0411_));
 sky130_fd_sc_hd__mux2_1 _6478_ (.A0(net11),
    .A1(net133),
    .S(_2897_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2899_));
 sky130_fd_sc_hd__clkbuf_1 _6479_ (.A(_2899_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0412_));
 sky130_fd_sc_hd__mux2_1 _6480_ (.A0(net12),
    .A1(\i_tinyqv.mem.q_ctrl.spi_in_buffer[2] ),
    .S(_2897_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2900_));
 sky130_fd_sc_hd__clkbuf_1 _6481_ (.A(_2900_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0413_));
 sky130_fd_sc_hd__mux2_1 _6482_ (.A0(net13),
    .A1(\i_tinyqv.mem.q_ctrl.spi_in_buffer[3] ),
    .S(_2897_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2901_));
 sky130_fd_sc_hd__clkbuf_1 _6483_ (.A(_2901_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0414_));
 sky130_fd_sc_hd__mux2_1 _6484_ (.A0(net167),
    .A1(\i_tinyqv.mem.q_ctrl.spi_in_buffer[4] ),
    .S(_2897_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2902_));
 sky130_fd_sc_hd__clkbuf_1 _6485_ (.A(net168),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0415_));
 sky130_fd_sc_hd__mux2_1 _6486_ (.A0(net133),
    .A1(\i_tinyqv.mem.q_ctrl.spi_in_buffer[5] ),
    .S(_2897_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2903_));
 sky130_fd_sc_hd__clkbuf_1 _6487_ (.A(net134),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0416_));
 sky130_fd_sc_hd__mux2_1 _6488_ (.A0(\i_tinyqv.mem.q_ctrl.spi_in_buffer[2] ),
    .A1(net271),
    .S(_2897_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2904_));
 sky130_fd_sc_hd__clkbuf_1 _6489_ (.A(_2904_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0417_));
 sky130_fd_sc_hd__mux2_1 _6490_ (.A0(\i_tinyqv.mem.q_ctrl.spi_in_buffer[3] ),
    .A1(net274),
    .S(_2897_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2905_));
 sky130_fd_sc_hd__clkbuf_1 _6491_ (.A(_2905_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0418_));
 sky130_fd_sc_hd__nand2_4 _6492_ (.A(_0868_),
    .B(\i_tinyqv.mem.q_ctrl.data_req ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2906_));
 sky130_fd_sc_hd__or2_1 _6493_ (.A(_0868_),
    .B(\i_tinyqv.mem.q_ctrl.data_req ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2907_));
 sky130_fd_sc_hd__and2_1 _6494_ (.A(_2906_),
    .B(_2907_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2908_));
 sky130_fd_sc_hd__buf_2 _6495_ (.A(_2908_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2909_));
 sky130_fd_sc_hd__mux2_1 _6496_ (.A0(\i_debug_uart_tx.uart_tx_data[0] ),
    .A1(\i_spi.end_txn ),
    .S(_2909_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2910_));
 sky130_fd_sc_hd__nand2_1 _6497_ (.A(_2906_),
    .B(_2907_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2911_));
 sky130_fd_sc_hd__clkbuf_4 _6498_ (.A(_2911_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2912_));
 sky130_fd_sc_hd__mux2_1 _6499_ (.A0(\i_tinyqv.cpu.data_out[24] ),
    .A1(\i_tinyqv.cpu.data_out[16] ),
    .S(_2912_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2913_));
 sky130_fd_sc_hd__xnor2_4 _6500_ (.A(\i_tinyqv.mem.qspi_data_byte_idx[1] ),
    .B(_2906_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2914_));
 sky130_fd_sc_hd__mux2_1 _6501_ (.A0(_2910_),
    .A1(_2913_),
    .S(_2914_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2915_));
 sky130_fd_sc_hd__nand2_2 _6502_ (.A(_2787_),
    .B(_2795_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2916_));
 sky130_fd_sc_hd__mux2_1 _6503_ (.A0(net10),
    .A1(_2915_),
    .S(_2916_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2917_));
 sky130_fd_sc_hd__or4bb_4 _6504_ (.A(\i_tinyqv.mem.q_ctrl.read_cycles_count[0] ),
    .B(\i_tinyqv.mem.q_ctrl.read_cycles_count[2] ),
    .C_N(_2789_),
    .D_N(\i_tinyqv.mem.q_ctrl.read_cycles_count[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2918_));
 sky130_fd_sc_hd__mux2_1 _6505_ (.A0(\i_tinyqv.mem.q_ctrl.spi_in_buffer[4] ),
    .A1(\i_tinyqv.mem.q_ctrl.spi_in_buffer[0] ),
    .S(_2918_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2919_));
 sky130_fd_sc_hd__or3b_2 _6506_ (.A(_2782_),
    .B(\i_tinyqv.mem.q_ctrl.read_cycles_count[0] ),
    .C_N(_1711_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2920_));
 sky130_fd_sc_hd__mux2_1 _6507_ (.A0(net10),
    .A1(_2919_),
    .S(_2920_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2921_));
 sky130_fd_sc_hd__mux2_1 _6508_ (.A0(_2917_),
    .A1(_2921_),
    .S(_2792_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2922_));
 sky130_fd_sc_hd__o21a_1 _6509_ (.A1(_2791_),
    .A2(_2800_),
    .B1(_2918_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2923_));
 sky130_fd_sc_hd__o221a_1 _6510_ (.A1(\i_tinyqv.mem.q_ctrl.spi_clk_out ),
    .A2(_2813_),
    .B1(_2916_),
    .B2(_1711_),
    .C1(_1713_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2924_));
 sky130_fd_sc_hd__o21ba_4 _6511_ (.A1(_1713_),
    .A2(_2923_),
    .B1_N(_2924_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2925_));
 sky130_fd_sc_hd__mux2_1 _6512_ (.A0(_2922_),
    .A1(_2316_),
    .S(_2925_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2926_));
 sky130_fd_sc_hd__clkbuf_1 _6513_ (.A(_2926_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0419_));
 sky130_fd_sc_hd__mux2_1 _6514_ (.A0(\i_tinyqv.cpu.data_out[25] ),
    .A1(\i_tinyqv.cpu.data_out[17] ),
    .S(_2912_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2927_));
 sky130_fd_sc_hd__mux2_1 _6515_ (.A0(\i_debug_uart_tx.uart_tx_data[1] ),
    .A1(\i_spi.dc_in ),
    .S(_2909_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2928_));
 sky130_fd_sc_hd__xnor2_4 _6516_ (.A(_0864_),
    .B(_2906_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2929_));
 sky130_fd_sc_hd__mux2_1 _6517_ (.A0(_2927_),
    .A1(_2928_),
    .S(_2929_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2930_));
 sky130_fd_sc_hd__mux2_1 _6518_ (.A0(net11),
    .A1(_2930_),
    .S(_2916_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2931_));
 sky130_fd_sc_hd__mux2_1 _6519_ (.A0(\i_tinyqv.mem.q_ctrl.spi_in_buffer[5] ),
    .A1(\i_tinyqv.mem.q_ctrl.spi_in_buffer[1] ),
    .S(_2918_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2932_));
 sky130_fd_sc_hd__mux2_1 _6520_ (.A0(net11),
    .A1(_2932_),
    .S(_2920_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2933_));
 sky130_fd_sc_hd__mux2_1 _6521_ (.A0(_2931_),
    .A1(_2933_),
    .S(_2792_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2934_));
 sky130_fd_sc_hd__mux2_1 _6522_ (.A0(_2934_),
    .A1(_2318_),
    .S(_2925_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2935_));
 sky130_fd_sc_hd__clkbuf_1 _6523_ (.A(_2935_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0420_));
 sky130_fd_sc_hd__mux2_1 _6524_ (.A0(\i_debug_uart_tx.uart_tx_data[2] ),
    .A1(\i_tinyqv.cpu.data_out[10] ),
    .S(_2909_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2936_));
 sky130_fd_sc_hd__mux2_1 _6525_ (.A0(\i_tinyqv.cpu.data_out[26] ),
    .A1(\i_tinyqv.cpu.data_out[18] ),
    .S(_2911_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2937_));
 sky130_fd_sc_hd__mux2_1 _6526_ (.A0(_2936_),
    .A1(_2937_),
    .S(_2914_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2938_));
 sky130_fd_sc_hd__mux2_1 _6527_ (.A0(net12),
    .A1(_2938_),
    .S(_2916_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2939_));
 sky130_fd_sc_hd__mux2_1 _6528_ (.A0(\i_tinyqv.mem.q_ctrl.spi_in_buffer[6] ),
    .A1(\i_tinyqv.mem.q_ctrl.spi_in_buffer[2] ),
    .S(_2918_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2940_));
 sky130_fd_sc_hd__mux2_1 _6529_ (.A0(net12),
    .A1(_2940_),
    .S(_2920_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2941_));
 sky130_fd_sc_hd__mux2_1 _6530_ (.A0(_2939_),
    .A1(_2941_),
    .S(_2792_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2942_));
 sky130_fd_sc_hd__mux2_1 _6531_ (.A0(_2942_),
    .A1(_2320_),
    .S(_2925_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2943_));
 sky130_fd_sc_hd__clkbuf_1 _6532_ (.A(_2943_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0421_));
 sky130_fd_sc_hd__mux2_1 _6533_ (.A0(\i_tinyqv.cpu.data_out[27] ),
    .A1(\i_tinyqv.cpu.data_out[19] ),
    .S(_2912_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2944_));
 sky130_fd_sc_hd__mux2_1 _6534_ (.A0(\i_debug_uart_tx.uart_tx_data[3] ),
    .A1(\i_tinyqv.cpu.data_out[11] ),
    .S(_2909_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2945_));
 sky130_fd_sc_hd__mux2_1 _6535_ (.A0(_2944_),
    .A1(_2945_),
    .S(_2929_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2946_));
 sky130_fd_sc_hd__mux2_1 _6536_ (.A0(net13),
    .A1(_2946_),
    .S(_2916_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2947_));
 sky130_fd_sc_hd__mux2_1 _6537_ (.A0(\i_tinyqv.mem.q_ctrl.spi_in_buffer[7] ),
    .A1(\i_tinyqv.mem.q_ctrl.spi_in_buffer[3] ),
    .S(_2918_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2948_));
 sky130_fd_sc_hd__mux2_1 _6538_ (.A0(net13),
    .A1(_2948_),
    .S(_2920_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2949_));
 sky130_fd_sc_hd__mux2_1 _6539_ (.A0(_2947_),
    .A1(_2949_),
    .S(_2792_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2950_));
 sky130_fd_sc_hd__mux2_1 _6540_ (.A0(_2950_),
    .A1(_2322_),
    .S(_2925_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2951_));
 sky130_fd_sc_hd__clkbuf_1 _6541_ (.A(_2951_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0422_));
 sky130_fd_sc_hd__and2_1 _6542_ (.A(_1713_),
    .B(_2916_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2952_));
 sky130_fd_sc_hd__mux2_1 _6543_ (.A0(\i_tinyqv.cpu.data_out[28] ),
    .A1(\i_tinyqv.cpu.data_out[20] ),
    .S(_2912_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2953_));
 sky130_fd_sc_hd__or2_1 _6544_ (.A(\i_debug_uart_tx.uart_tx_data[4] ),
    .B(_2909_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2954_));
 sky130_fd_sc_hd__o211a_1 _6545_ (.A1(\i_tinyqv.cpu.data_out[12] ),
    .A2(_2912_),
    .B1(_2929_),
    .C1(_2954_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2955_));
 sky130_fd_sc_hd__nand2_2 _6546_ (.A(_1713_),
    .B(_2916_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2956_));
 sky130_fd_sc_hd__a211o_1 _6547_ (.A1(_2914_),
    .A2(_2953_),
    .B1(_2955_),
    .C1(_2956_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2957_));
 sky130_fd_sc_hd__o21a_1 _6548_ (.A1(_2316_),
    .A2(_2952_),
    .B1(_2957_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2958_));
 sky130_fd_sc_hd__mux2_1 _6549_ (.A0(_2958_),
    .A1(_1712_),
    .S(_2925_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2959_));
 sky130_fd_sc_hd__clkbuf_1 _6550_ (.A(_2959_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0423_));
 sky130_fd_sc_hd__mux2_1 _6551_ (.A0(\i_tinyqv.cpu.data_out[29] ),
    .A1(\i_tinyqv.cpu.data_out[21] ),
    .S(_2912_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2960_));
 sky130_fd_sc_hd__or2_1 _6552_ (.A(\i_debug_uart_tx.uart_tx_data[5] ),
    .B(_2909_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2961_));
 sky130_fd_sc_hd__o211a_1 _6553_ (.A1(\i_tinyqv.cpu.data_out[13] ),
    .A2(_2912_),
    .B1(_2929_),
    .C1(_2961_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2962_));
 sky130_fd_sc_hd__a211o_1 _6554_ (.A1(_2914_),
    .A2(_2960_),
    .B1(_2962_),
    .C1(_2956_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2963_));
 sky130_fd_sc_hd__o21a_1 _6555_ (.A1(_2318_),
    .A2(_2952_),
    .B1(_2963_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2964_));
 sky130_fd_sc_hd__mux2_1 _6556_ (.A0(_2964_),
    .A1(_1717_),
    .S(_2925_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2965_));
 sky130_fd_sc_hd__clkbuf_1 _6557_ (.A(_2965_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0424_));
 sky130_fd_sc_hd__mux2_1 _6558_ (.A0(\i_debug_uart_tx.uart_tx_data[6] ),
    .A1(\i_tinyqv.cpu.data_out[14] ),
    .S(_2909_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2966_));
 sky130_fd_sc_hd__or2_1 _6559_ (.A(\i_tinyqv.cpu.data_out[30] ),
    .B(_2912_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2967_));
 sky130_fd_sc_hd__o211a_1 _6560_ (.A1(\i_tinyqv.cpu.data_out[22] ),
    .A2(_2909_),
    .B1(_2914_),
    .C1(_2967_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2968_));
 sky130_fd_sc_hd__a211o_1 _6561_ (.A1(_2929_),
    .A2(_2966_),
    .B1(_2968_),
    .C1(_2956_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2969_));
 sky130_fd_sc_hd__o21a_1 _6562_ (.A1(_2320_),
    .A2(_2952_),
    .B1(_2969_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2970_));
 sky130_fd_sc_hd__mux2_1 _6563_ (.A0(_2970_),
    .A1(_1720_),
    .S(_2925_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2971_));
 sky130_fd_sc_hd__clkbuf_1 _6564_ (.A(_2971_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0425_));
 sky130_fd_sc_hd__mux2_1 _6565_ (.A0(\i_tinyqv.cpu.data_out[31] ),
    .A1(\i_tinyqv.cpu.data_out[23] ),
    .S(_2912_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2972_));
 sky130_fd_sc_hd__or2_1 _6566_ (.A(\i_debug_uart_tx.uart_tx_data[7] ),
    .B(_2909_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2973_));
 sky130_fd_sc_hd__o211a_1 _6567_ (.A1(\i_tinyqv.cpu.data_out[15] ),
    .A2(_2912_),
    .B1(_2929_),
    .C1(_2973_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2974_));
 sky130_fd_sc_hd__a211o_1 _6568_ (.A1(_2914_),
    .A2(_2972_),
    .B1(_2974_),
    .C1(_2956_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2975_));
 sky130_fd_sc_hd__o21a_1 _6569_ (.A1(_2322_),
    .A2(_2952_),
    .B1(_2975_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2976_));
 sky130_fd_sc_hd__mux2_1 _6570_ (.A0(_2976_),
    .A1(_1721_),
    .S(_2925_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2977_));
 sky130_fd_sc_hd__clkbuf_1 _6571_ (.A(_2977_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0426_));
 sky130_fd_sc_hd__or2_1 _6572_ (.A(net311),
    .B(_2229_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2978_));
 sky130_fd_sc_hd__clkbuf_1 _6573_ (.A(_2978_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0427_));
 sky130_fd_sc_hd__or2_1 _6574_ (.A(\i_tinyqv.mem.q_ctrl.spi_ram_a_select ),
    .B(_2229_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2979_));
 sky130_fd_sc_hd__clkbuf_1 _6575_ (.A(_2979_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0428_));
 sky130_fd_sc_hd__nor2_1 _6576_ (.A(_2229_),
    .B(_1543_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0429_));
 sky130_fd_sc_hd__or2_1 _6577_ (.A(_1400_),
    .B(\i_tinyqv.cpu.instr_data[2][0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2980_));
 sky130_fd_sc_hd__mux2_1 _6578_ (.A0(\i_tinyqv.cpu.instr_data_in[0] ),
    .A1(_2980_),
    .S(_2562_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2981_));
 sky130_fd_sc_hd__clkbuf_1 _6579_ (.A(_2981_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0430_));
 sky130_fd_sc_hd__or2_1 _6580_ (.A(_1400_),
    .B(\i_tinyqv.cpu.instr_data[2][1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2982_));
 sky130_fd_sc_hd__mux2_1 _6581_ (.A0(\i_tinyqv.cpu.instr_data_in[1] ),
    .A1(_2982_),
    .S(_2562_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2983_));
 sky130_fd_sc_hd__clkbuf_1 _6582_ (.A(_2983_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0431_));
 sky130_fd_sc_hd__mux2_1 _6583_ (.A0(net10),
    .A1(\i_tinyqv.mem.q_ctrl.delay_cycles_cfg[0] ),
    .S(_1737_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2984_));
 sky130_fd_sc_hd__clkbuf_1 _6584_ (.A(_2984_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0432_));
 sky130_fd_sc_hd__mux2_1 _6585_ (.A0(net11),
    .A1(\i_tinyqv.mem.q_ctrl.delay_cycles_cfg[1] ),
    .S(_1728_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2985_));
 sky130_fd_sc_hd__clkbuf_1 _6586_ (.A(_2985_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0433_));
 sky130_fd_sc_hd__mux2_1 _6587_ (.A0(net12),
    .A1(\i_tinyqv.mem.q_ctrl.delay_cycles_cfg[2] ),
    .S(_1728_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2986_));
 sky130_fd_sc_hd__clkbuf_1 _6588_ (.A(_2986_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0434_));
 sky130_fd_sc_hd__clkbuf_4 _6589_ (.A(net31),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2987_));
 sky130_fd_sc_hd__xor2_1 _6590_ (.A(_0749_),
    .B(\i_tinyqv.cpu.i_core.imm_lo[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2988_));
 sky130_fd_sc_hd__and2_1 _6591_ (.A(_0653_),
    .B(\i_tinyqv.cpu.is_branch ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2989_));
 sky130_fd_sc_hd__clkbuf_4 _6592_ (.A(_2989_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2990_));
 sky130_fd_sc_hd__buf_4 _6593_ (.A(_2990_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2991_));
 sky130_fd_sc_hd__mux2_1 _6594_ (.A0(_2505_),
    .A1(_2988_),
    .S(_2991_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2992_));
 sky130_fd_sc_hd__clkbuf_4 _6595_ (.A(net40),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2993_));
 sky130_fd_sc_hd__a22o_1 _6596_ (.A1(\i_tinyqv.cpu.i_core.i_registers.registers[1][9] ),
    .A2(_2987_),
    .B1(_2992_),
    .B2(_2993_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2994_));
 sky130_fd_sc_hd__clkbuf_4 _6597_ (.A(_2306_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2995_));
 sky130_fd_sc_hd__and2b_1 _6598_ (.A_N(_1521_),
    .B(_2995_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2996_));
 sky130_fd_sc_hd__o21a_1 _6599_ (.A1(_2994_),
    .A2(_2996_),
    .B1(_2061_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0435_));
 sky130_fd_sc_hd__xor2_1 _6600_ (.A(net85),
    .B(\i_tinyqv.cpu.i_core.imm_lo[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2997_));
 sky130_fd_sc_hd__and3_1 _6601_ (.A(_0749_),
    .B(\i_tinyqv.cpu.i_core.imm_lo[1] ),
    .C(_2997_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_2998_));
 sky130_fd_sc_hd__a21oi_1 _6602_ (.A1(_0749_),
    .A2(\i_tinyqv.cpu.i_core.imm_lo[1] ),
    .B1(_2997_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_2999_));
 sky130_fd_sc_hd__nor2_1 _6603_ (.A(_2998_),
    .B(_2999_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3000_));
 sky130_fd_sc_hd__mux2_1 _6604_ (.A0(_2507_),
    .A1(_3000_),
    .S(_2991_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3001_));
 sky130_fd_sc_hd__a22o_1 _6605_ (.A1(\i_tinyqv.cpu.i_core.i_registers.registers[1][10] ),
    .A2(_2987_),
    .B1(_3001_),
    .B2(_2993_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3002_));
 sky130_fd_sc_hd__and2b_1 _6606_ (.A_N(_1524_),
    .B(_2995_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3003_));
 sky130_fd_sc_hd__o21a_1 _6607_ (.A1(_3002_),
    .A2(_3003_),
    .B1(_2061_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0436_));
 sky130_fd_sc_hd__a21oi_4 _6608_ (.A1(_1551_),
    .A2(_1536_),
    .B1(_1541_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3004_));
 sky130_fd_sc_hd__clkbuf_4 _6609_ (.A(_3004_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3005_));
 sky130_fd_sc_hd__and2_2 _6610_ (.A(\i_tinyqv.mem.q_ctrl.spi_clk_out ),
    .B(_1709_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3006_));
 sky130_fd_sc_hd__clkbuf_4 _6611_ (.A(_3006_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3007_));
 sky130_fd_sc_hd__nor2_1 _6612_ (.A(_3004_),
    .B(_3007_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3008_));
 sky130_fd_sc_hd__clkbuf_4 _6613_ (.A(_3008_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3009_));
 sky130_fd_sc_hd__a32o_1 _6614_ (.A1(net300),
    .A2(_2878_),
    .A3(_3005_),
    .B1(_3009_),
    .B2(net122),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0437_));
 sky130_fd_sc_hd__clkbuf_4 _6615_ (.A(\i_tinyqv.cpu.was_early_branch ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3010_));
 sky130_fd_sc_hd__mux2_1 _6616_ (.A0(_1406_),
    .A1(_2988_),
    .S(_3010_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3011_));
 sky130_fd_sc_hd__clkbuf_4 _6617_ (.A(_2681_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3012_));
 sky130_fd_sc_hd__mux2_1 _6618_ (.A0(\i_tinyqv.cpu.data_addr[1] ),
    .A1(_3011_),
    .S(_3012_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3013_));
 sky130_fd_sc_hd__a22o_1 _6619_ (.A1(net93),
    .A2(_3009_),
    .B1(_3013_),
    .B2(_3005_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0438_));
 sky130_fd_sc_hd__mux2_1 _6620_ (.A0(\i_tinyqv.cpu.instr_write_offset[2] ),
    .A1(_3000_),
    .S(_3010_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3014_));
 sky130_fd_sc_hd__mux2_1 _6621_ (.A0(\i_tinyqv.cpu.data_addr[2] ),
    .A1(_3014_),
    .S(_3012_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3015_));
 sky130_fd_sc_hd__a22o_1 _6622_ (.A1(net126),
    .A2(_3009_),
    .B1(_3015_),
    .B2(_3005_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0439_));
 sky130_fd_sc_hd__or2_1 _6623_ (.A(_0884_),
    .B(\i_tinyqv.cpu.instr_write_offset[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3016_));
 sky130_fd_sc_hd__clkbuf_4 _6624_ (.A(\i_tinyqv.cpu.was_early_branch ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3017_));
 sky130_fd_sc_hd__a21oi_1 _6625_ (.A1(_0884_),
    .A2(\i_tinyqv.cpu.instr_write_offset[3] ),
    .B1(_3017_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3018_));
 sky130_fd_sc_hd__nand2_1 _6626_ (.A(\i_tinyqv.cpu.instr_data_start[3] ),
    .B(\i_tinyqv.cpu.i_core.imm_lo[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3019_));
 sky130_fd_sc_hd__or2_1 _6627_ (.A(\i_tinyqv.cpu.instr_data_start[3] ),
    .B(\i_tinyqv.cpu.i_core.imm_lo[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3020_));
 sky130_fd_sc_hd__nand2_1 _6628_ (.A(_3019_),
    .B(_3020_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3021_));
 sky130_fd_sc_hd__a21oi_1 _6629_ (.A1(net60),
    .A2(\i_tinyqv.cpu.i_core.imm_lo[2] ),
    .B1(_2998_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3022_));
 sky130_fd_sc_hd__xor2_1 _6630_ (.A(_3021_),
    .B(_3022_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3023_));
 sky130_fd_sc_hd__a221o_1 _6631_ (.A1(_3016_),
    .A2(_3018_),
    .B1(_3023_),
    .B2(_3017_),
    .C1(_2878_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3024_));
 sky130_fd_sc_hd__or2_1 _6632_ (.A(\i_tinyqv.cpu.data_addr[3] ),
    .B(_3012_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3025_));
 sky130_fd_sc_hd__a32o_1 _6633_ (.A1(_3005_),
    .A2(_3024_),
    .A3(_3025_),
    .B1(_3009_),
    .B2(net95),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0440_));
 sky130_fd_sc_hd__nand2_1 _6634_ (.A(_1442_),
    .B(_2306_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3026_));
 sky130_fd_sc_hd__clkbuf_4 _6635_ (.A(_3026_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3027_));
 sky130_fd_sc_hd__and2_1 _6636_ (.A(_1442_),
    .B(_2306_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3028_));
 sky130_fd_sc_hd__clkbuf_4 _6637_ (.A(_3028_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3029_));
 sky130_fd_sc_hd__a211o_1 _6638_ (.A1(_1415_),
    .A2(_2995_),
    .B1(_2994_),
    .C1(_3029_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3030_));
 sky130_fd_sc_hd__o211a_1 _6639_ (.A1(_0749_),
    .A2(_3027_),
    .B1(_3030_),
    .C1(_2061_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0441_));
 sky130_fd_sc_hd__a211o_1 _6640_ (.A1(_1339_),
    .A2(_2995_),
    .B1(_3002_),
    .C1(_3029_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3031_));
 sky130_fd_sc_hd__o211a_1 _6641_ (.A1(net60),
    .A2(_3027_),
    .B1(_3031_),
    .C1(_2061_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0442_));
 sky130_fd_sc_hd__mux2_1 _6642_ (.A0(\i_spi.end_txn ),
    .A1(net308),
    .S(_2415_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3032_));
 sky130_fd_sc_hd__clkbuf_1 _6643_ (.A(_3032_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0443_));
 sky130_fd_sc_hd__mux2_1 _6644_ (.A0(_1591_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.registers[1][11] ),
    .S(net31),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3033_));
 sky130_fd_sc_hd__mux2_1 _6645_ (.A0(_2509_),
    .A1(_3023_),
    .S(_2991_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3034_));
 sky130_fd_sc_hd__mux2_1 _6646_ (.A0(_3033_),
    .A1(_3034_),
    .S(_2993_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3035_));
 sky130_fd_sc_hd__or2_1 _6647_ (.A(_3029_),
    .B(_3035_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3036_));
 sky130_fd_sc_hd__o211a_1 _6648_ (.A1(_0884_),
    .A2(_3027_),
    .B1(_3036_),
    .C1(_2061_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0444_));
 sky130_fd_sc_hd__buf_2 _6649_ (.A(_3026_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3037_));
 sky130_fd_sc_hd__inv_2 _6650_ (.A(\i_tinyqv.cpu.i_core.i_registers.registers[1][12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3038_));
 sky130_fd_sc_hd__clkbuf_4 _6651_ (.A(_2987_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3039_));
 sky130_fd_sc_hd__clkbuf_4 _6652_ (.A(_1390_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3040_));
 sky130_fd_sc_hd__nand2_1 _6653_ (.A(\i_tinyqv.cpu.instr_data_start[4] ),
    .B(\i_tinyqv.cpu.i_core.imm_lo[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3041_));
 sky130_fd_sc_hd__or2_1 _6654_ (.A(\i_tinyqv.cpu.instr_data_start[4] ),
    .B(\i_tinyqv.cpu.i_core.imm_lo[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3042_));
 sky130_fd_sc_hd__nand2_1 _6655_ (.A(_3041_),
    .B(_3042_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3043_));
 sky130_fd_sc_hd__o21a_1 _6656_ (.A1(_3021_),
    .A2(_3022_),
    .B1(_3019_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3044_));
 sky130_fd_sc_hd__xnor2_2 _6657_ (.A(_3043_),
    .B(_3044_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3045_));
 sky130_fd_sc_hd__nand2_1 _6658_ (.A(_1390_),
    .B(_2511_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3046_));
 sky130_fd_sc_hd__clkbuf_4 _6659_ (.A(net40),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3047_));
 sky130_fd_sc_hd__o211a_1 _6660_ (.A1(_3040_),
    .A2(_3045_),
    .B1(_3046_),
    .C1(_3047_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3048_));
 sky130_fd_sc_hd__a221o_1 _6661_ (.A1(_3038_),
    .A2(_3039_),
    .B1(_2995_),
    .B2(_0905_),
    .C1(_3048_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3049_));
 sky130_fd_sc_hd__nand2_1 _6662_ (.A(_3037_),
    .B(_3049_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3050_));
 sky130_fd_sc_hd__o211a_1 _6663_ (.A1(\i_tinyqv.cpu.instr_data_start[4] ),
    .A2(_3027_),
    .B1(_3050_),
    .C1(_2061_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0445_));
 sky130_fd_sc_hd__clkbuf_4 _6664_ (.A(_2993_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3051_));
 sky130_fd_sc_hd__and2_1 _6665_ (.A(\i_tinyqv.cpu.instr_data_start[5] ),
    .B(\i_tinyqv.cpu.i_core.imm_lo[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3052_));
 sky130_fd_sc_hd__nor2_1 _6666_ (.A(\i_tinyqv.cpu.instr_data_start[5] ),
    .B(\i_tinyqv.cpu.i_core.imm_lo[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3053_));
 sky130_fd_sc_hd__nor2_1 _6667_ (.A(_3052_),
    .B(_3053_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3054_));
 sky130_fd_sc_hd__o21a_1 _6668_ (.A1(_3043_),
    .A2(_3044_),
    .B1(_3041_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3055_));
 sky130_fd_sc_hd__xnor2_1 _6669_ (.A(_3054_),
    .B(_3055_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3056_));
 sky130_fd_sc_hd__mux2_1 _6670_ (.A0(_2513_),
    .A1(_3056_),
    .S(_2991_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3057_));
 sky130_fd_sc_hd__inv_2 _6671_ (.A(\i_tinyqv.cpu.i_core.i_registers.registers[1][13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3058_));
 sky130_fd_sc_hd__mux2_1 _6672_ (.A0(_1205_),
    .A1(_3058_),
    .S(_2987_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3059_));
 sky130_fd_sc_hd__nor2_1 _6673_ (.A(_3051_),
    .B(_3059_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3060_));
 sky130_fd_sc_hd__a211o_1 _6674_ (.A1(_3051_),
    .A2(_3057_),
    .B1(_3060_),
    .C1(_3029_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3061_));
 sky130_fd_sc_hd__o211a_1 _6675_ (.A1(\i_tinyqv.cpu.instr_data_start[5] ),
    .A2(_3027_),
    .B1(_3061_),
    .C1(_2061_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0446_));
 sky130_fd_sc_hd__inv_2 _6676_ (.A(\i_tinyqv.cpu.i_core.i_registers.registers[1][14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3062_));
 sky130_fd_sc_hd__nand2_1 _6677_ (.A(_0883_),
    .B(\i_tinyqv.cpu.i_core.imm_lo[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3063_));
 sky130_fd_sc_hd__or2_1 _6678_ (.A(_0883_),
    .B(\i_tinyqv.cpu.i_core.imm_lo[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3064_));
 sky130_fd_sc_hd__nand2_1 _6679_ (.A(_3063_),
    .B(_3064_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3065_));
 sky130_fd_sc_hd__o21ba_1 _6680_ (.A1(_3053_),
    .A2(_3055_),
    .B1_N(_3052_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3066_));
 sky130_fd_sc_hd__xnor2_1 _6681_ (.A(_3065_),
    .B(_3066_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3067_));
 sky130_fd_sc_hd__nand2_1 _6682_ (.A(_1390_),
    .B(_2515_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3068_));
 sky130_fd_sc_hd__o211a_1 _6683_ (.A1(_3040_),
    .A2(_3067_),
    .B1(_3068_),
    .C1(_3047_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3069_));
 sky130_fd_sc_hd__a221o_1 _6684_ (.A1(_3062_),
    .A2(_3039_),
    .B1(_2995_),
    .B2(_1340_),
    .C1(_3069_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3070_));
 sky130_fd_sc_hd__nand2_1 _6685_ (.A(_3037_),
    .B(_3070_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3071_));
 sky130_fd_sc_hd__o211a_1 _6686_ (.A1(_0883_),
    .A2(_3027_),
    .B1(_3071_),
    .C1(_2061_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0447_));
 sky130_fd_sc_hd__inv_2 _6687_ (.A(\i_tinyqv.cpu.i_core.i_registers.registers[1][15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3072_));
 sky130_fd_sc_hd__mux2_1 _6688_ (.A0(_1593_),
    .A1(_3072_),
    .S(_2987_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3073_));
 sky130_fd_sc_hd__nor2_1 _6689_ (.A(_3051_),
    .B(_3073_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3074_));
 sky130_fd_sc_hd__or2_1 _6690_ (.A(_2991_),
    .B(_2517_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3075_));
 sky130_fd_sc_hd__nand2_1 _6691_ (.A(\i_tinyqv.cpu.instr_data_start[7] ),
    .B(\i_tinyqv.cpu.i_core.imm_lo[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3076_));
 sky130_fd_sc_hd__or2_1 _6692_ (.A(\i_tinyqv.cpu.instr_data_start[7] ),
    .B(\i_tinyqv.cpu.i_core.imm_lo[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3077_));
 sky130_fd_sc_hd__nand2_1 _6693_ (.A(_3076_),
    .B(_3077_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3078_));
 sky130_fd_sc_hd__o21ai_1 _6694_ (.A1(_3065_),
    .A2(_3066_),
    .B1(_3063_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3079_));
 sky130_fd_sc_hd__xor2_1 _6695_ (.A(_3078_),
    .B(_3079_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3080_));
 sky130_fd_sc_hd__nand2_1 _6696_ (.A(_2991_),
    .B(_3080_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3081_));
 sky130_fd_sc_hd__a31o_1 _6697_ (.A1(_3051_),
    .A2(_3075_),
    .A3(_3081_),
    .B1(_3028_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3082_));
 sky130_fd_sc_hd__o221a_1 _6698_ (.A1(\i_tinyqv.cpu.instr_data_start[7] ),
    .A2(_3037_),
    .B1(_3074_),
    .B2(_3082_),
    .C1(_1753_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0448_));
 sky130_fd_sc_hd__inv_2 _6699_ (.A(\i_tinyqv.cpu.i_core.i_registers.registers[1][16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3083_));
 sky130_fd_sc_hd__nand2_1 _6700_ (.A(\i_tinyqv.cpu.instr_data_start[8] ),
    .B(\i_tinyqv.cpu.i_core.imm_lo[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3084_));
 sky130_fd_sc_hd__or2_1 _6701_ (.A(\i_tinyqv.cpu.instr_data_start[8] ),
    .B(\i_tinyqv.cpu.i_core.imm_lo[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3085_));
 sky130_fd_sc_hd__nand2_1 _6702_ (.A(_3084_),
    .B(_3085_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3086_));
 sky130_fd_sc_hd__a21bo_1 _6703_ (.A1(_3077_),
    .A2(_3079_),
    .B1_N(_3076_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3087_));
 sky130_fd_sc_hd__xnor2_1 _6704_ (.A(_3086_),
    .B(_3087_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3088_));
 sky130_fd_sc_hd__mux2_1 _6705_ (.A0(_2519_),
    .A1(_3088_),
    .S(_2990_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3089_));
 sky130_fd_sc_hd__and2b_1 _6706_ (.A_N(_3089_),
    .B(net40),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3090_));
 sky130_fd_sc_hd__a221o_1 _6707_ (.A1(_3083_),
    .A2(_3039_),
    .B1(_2995_),
    .B2(_0911_),
    .C1(_3090_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3091_));
 sky130_fd_sc_hd__nand2_1 _6708_ (.A(_3037_),
    .B(_3091_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3092_));
 sky130_fd_sc_hd__clkbuf_4 _6709_ (.A(_1752_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3093_));
 sky130_fd_sc_hd__o211a_1 _6710_ (.A1(\i_tinyqv.cpu.instr_data_start[8] ),
    .A2(_3027_),
    .B1(_3092_),
    .C1(_3093_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0449_));
 sky130_fd_sc_hd__mux2_1 _6711_ (.A0(_1202_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.registers[1][17] ),
    .S(net31),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3094_));
 sky130_fd_sc_hd__a21boi_2 _6712_ (.A1(_3085_),
    .A2(_3087_),
    .B1_N(_3084_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3095_));
 sky130_fd_sc_hd__nand2_1 _6713_ (.A(_0882_),
    .B(\i_tinyqv.cpu.i_core.imm_lo[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3096_));
 sky130_fd_sc_hd__or2_1 _6714_ (.A(_0882_),
    .B(\i_tinyqv.cpu.i_core.imm_lo[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3097_));
 sky130_fd_sc_hd__nand2_1 _6715_ (.A(_3096_),
    .B(_3097_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3098_));
 sky130_fd_sc_hd__xor2_1 _6716_ (.A(_3095_),
    .B(_3098_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3099_));
 sky130_fd_sc_hd__mux2_1 _6717_ (.A0(_2521_),
    .A1(_3099_),
    .S(_2990_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3100_));
 sky130_fd_sc_hd__mux2_1 _6718_ (.A0(_3094_),
    .A1(_3100_),
    .S(_2993_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3101_));
 sky130_fd_sc_hd__or2_1 _6719_ (.A(_3029_),
    .B(_3101_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3102_));
 sky130_fd_sc_hd__o211a_1 _6720_ (.A1(_0882_),
    .A2(_3027_),
    .B1(_3102_),
    .C1(_3093_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0450_));
 sky130_fd_sc_hd__inv_2 _6721_ (.A(\i_tinyqv.cpu.i_core.i_registers.registers[1][18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3103_));
 sky130_fd_sc_hd__o21a_1 _6722_ (.A1(_3095_),
    .A2(_3098_),
    .B1(_3096_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3104_));
 sky130_fd_sc_hd__nor2_1 _6723_ (.A(\i_tinyqv.cpu.instr_data_start[10] ),
    .B(\i_tinyqv.cpu.i_core.imm_lo[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3105_));
 sky130_fd_sc_hd__nand2_1 _6724_ (.A(\i_tinyqv.cpu.instr_data_start[10] ),
    .B(\i_tinyqv.cpu.i_core.imm_lo[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3106_));
 sky130_fd_sc_hd__and2b_1 _6725_ (.A_N(_3105_),
    .B(_3106_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3107_));
 sky130_fd_sc_hd__xor2_1 _6726_ (.A(_3104_),
    .B(_3107_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3108_));
 sky130_fd_sc_hd__nand2_1 _6727_ (.A(_1390_),
    .B(_2523_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3109_));
 sky130_fd_sc_hd__o211a_1 _6728_ (.A1(_3040_),
    .A2(_3108_),
    .B1(_3109_),
    .C1(_3047_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3110_));
 sky130_fd_sc_hd__a221o_1 _6729_ (.A1(_3103_),
    .A2(_3039_),
    .B1(_2995_),
    .B2(_1342_),
    .C1(_3110_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3111_));
 sky130_fd_sc_hd__nand2_1 _6730_ (.A(_3037_),
    .B(_3111_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3112_));
 sky130_fd_sc_hd__o211a_1 _6731_ (.A1(\i_tinyqv.cpu.instr_data_start[10] ),
    .A2(_3027_),
    .B1(_3112_),
    .C1(_3093_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0451_));
 sky130_fd_sc_hd__mux2_1 _6732_ (.A0(_1596_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.registers[1][19] ),
    .S(net31),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3113_));
 sky130_fd_sc_hd__nand2_1 _6733_ (.A(\i_tinyqv.cpu.instr_data_start[11] ),
    .B(\i_tinyqv.cpu.i_core.imm_lo[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3114_));
 sky130_fd_sc_hd__or2_1 _6734_ (.A(\i_tinyqv.cpu.instr_data_start[11] ),
    .B(\i_tinyqv.cpu.i_core.imm_lo[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3115_));
 sky130_fd_sc_hd__nand2_1 _6735_ (.A(_3114_),
    .B(_3115_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3116_));
 sky130_fd_sc_hd__o211a_1 _6736_ (.A1(_3095_),
    .A2(_3098_),
    .B1(_3106_),
    .C1(_3096_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3117_));
 sky130_fd_sc_hd__nor2_1 _6737_ (.A(_3105_),
    .B(_3117_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3118_));
 sky130_fd_sc_hd__xnor2_1 _6738_ (.A(_3116_),
    .B(_3118_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3119_));
 sky130_fd_sc_hd__mux2_1 _6739_ (.A0(_2526_),
    .A1(_3119_),
    .S(_2990_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3120_));
 sky130_fd_sc_hd__mux2_1 _6740_ (.A0(_3113_),
    .A1(_3120_),
    .S(_3047_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3121_));
 sky130_fd_sc_hd__or2_1 _6741_ (.A(_3029_),
    .B(_3121_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3122_));
 sky130_fd_sc_hd__o211a_1 _6742_ (.A1(\i_tinyqv.cpu.instr_data_start[11] ),
    .A2(_3027_),
    .B1(_3122_),
    .C1(_3093_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0452_));
 sky130_fd_sc_hd__buf_2 _6743_ (.A(_3026_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3123_));
 sky130_fd_sc_hd__inv_2 _6744_ (.A(\i_tinyqv.cpu.i_core.i_registers.registers[1][20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3124_));
 sky130_fd_sc_hd__o31a_1 _6745_ (.A1(_3116_),
    .A2(_3105_),
    .A3(_3117_),
    .B1(_3114_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3125_));
 sky130_fd_sc_hd__nor2_1 _6746_ (.A(_0726_),
    .B(\i_tinyqv.cpu.imm[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3126_));
 sky130_fd_sc_hd__nand2_1 _6747_ (.A(_0726_),
    .B(\i_tinyqv.cpu.imm[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3127_));
 sky130_fd_sc_hd__or2b_1 _6748_ (.A(_3126_),
    .B_N(_3127_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3128_));
 sky130_fd_sc_hd__xnor2_1 _6749_ (.A(_3125_),
    .B(_3128_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3129_));
 sky130_fd_sc_hd__nand2_1 _6750_ (.A(_1390_),
    .B(_2528_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3130_));
 sky130_fd_sc_hd__o211a_1 _6751_ (.A1(_3040_),
    .A2(_3129_),
    .B1(_3130_),
    .C1(_3047_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3131_));
 sky130_fd_sc_hd__a221o_1 _6752_ (.A1(_3124_),
    .A2(_3039_),
    .B1(_2306_),
    .B2(_0906_),
    .C1(_3131_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3132_));
 sky130_fd_sc_hd__nand2_1 _6753_ (.A(_3037_),
    .B(_3132_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3133_));
 sky130_fd_sc_hd__o211a_1 _6754_ (.A1(_0726_),
    .A2(_3123_),
    .B1(_3133_),
    .C1(_3093_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0453_));
 sky130_fd_sc_hd__nand2_1 _6755_ (.A(\i_tinyqv.cpu.i_core.i_registers.registers[1][21] ),
    .B(net31),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3134_));
 sky130_fd_sc_hd__o21ai_1 _6756_ (.A1(_1201_),
    .A2(_2987_),
    .B1(_3134_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3135_));
 sky130_fd_sc_hd__nand2_1 _6757_ (.A(\i_tinyqv.cpu.instr_data_start[13] ),
    .B(\i_tinyqv.cpu.imm[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3136_));
 sky130_fd_sc_hd__or2_1 _6758_ (.A(\i_tinyqv.cpu.instr_data_start[13] ),
    .B(\i_tinyqv.cpu.imm[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3137_));
 sky130_fd_sc_hd__nand2_1 _6759_ (.A(_3136_),
    .B(_3137_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3138_));
 sky130_fd_sc_hd__o311a_1 _6760_ (.A1(_3116_),
    .A2(_3105_),
    .A3(_3117_),
    .B1(_3114_),
    .C1(_3127_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3139_));
 sky130_fd_sc_hd__nor2_1 _6761_ (.A(_3126_),
    .B(_3139_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3140_));
 sky130_fd_sc_hd__xnor2_1 _6762_ (.A(_3138_),
    .B(_3140_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3141_));
 sky130_fd_sc_hd__mux2_1 _6763_ (.A0(_2530_),
    .A1(_3141_),
    .S(_2990_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3142_));
 sky130_fd_sc_hd__mux2_1 _6764_ (.A0(_3135_),
    .A1(_3142_),
    .S(_3047_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3143_));
 sky130_fd_sc_hd__or2_1 _6765_ (.A(_3029_),
    .B(_3143_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3144_));
 sky130_fd_sc_hd__o211a_1 _6766_ (.A1(\i_tinyqv.cpu.instr_data_start[13] ),
    .A2(_3123_),
    .B1(_3144_),
    .C1(_3093_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0454_));
 sky130_fd_sc_hd__and2_1 _6767_ (.A(_1338_),
    .B(_2995_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3145_));
 sky130_fd_sc_hd__o31a_1 _6768_ (.A1(_3138_),
    .A2(_3126_),
    .A3(_3139_),
    .B1(_3136_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3146_));
 sky130_fd_sc_hd__nor2_1 _6769_ (.A(\i_tinyqv.cpu.instr_data_start[14] ),
    .B(\i_tinyqv.cpu.imm[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3147_));
 sky130_fd_sc_hd__nand2_1 _6770_ (.A(\i_tinyqv.cpu.instr_data_start[14] ),
    .B(\i_tinyqv.cpu.imm[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3148_));
 sky130_fd_sc_hd__and2b_1 _6771_ (.A_N(_3147_),
    .B(_3148_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3149_));
 sky130_fd_sc_hd__xnor2_1 _6772_ (.A(_3146_),
    .B(_3149_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3150_));
 sky130_fd_sc_hd__mux2_1 _6773_ (.A0(_2532_),
    .A1(_3150_),
    .S(_2991_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3151_));
 sky130_fd_sc_hd__a221o_1 _6774_ (.A1(\i_tinyqv.cpu.i_core.i_registers.registers[1][22] ),
    .A2(_3039_),
    .B1(_3151_),
    .B2(_3051_),
    .C1(_3028_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3152_));
 sky130_fd_sc_hd__o221a_1 _6775_ (.A1(\i_tinyqv.cpu.instr_data_start[14] ),
    .A2(_3037_),
    .B1(_3145_),
    .B2(_3152_),
    .C1(_1753_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0455_));
 sky130_fd_sc_hd__nand2_1 _6776_ (.A(_0881_),
    .B(\i_tinyqv.cpu.imm[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3153_));
 sky130_fd_sc_hd__or2_1 _6777_ (.A(_0881_),
    .B(\i_tinyqv.cpu.imm[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3154_));
 sky130_fd_sc_hd__nand2_1 _6778_ (.A(_3153_),
    .B(_3154_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3155_));
 sky130_fd_sc_hd__and2_1 _6779_ (.A(_3148_),
    .B(_3146_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3156_));
 sky130_fd_sc_hd__nor2_1 _6780_ (.A(_3147_),
    .B(_3156_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3157_));
 sky130_fd_sc_hd__xnor2_1 _6781_ (.A(_3155_),
    .B(_3157_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3158_));
 sky130_fd_sc_hd__mux2_1 _6782_ (.A0(_2534_),
    .A1(_3158_),
    .S(_2991_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3159_));
 sky130_fd_sc_hd__inv_2 _6783_ (.A(\i_tinyqv.cpu.i_core.i_registers.registers[1][23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3160_));
 sky130_fd_sc_hd__mux2_1 _6784_ (.A0(_1590_),
    .A1(_3160_),
    .S(_2987_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3161_));
 sky130_fd_sc_hd__nor2_1 _6785_ (.A(_2993_),
    .B(_3161_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3162_));
 sky130_fd_sc_hd__a211o_1 _6786_ (.A1(_3051_),
    .A2(_3159_),
    .B1(_3162_),
    .C1(_3029_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3163_));
 sky130_fd_sc_hd__o211a_1 _6787_ (.A1(_0881_),
    .A2(_3123_),
    .B1(_3163_),
    .C1(_3093_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0456_));
 sky130_fd_sc_hd__inv_2 _6788_ (.A(net105),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3164_));
 sky130_fd_sc_hd__o31a_1 _6789_ (.A1(_3155_),
    .A2(_3147_),
    .A3(_3156_),
    .B1(_3153_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3165_));
 sky130_fd_sc_hd__or2_1 _6790_ (.A(\i_tinyqv.cpu.instr_data_start[16] ),
    .B(\i_tinyqv.cpu.imm[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3166_));
 sky130_fd_sc_hd__nand2_1 _6791_ (.A(\i_tinyqv.cpu.instr_data_start[16] ),
    .B(\i_tinyqv.cpu.imm[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3167_));
 sky130_fd_sc_hd__nand2_1 _6792_ (.A(_3166_),
    .B(_3167_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3168_));
 sky130_fd_sc_hd__xnor2_1 _6793_ (.A(_3165_),
    .B(_3168_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3169_));
 sky130_fd_sc_hd__nand2_1 _6794_ (.A(_1390_),
    .B(_2536_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3170_));
 sky130_fd_sc_hd__o211a_1 _6795_ (.A1(_3040_),
    .A2(_3169_),
    .B1(_3170_),
    .C1(_3047_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3171_));
 sky130_fd_sc_hd__a221o_1 _6796_ (.A1(_3164_),
    .A2(_3039_),
    .B1(_2306_),
    .B2(_0915_),
    .C1(_3171_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3172_));
 sky130_fd_sc_hd__nand2_1 _6797_ (.A(_3037_),
    .B(_3172_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3173_));
 sky130_fd_sc_hd__o211a_1 _6798_ (.A1(\i_tinyqv.cpu.instr_data_start[16] ),
    .A2(_3123_),
    .B1(_3173_),
    .C1(_3093_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0457_));
 sky130_fd_sc_hd__inv_2 _6799_ (.A(net203),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3174_));
 sky130_fd_sc_hd__nand2_1 _6800_ (.A(\i_tinyqv.cpu.instr_data_start[17] ),
    .B(\i_tinyqv.cpu.imm[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3175_));
 sky130_fd_sc_hd__or2_1 _6801_ (.A(\i_tinyqv.cpu.instr_data_start[17] ),
    .B(\i_tinyqv.cpu.imm[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3176_));
 sky130_fd_sc_hd__nand2_1 _6802_ (.A(_3175_),
    .B(_3176_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3177_));
 sky130_fd_sc_hd__nand2_1 _6803_ (.A(_3167_),
    .B(_3165_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3178_));
 sky130_fd_sc_hd__nand2_1 _6804_ (.A(_3166_),
    .B(_3178_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3179_));
 sky130_fd_sc_hd__xnor2_1 _6805_ (.A(_3177_),
    .B(_3179_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3180_));
 sky130_fd_sc_hd__nand2_1 _6806_ (.A(_1390_),
    .B(_2538_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3181_));
 sky130_fd_sc_hd__o211a_1 _6807_ (.A1(_3040_),
    .A2(_3180_),
    .B1(_3181_),
    .C1(_3047_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3182_));
 sky130_fd_sc_hd__a221o_1 _6808_ (.A1(_3174_),
    .A2(_3039_),
    .B1(_2306_),
    .B2(_1213_),
    .C1(_3182_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3183_));
 sky130_fd_sc_hd__nand2_1 _6809_ (.A(_3037_),
    .B(_3183_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3184_));
 sky130_fd_sc_hd__o211a_1 _6810_ (.A1(\i_tinyqv.cpu.instr_data_start[17] ),
    .A2(_3123_),
    .B1(_3184_),
    .C1(_3093_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0458_));
 sky130_fd_sc_hd__inv_2 _6811_ (.A(\i_tinyqv.cpu.i_core.i_registers.registers[1][26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3185_));
 sky130_fd_sc_hd__o21a_1 _6812_ (.A1(_3177_),
    .A2(_3179_),
    .B1(_3175_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3186_));
 sky130_fd_sc_hd__nor2_1 _6813_ (.A(_0784_),
    .B(\i_tinyqv.cpu.imm[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3187_));
 sky130_fd_sc_hd__nand2_1 _6814_ (.A(_0784_),
    .B(\i_tinyqv.cpu.imm[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3188_));
 sky130_fd_sc_hd__or2b_1 _6815_ (.A(_3187_),
    .B_N(_3188_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3189_));
 sky130_fd_sc_hd__xnor2_1 _6816_ (.A(_3186_),
    .B(_3189_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3190_));
 sky130_fd_sc_hd__nand2_1 _6817_ (.A(_1390_),
    .B(_2540_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3191_));
 sky130_fd_sc_hd__o211a_1 _6818_ (.A1(_3040_),
    .A2(_3190_),
    .B1(_3191_),
    .C1(net40),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3192_));
 sky130_fd_sc_hd__a221o_1 _6819_ (.A1(_3185_),
    .A2(_3039_),
    .B1(_2306_),
    .B2(_1345_),
    .C1(_3192_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3193_));
 sky130_fd_sc_hd__nand2_1 _6820_ (.A(_3026_),
    .B(_3193_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3194_));
 sky130_fd_sc_hd__o211a_1 _6821_ (.A1(_0784_),
    .A2(_3123_),
    .B1(_3194_),
    .C1(_3093_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0459_));
 sky130_fd_sc_hd__nand2_1 _6822_ (.A(\i_tinyqv.cpu.instr_data_start[19] ),
    .B(\i_tinyqv.cpu.imm[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3195_));
 sky130_fd_sc_hd__or2_1 _6823_ (.A(\i_tinyqv.cpu.instr_data_start[19] ),
    .B(\i_tinyqv.cpu.imm[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3196_));
 sky130_fd_sc_hd__nand2_1 _6824_ (.A(_3195_),
    .B(_3196_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3197_));
 sky130_fd_sc_hd__o21ai_1 _6825_ (.A1(_3187_),
    .A2(_3186_),
    .B1(_3188_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3198_));
 sky130_fd_sc_hd__xor2_1 _6826_ (.A(_3197_),
    .B(_3198_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3199_));
 sky130_fd_sc_hd__nand2_1 _6827_ (.A(_3040_),
    .B(_2542_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3200_));
 sky130_fd_sc_hd__o211ai_1 _6828_ (.A1(_3040_),
    .A2(_3199_),
    .B1(_3200_),
    .C1(_3051_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3201_));
 sky130_fd_sc_hd__nor2_1 _6829_ (.A(_2987_),
    .B(_1601_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3202_));
 sky130_fd_sc_hd__a211o_1 _6830_ (.A1(\i_tinyqv.cpu.i_core.i_registers.registers[1][27] ),
    .A2(_2987_),
    .B1(_3202_),
    .C1(_2993_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3203_));
 sky130_fd_sc_hd__a21o_1 _6831_ (.A1(_3201_),
    .A2(_3203_),
    .B1(_3029_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3204_));
 sky130_fd_sc_hd__clkbuf_4 _6832_ (.A(_1752_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3205_));
 sky130_fd_sc_hd__o211a_1 _6833_ (.A1(\i_tinyqv.cpu.instr_data_start[19] ),
    .A2(_3123_),
    .B1(_3204_),
    .C1(_3205_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0460_));
 sky130_fd_sc_hd__mux2_1 _6834_ (.A0(_0902_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.registers[1][28] ),
    .S(net31),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3206_));
 sky130_fd_sc_hd__a21boi_1 _6835_ (.A1(_3196_),
    .A2(_3198_),
    .B1_N(_3195_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3207_));
 sky130_fd_sc_hd__nor2_1 _6836_ (.A(\i_tinyqv.cpu.instr_data_start[20] ),
    .B(\i_tinyqv.cpu.imm[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3208_));
 sky130_fd_sc_hd__nand2_1 _6837_ (.A(\i_tinyqv.cpu.instr_data_start[20] ),
    .B(\i_tinyqv.cpu.imm[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3209_));
 sky130_fd_sc_hd__or2b_1 _6838_ (.A(_3208_),
    .B_N(_3209_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3210_));
 sky130_fd_sc_hd__xor2_1 _6839_ (.A(_3207_),
    .B(_3210_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3211_));
 sky130_fd_sc_hd__mux2_1 _6840_ (.A0(_2544_),
    .A1(_3211_),
    .S(_2990_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3212_));
 sky130_fd_sc_hd__mux2_1 _6841_ (.A0(_3206_),
    .A1(_3212_),
    .S(_3047_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3213_));
 sky130_fd_sc_hd__or2_1 _6842_ (.A(_3029_),
    .B(_3213_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3214_));
 sky130_fd_sc_hd__o211a_1 _6843_ (.A1(\i_tinyqv.cpu.instr_data_start[20] ),
    .A2(_3123_),
    .B1(_3214_),
    .C1(_3205_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0461_));
 sky130_fd_sc_hd__nand2_1 _6844_ (.A(\i_tinyqv.cpu.instr_data_start[21] ),
    .B(\i_tinyqv.cpu.imm[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3215_));
 sky130_fd_sc_hd__or2_1 _6845_ (.A(\i_tinyqv.cpu.instr_data_start[21] ),
    .B(\i_tinyqv.cpu.imm[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3216_));
 sky130_fd_sc_hd__nand2_1 _6846_ (.A(_3215_),
    .B(_3216_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3217_));
 sky130_fd_sc_hd__o21ai_1 _6847_ (.A1(_3208_),
    .A2(_3207_),
    .B1(_3209_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3218_));
 sky130_fd_sc_hd__xnor2_1 _6848_ (.A(_3217_),
    .B(_3218_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3219_));
 sky130_fd_sc_hd__mux2_1 _6849_ (.A0(_2546_),
    .A1(_3219_),
    .S(_2991_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3220_));
 sky130_fd_sc_hd__a221o_1 _6850_ (.A1(\i_tinyqv.cpu.i_core.i_registers.registers[1][29] ),
    .A2(_2987_),
    .B1(_2306_),
    .B2(_1211_),
    .C1(_3028_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3221_));
 sky130_fd_sc_hd__a21o_1 _6851_ (.A1(_3051_),
    .A2(_3220_),
    .B1(_3221_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3222_));
 sky130_fd_sc_hd__o211a_1 _6852_ (.A1(\i_tinyqv.cpu.instr_data_start[21] ),
    .A2(_3123_),
    .B1(_3222_),
    .C1(_3205_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0462_));
 sky130_fd_sc_hd__mux2_1 _6853_ (.A0(_1335_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.registers[1][30] ),
    .S(net31),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3223_));
 sky130_fd_sc_hd__a21boi_1 _6854_ (.A1(_3216_),
    .A2(_3218_),
    .B1_N(_3215_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3224_));
 sky130_fd_sc_hd__nor2_1 _6855_ (.A(\i_tinyqv.cpu.instr_data_start[22] ),
    .B(\i_tinyqv.cpu.imm[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3225_));
 sky130_fd_sc_hd__nand2_1 _6856_ (.A(\i_tinyqv.cpu.instr_data_start[22] ),
    .B(\i_tinyqv.cpu.imm[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3226_));
 sky130_fd_sc_hd__or2b_1 _6857_ (.A(_3225_),
    .B_N(_3226_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3227_));
 sky130_fd_sc_hd__xor2_1 _6858_ (.A(_3224_),
    .B(_3227_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3228_));
 sky130_fd_sc_hd__mux2_1 _6859_ (.A0(_2548_),
    .A1(_3228_),
    .S(_2990_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3229_));
 sky130_fd_sc_hd__mux2_1 _6860_ (.A0(_3223_),
    .A1(_3229_),
    .S(_3047_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3230_));
 sky130_fd_sc_hd__or2_1 _6861_ (.A(_3028_),
    .B(_3230_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3231_));
 sky130_fd_sc_hd__o211a_1 _6862_ (.A1(\i_tinyqv.cpu.instr_data_start[22] ),
    .A2(_3123_),
    .B1(_3231_),
    .C1(_3205_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0463_));
 sky130_fd_sc_hd__o21ai_1 _6863_ (.A1(_3225_),
    .A2(_3224_),
    .B1(_3226_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3232_));
 sky130_fd_sc_hd__xnor2_1 _6864_ (.A(\i_tinyqv.cpu.instr_data_start[23] ),
    .B(\i_tinyqv.cpu.imm[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3233_));
 sky130_fd_sc_hd__xnor2_1 _6865_ (.A(_3232_),
    .B(_3233_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3234_));
 sky130_fd_sc_hd__or2_1 _6866_ (.A(_2991_),
    .B(_2550_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3235_));
 sky130_fd_sc_hd__o211a_1 _6867_ (.A1(_3040_),
    .A2(_3234_),
    .B1(_3235_),
    .C1(_2993_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3236_));
 sky130_fd_sc_hd__o21a_1 _6868_ (.A1(_1442_),
    .A2(_1599_),
    .B1(_2306_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3237_));
 sky130_fd_sc_hd__a211o_1 _6869_ (.A1(\i_tinyqv.cpu.i_core.i_registers.registers[1][31] ),
    .A2(_3039_),
    .B1(_3236_),
    .C1(_3237_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3238_));
 sky130_fd_sc_hd__o211a_1 _6870_ (.A1(\i_tinyqv.cpu.instr_data_start[23] ),
    .A2(_3037_),
    .B1(_3238_),
    .C1(_3205_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0464_));
 sky130_fd_sc_hd__clkbuf_4 _6871_ (.A(_1437_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3239_));
 sky130_fd_sc_hd__inv_2 _6872_ (.A(\i_tinyqv.cpu.instr_fetch_stopped ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3240_));
 sky130_fd_sc_hd__a21oi_1 _6873_ (.A1(\i_tinyqv.cpu.instr_fetch_running ),
    .A2(_3240_),
    .B1(net183),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3241_));
 sky130_fd_sc_hd__o21ba_1 _6874_ (.A1(_1550_),
    .A2(_3241_),
    .B1_N(_3051_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3242_));
 sky130_fd_sc_hd__a211oi_1 _6875_ (.A1(_3239_),
    .A2(_3051_),
    .B1(_3242_),
    .C1(_2066_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0465_));
 sky130_fd_sc_hd__a31o_1 _6876_ (.A1(_3017_),
    .A2(_2049_),
    .A3(_1604_),
    .B1(_1480_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0466_));
 sky130_fd_sc_hd__nand2_1 _6877_ (.A(\i_tinyqv.cpu.is_store ),
    .B(_1761_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3243_));
 sky130_fd_sc_hd__o21a_1 _6878_ (.A1(\i_tinyqv.cpu.data_write_n[0] ),
    .A2(_1556_),
    .B1(_3243_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3244_));
 sky130_fd_sc_hd__a211o_1 _6879_ (.A1(\i_tinyqv.cpu.i_core.mem_op[0] ),
    .A2(_1762_),
    .B1(_3244_),
    .C1(_2067_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0467_));
 sky130_fd_sc_hd__o21a_1 _6880_ (.A1(\i_tinyqv.cpu.data_write_n[1] ),
    .A2(_1556_),
    .B1(_3243_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3245_));
 sky130_fd_sc_hd__a211o_1 _6881_ (.A1(net258),
    .A2(_1762_),
    .B1(_3245_),
    .C1(_2067_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0468_));
 sky130_fd_sc_hd__a21o_1 _6882_ (.A1(\i_tinyqv.cpu.load_started ),
    .A2(_1556_),
    .B1(_1759_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3246_));
 sky130_fd_sc_hd__mux2_1 _6883_ (.A0(\i_tinyqv.cpu.data_read_n[0] ),
    .A1(\i_tinyqv.cpu.i_core.mem_op[0] ),
    .S(_1761_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3247_));
 sky130_fd_sc_hd__or2_1 _6884_ (.A(_3246_),
    .B(_3247_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3248_));
 sky130_fd_sc_hd__clkbuf_1 _6885_ (.A(_3248_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0469_));
 sky130_fd_sc_hd__mux2_1 _6886_ (.A0(\i_tinyqv.cpu.data_read_n[1] ),
    .A1(\i_tinyqv.cpu.i_core.mem_op[1] ),
    .S(_1761_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3249_));
 sky130_fd_sc_hd__or2_1 _6887_ (.A(_3246_),
    .B(_3249_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3250_));
 sky130_fd_sc_hd__clkbuf_1 _6888_ (.A(_3250_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0470_));
 sky130_fd_sc_hd__a211o_1 _6889_ (.A1(\i_tinyqv.cpu.data_write_n[1] ),
    .A2(net294),
    .B1(_0957_),
    .C1(_0979_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3251_));
 sky130_fd_sc_hd__a21o_1 _6890_ (.A1(\i_tinyqv.cpu.no_write_in_progress ),
    .A2(_1604_),
    .B1(_2066_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3252_));
 sky130_fd_sc_hd__a31o_1 _6891_ (.A1(_1387_),
    .A2(_3243_),
    .A3(_3251_),
    .B1(_3252_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0471_));
 sky130_fd_sc_hd__a31o_1 _6892_ (.A1(\i_tinyqv.cpu.is_load ),
    .A2(net144),
    .A3(_1442_),
    .B1(_1760_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0472_));
 sky130_fd_sc_hd__nor2_2 _6893_ (.A(_0612_),
    .B(_0854_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3253_));
 sky130_fd_sc_hd__and2_1 _6894_ (.A(_0752_),
    .B(_3253_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3254_));
 sky130_fd_sc_hd__mux2_1 _6895_ (.A0(\i_debug_uart_tx.uart_tx_data[0] ),
    .A1(_2641_),
    .S(_3254_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3255_));
 sky130_fd_sc_hd__clkbuf_1 _6896_ (.A(_3255_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0473_));
 sky130_fd_sc_hd__mux2_1 _6897_ (.A0(\i_debug_uart_tx.uart_tx_data[1] ),
    .A1(_2647_),
    .S(_3254_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3256_));
 sky130_fd_sc_hd__clkbuf_1 _6898_ (.A(_3256_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0474_));
 sky130_fd_sc_hd__inv_2 _6899_ (.A(net16),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3257_));
 sky130_fd_sc_hd__mux2_1 _6900_ (.A0(\i_debug_uart_tx.uart_tx_data[2] ),
    .A1(_3257_),
    .S(_3254_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3258_));
 sky130_fd_sc_hd__clkbuf_1 _6901_ (.A(_3258_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0475_));
 sky130_fd_sc_hd__mux2_1 _6902_ (.A0(\i_debug_uart_tx.uart_tx_data[3] ),
    .A1(_2631_),
    .S(_3254_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3259_));
 sky130_fd_sc_hd__clkbuf_1 _6903_ (.A(_3259_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0476_));
 sky130_fd_sc_hd__nand2_2 _6904_ (.A(_1026_),
    .B(_0955_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3260_));
 sky130_fd_sc_hd__nor2_2 _6905_ (.A(_2640_),
    .B(_3260_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3261_));
 sky130_fd_sc_hd__nand2_1 _6906_ (.A(_0956_),
    .B(_0612_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3262_));
 sky130_fd_sc_hd__and2_1 _6907_ (.A(_1026_),
    .B(_3262_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3263_));
 sky130_fd_sc_hd__and3_1 _6908_ (.A(\i_tinyqv.cpu.is_store ),
    .B(\i_tinyqv.cpu.no_write_in_progress ),
    .C(_3263_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3264_));
 sky130_fd_sc_hd__buf_2 _6909_ (.A(_3264_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3265_));
 sky130_fd_sc_hd__or2_1 _6910_ (.A(_0939_),
    .B(_0854_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3266_));
 sky130_fd_sc_hd__a32o_1 _6911_ (.A1(_1619_),
    .A2(_3261_),
    .A3(_3265_),
    .B1(_3266_),
    .B2(net309),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0477_));
 sky130_fd_sc_hd__nor2_2 _6912_ (.A(_0772_),
    .B(_3260_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3267_));
 sky130_fd_sc_hd__a32o_1 _6913_ (.A1(_1619_),
    .A2(_3265_),
    .A3(_3267_),
    .B1(_3266_),
    .B2(net313),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0478_));
 sky130_fd_sc_hd__nor2_2 _6914_ (.A(net16),
    .B(_3260_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3268_));
 sky130_fd_sc_hd__a32o_1 _6915_ (.A1(_1619_),
    .A2(_3265_),
    .A3(_3268_),
    .B1(_3266_),
    .B2(net234),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0479_));
 sky130_fd_sc_hd__nor2_2 _6916_ (.A(net50),
    .B(_3260_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3269_));
 sky130_fd_sc_hd__a32o_1 _6917_ (.A1(_1619_),
    .A2(_3265_),
    .A3(_3269_),
    .B1(_3266_),
    .B2(net273),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0480_));
 sky130_fd_sc_hd__or3_2 _6918_ (.A(_0956_),
    .B(_0909_),
    .C(_0854_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3270_));
 sky130_fd_sc_hd__a32o_1 _6919_ (.A1(_0691_),
    .A2(_3261_),
    .A3(_3265_),
    .B1(_3270_),
    .B2(net186),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0481_));
 sky130_fd_sc_hd__a32o_1 _6920_ (.A1(_0691_),
    .A2(_3265_),
    .A3(_3267_),
    .B1(_3270_),
    .B2(net169),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0482_));
 sky130_fd_sc_hd__a32o_1 _6921_ (.A1(_0691_),
    .A2(_3265_),
    .A3(_3268_),
    .B1(_3270_),
    .B2(net132),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0483_));
 sky130_fd_sc_hd__a32o_1 _6922_ (.A1(_0691_),
    .A2(_3265_),
    .A3(_3269_),
    .B1(_3270_),
    .B2(net131),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0484_));
 sky130_fd_sc_hd__or3_2 _6923_ (.A(_0956_),
    .B(_0724_),
    .C(_0854_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3271_));
 sky130_fd_sc_hd__a32o_1 _6924_ (.A1(_1589_),
    .A2(_3261_),
    .A3(_3265_),
    .B1(_3271_),
    .B2(net149),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0485_));
 sky130_fd_sc_hd__a32o_1 _6925_ (.A1(_1589_),
    .A2(_3265_),
    .A3(_3267_),
    .B1(_3271_),
    .B2(net136),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0486_));
 sky130_fd_sc_hd__a32o_1 _6926_ (.A1(_1589_),
    .A2(_3264_),
    .A3(_3268_),
    .B1(_3271_),
    .B2(net130),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0487_));
 sky130_fd_sc_hd__a32o_1 _6927_ (.A1(_1589_),
    .A2(_3264_),
    .A3(_3269_),
    .B1(_3271_),
    .B2(net125),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0488_));
 sky130_fd_sc_hd__or2_1 _6928_ (.A(_0916_),
    .B(_0854_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3272_));
 sky130_fd_sc_hd__a22o_1 _6929_ (.A1(_3253_),
    .A2(_3261_),
    .B1(_3272_),
    .B2(net156),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0489_));
 sky130_fd_sc_hd__a22o_1 _6930_ (.A1(_3253_),
    .A2(_3267_),
    .B1(_3272_),
    .B2(net140),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0490_));
 sky130_fd_sc_hd__a22o_1 _6931_ (.A1(_3253_),
    .A2(_3268_),
    .B1(_3272_),
    .B2(net175),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0491_));
 sky130_fd_sc_hd__a22o_1 _6932_ (.A1(_3253_),
    .A2(_3269_),
    .B1(_3272_),
    .B2(net143),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0492_));
 sky130_fd_sc_hd__nor2_1 _6933_ (.A(_0854_),
    .B(_3263_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3273_));
 sky130_fd_sc_hd__buf_2 _6934_ (.A(_3273_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3274_));
 sky130_fd_sc_hd__or2_1 _6935_ (.A(_2081_),
    .B(_0854_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3275_));
 sky130_fd_sc_hd__a32o_1 _6936_ (.A1(_1619_),
    .A2(_3261_),
    .A3(_3274_),
    .B1(_3275_),
    .B2(net129),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0493_));
 sky130_fd_sc_hd__a32o_1 _6937_ (.A1(_1619_),
    .A2(_3267_),
    .A3(_3274_),
    .B1(_3275_),
    .B2(net112),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0494_));
 sky130_fd_sc_hd__a32o_1 _6938_ (.A1(_1619_),
    .A2(_3268_),
    .A3(_3274_),
    .B1(_3275_),
    .B2(net115),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0495_));
 sky130_fd_sc_hd__a32o_1 _6939_ (.A1(_1619_),
    .A2(_3269_),
    .A3(_3274_),
    .B1(_3275_),
    .B2(net113),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0496_));
 sky130_fd_sc_hd__or2_1 _6940_ (.A(_0630_),
    .B(_0854_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3276_));
 sky130_fd_sc_hd__a32o_1 _6941_ (.A1(_0691_),
    .A2(_3261_),
    .A3(_3274_),
    .B1(_3276_),
    .B2(net107),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0497_));
 sky130_fd_sc_hd__a32o_1 _6942_ (.A1(_0691_),
    .A2(_3267_),
    .A3(_3274_),
    .B1(_3276_),
    .B2(net118),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0498_));
 sky130_fd_sc_hd__a32o_1 _6943_ (.A1(_0691_),
    .A2(_3268_),
    .A3(_3274_),
    .B1(_3276_),
    .B2(net119),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0499_));
 sky130_fd_sc_hd__a32o_1 _6944_ (.A1(_0691_),
    .A2(_3269_),
    .A3(_3274_),
    .B1(_3276_),
    .B2(net124),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0500_));
 sky130_fd_sc_hd__or2_1 _6945_ (.A(_1604_),
    .B(_0854_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3277_));
 sky130_fd_sc_hd__a32o_1 _6946_ (.A1(_1589_),
    .A2(_3261_),
    .A3(_3274_),
    .B1(_3277_),
    .B2(net114),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0501_));
 sky130_fd_sc_hd__a32o_1 _6947_ (.A1(_1589_),
    .A2(_3267_),
    .A3(_3274_),
    .B1(_3277_),
    .B2(net109),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0502_));
 sky130_fd_sc_hd__a32o_1 _6948_ (.A1(_1589_),
    .A2(_3268_),
    .A3(_3273_),
    .B1(_3277_),
    .B2(net120),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0503_));
 sky130_fd_sc_hd__a32o_1 _6949_ (.A1(_1589_),
    .A2(_3269_),
    .A3(_3273_),
    .B1(_3277_),
    .B2(net110),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0504_));
 sky130_fd_sc_hd__nor2_1 _6950_ (.A(_2066_),
    .B(_0974_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0505_));
 sky130_fd_sc_hd__and3_1 _6951_ (.A(_2079_),
    .B(_0612_),
    .C(_0724_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3278_));
 sky130_fd_sc_hd__clkbuf_1 _6952_ (.A(_3278_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0506_));
 sky130_fd_sc_hd__o22a_1 _6953_ (.A1(_0956_),
    .A2(_1589_),
    .B1(_2087_),
    .B2(_0505_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0507_));
 sky130_fd_sc_hd__or3_1 _6954_ (.A(\i_tinyqv.cpu.data_ready_latch ),
    .B(_1604_),
    .C(_1556_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3279_));
 sky130_fd_sc_hd__o211a_1 _6955_ (.A1(net236),
    .A2(_1387_),
    .B1(_3279_),
    .C1(_3205_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0508_));
 sky130_fd_sc_hd__o211a_1 _6956_ (.A1(net180),
    .A2(_1556_),
    .B1(_1604_),
    .C1(_3205_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0509_));
 sky130_fd_sc_hd__and2_1 _6957_ (.A(_2146_),
    .B(_2151_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3280_));
 sky130_fd_sc_hd__buf_2 _6958_ (.A(_3280_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3281_));
 sky130_fd_sc_hd__clkbuf_4 _6959_ (.A(_3281_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3282_));
 sky130_fd_sc_hd__or3_1 _6960_ (.A(_1468_),
    .B(_1483_),
    .C(_1487_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3283_));
 sky130_fd_sc_hd__inv_2 _6961_ (.A(_3283_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3284_));
 sky130_fd_sc_hd__mux2_1 _6962_ (.A0(\i_tinyqv.cpu.instr_data[1][11] ),
    .A1(\i_tinyqv.cpu.instr_data[3][11] ),
    .S(_1504_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3285_));
 sky130_fd_sc_hd__mux2_1 _6963_ (.A0(\i_tinyqv.cpu.instr_data[0][11] ),
    .A1(\i_tinyqv.cpu.instr_data[2][11] ),
    .S(_1504_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3286_));
 sky130_fd_sc_hd__mux2_4 _6964_ (.A0(_3285_),
    .A1(_3286_),
    .S(_1432_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3287_));
 sky130_fd_sc_hd__inv_2 _6965_ (.A(_3287_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3288_));
 sky130_fd_sc_hd__nor2_2 _6966_ (.A(_1420_),
    .B(_1426_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3289_));
 sky130_fd_sc_hd__buf_2 _6967_ (.A(_3289_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3290_));
 sky130_fd_sc_hd__clkbuf_4 _6968_ (.A(_3290_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3291_));
 sky130_fd_sc_hd__and4_2 _6969_ (.A(_1420_),
    .B(_1426_),
    .C(_1473_),
    .D(_2124_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3292_));
 sky130_fd_sc_hd__a22o_1 _6970_ (.A1(_1483_),
    .A2(_2132_),
    .B1(_3292_),
    .B2(_2118_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3293_));
 sky130_fd_sc_hd__a21o_1 _6971_ (.A1(_3291_),
    .A2(_2135_),
    .B1(_3293_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3294_));
 sky130_fd_sc_hd__nand2_2 _6972_ (.A(_2147_),
    .B(_2151_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3295_));
 sky130_fd_sc_hd__a211o_1 _6973_ (.A1(_3284_),
    .A2(_3288_),
    .B1(_3294_),
    .C1(_3295_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3296_));
 sky130_fd_sc_hd__o211a_1 _6974_ (.A1(\i_tinyqv.cpu.is_load ),
    .A2(_3282_),
    .B1(_3296_),
    .C1(_3205_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0510_));
 sky130_fd_sc_hd__or2_1 _6975_ (.A(_1483_),
    .B(_2127_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3297_));
 sky130_fd_sc_hd__a21o_1 _6976_ (.A1(_1461_),
    .A2(_1503_),
    .B1(_1506_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3298_));
 sky130_fd_sc_hd__buf_2 _6977_ (.A(_3298_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3299_));
 sky130_fd_sc_hd__nand2_1 _6978_ (.A(_1498_),
    .B(_3287_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3300_));
 sky130_fd_sc_hd__nor2_1 _6979_ (.A(_3299_),
    .B(_3300_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3301_));
 sky130_fd_sc_hd__or3_1 _6980_ (.A(_1483_),
    .B(_2119_),
    .C(_3301_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3302_));
 sky130_fd_sc_hd__o211a_1 _6981_ (.A1(_2123_),
    .A2(_2122_),
    .B1(_3297_),
    .C1(_3302_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3303_));
 sky130_fd_sc_hd__clkbuf_4 _6982_ (.A(_1452_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3304_));
 sky130_fd_sc_hd__clkbuf_4 _6983_ (.A(_1455_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3305_));
 sky130_fd_sc_hd__or3_1 _6984_ (.A(_2140_),
    .B(_1465_),
    .C(_1492_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3306_));
 sky130_fd_sc_hd__or2_1 _6985_ (.A(_1502_),
    .B(_1510_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3307_));
 sky130_fd_sc_hd__nor2b_2 _6986_ (.A(_3307_),
    .B_N(_1514_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3308_));
 sky130_fd_sc_hd__nand2_1 _6987_ (.A(_2126_),
    .B(_3308_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3309_));
 sky130_fd_sc_hd__o31a_1 _6988_ (.A1(_3304_),
    .A2(_3305_),
    .A3(_3306_),
    .B1(_3309_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3310_));
 sky130_fd_sc_hd__a31o_1 _6989_ (.A1(_3281_),
    .A2(_3303_),
    .A3(_3310_),
    .B1(_2066_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3311_));
 sky130_fd_sc_hd__o21ba_1 _6990_ (.A1(net249),
    .A2(_3282_),
    .B1_N(_3311_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0511_));
 sky130_fd_sc_hd__nand2_2 _6991_ (.A(_3291_),
    .B(_3281_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3312_));
 sky130_fd_sc_hd__inv_2 _6992_ (.A(_1460_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3313_));
 sky130_fd_sc_hd__or3_2 _6993_ (.A(_2155_),
    .B(_3313_),
    .C(_1465_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3314_));
 sky130_fd_sc_hd__or2_4 _6994_ (.A(_3305_),
    .B(_3314_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3315_));
 sky130_fd_sc_hd__inv_2 _6995_ (.A(\i_tinyqv.cpu.is_auipc ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3316_));
 sky130_fd_sc_hd__o32a_1 _6996_ (.A1(_3304_),
    .A2(_3312_),
    .A3(_3315_),
    .B1(_3282_),
    .B2(_3316_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3317_));
 sky130_fd_sc_hd__nor2_1 _6997_ (.A(_2067_),
    .B(_3317_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0512_));
 sky130_fd_sc_hd__or3b_1 _6998_ (.A(_1491_),
    .B(_1492_),
    .C_N(_1452_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3318_));
 sky130_fd_sc_hd__buf_2 _6999_ (.A(_3318_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3319_));
 sky130_fd_sc_hd__nor2_1 _7000_ (.A(_3305_),
    .B(_3319_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3320_));
 sky130_fd_sc_hd__nand2_1 _7001_ (.A(_1420_),
    .B(_1476_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3321_));
 sky130_fd_sc_hd__nor2_2 _7002_ (.A(_2118_),
    .B(_3321_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3322_));
 sky130_fd_sc_hd__a211o_1 _7003_ (.A1(_3284_),
    .A2(_3287_),
    .B1(_3322_),
    .C1(_3290_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3323_));
 sky130_fd_sc_hd__mux2_1 _7004_ (.A0(\i_tinyqv.cpu.is_store ),
    .A1(_3323_),
    .S(_3281_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3324_));
 sky130_fd_sc_hd__o211a_1 _7005_ (.A1(_3312_),
    .A2(_3320_),
    .B1(_3324_),
    .C1(_3205_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0513_));
 sky130_fd_sc_hd__and4bb_1 _7006_ (.A_N(_3305_),
    .B_N(_1492_),
    .C(_1491_),
    .D(_1452_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3325_));
 sky130_fd_sc_hd__a211o_1 _7007_ (.A1(_2121_),
    .A2(_3301_),
    .B1(_2136_),
    .C1(_2131_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3326_));
 sky130_fd_sc_hd__mux2_1 _7008_ (.A0(\i_tinyqv.cpu.is_alu_reg ),
    .A1(_3326_),
    .S(_3281_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3327_));
 sky130_fd_sc_hd__o211a_1 _7009_ (.A1(_3312_),
    .A2(_3325_),
    .B1(_3327_),
    .C1(_3205_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0514_));
 sky130_fd_sc_hd__buf_2 _7010_ (.A(_3290_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3328_));
 sky130_fd_sc_hd__nor2_1 _7011_ (.A(_3305_),
    .B(_3314_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3329_));
 sky130_fd_sc_hd__buf_2 _7012_ (.A(_3329_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3330_));
 sky130_fd_sc_hd__and2b_2 _7013_ (.A_N(_3308_),
    .B(_2126_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3331_));
 sky130_fd_sc_hd__a311o_1 _7014_ (.A1(_3328_),
    .A2(_3304_),
    .A3(_3330_),
    .B1(_3331_),
    .C1(_3295_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3332_));
 sky130_fd_sc_hd__o211a_1 _7015_ (.A1(net212),
    .A2(_3282_),
    .B1(_3332_),
    .C1(_1753_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0515_));
 sky130_fd_sc_hd__nor2_1 _7016_ (.A(_2140_),
    .B(_3295_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3333_));
 sky130_fd_sc_hd__inv_2 _7017_ (.A(_1455_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3334_));
 sky130_fd_sc_hd__nor2_1 _7018_ (.A(_3334_),
    .B(_3319_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3335_));
 sky130_fd_sc_hd__and2b_1 _7019_ (.A_N(_2119_),
    .B(_1476_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3336_));
 sky130_fd_sc_hd__clkbuf_4 _7020_ (.A(_3336_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3337_));
 sky130_fd_sc_hd__mux2_1 _7021_ (.A0(\i_tinyqv.cpu.is_branch ),
    .A1(_3337_),
    .S(_3281_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3338_));
 sky130_fd_sc_hd__a21oi_1 _7022_ (.A1(_3333_),
    .A2(_3335_),
    .B1(_3338_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3339_));
 sky130_fd_sc_hd__nor2_1 _7023_ (.A(_2067_),
    .B(_3339_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0516_));
 sky130_fd_sc_hd__and2_1 _7024_ (.A(\i_tinyqv.cpu.is_jalr ),
    .B(_3295_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3340_));
 sky130_fd_sc_hd__nor2_1 _7025_ (.A(_1490_),
    .B(_1494_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3341_));
 sky130_fd_sc_hd__or3_1 _7026_ (.A(_1514_),
    .B(_3287_),
    .C(_3307_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3342_));
 sky130_fd_sc_hd__and3_1 _7027_ (.A(_3341_),
    .B(_3281_),
    .C(_3342_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3343_));
 sky130_fd_sc_hd__and3b_1 _7028_ (.A_N(_2155_),
    .B(_1466_),
    .C(_3333_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3344_));
 sky130_fd_sc_hd__o31a_1 _7029_ (.A1(_3340_),
    .A2(_3343_),
    .A3(_3344_),
    .B1(_2061_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0517_));
 sky130_fd_sc_hd__nand2_1 _7030_ (.A(_1479_),
    .B(_3282_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3345_));
 sky130_fd_sc_hd__o211a_1 _7031_ (.A1(\i_tinyqv.cpu.is_jal ),
    .A2(_3282_),
    .B1(_3345_),
    .C1(_1753_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0518_));
 sky130_fd_sc_hd__nor2_1 _7032_ (.A(_2120_),
    .B(_2130_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3346_));
 sky130_fd_sc_hd__nor2_1 _7033_ (.A(_1478_),
    .B(_3337_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3347_));
 sky130_fd_sc_hd__nand2_1 _7034_ (.A(_3346_),
    .B(_3347_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3348_));
 sky130_fd_sc_hd__nor2_1 _7035_ (.A(_1468_),
    .B(_3297_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3349_));
 sky130_fd_sc_hd__and2_1 _7036_ (.A(_1468_),
    .B(_3322_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3350_));
 sky130_fd_sc_hd__and3_2 _7037_ (.A(_1426_),
    .B(_2123_),
    .C(_3322_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3351_));
 sky130_fd_sc_hd__or3_2 _7038_ (.A(_3349_),
    .B(_3350_),
    .C(_3351_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3352_));
 sky130_fd_sc_hd__or2_1 _7039_ (.A(_3292_),
    .B(_3284_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3353_));
 sky130_fd_sc_hd__or4_1 _7040_ (.A(_2126_),
    .B(_2138_),
    .C(_3352_),
    .D(_3353_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3354_));
 sky130_fd_sc_hd__or2_1 _7041_ (.A(_3348_),
    .B(_3354_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3355_));
 sky130_fd_sc_hd__o22a_1 _7042_ (.A1(_1456_),
    .A2(_3306_),
    .B1(_3355_),
    .B2(_1468_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3356_));
 sky130_fd_sc_hd__o211ai_1 _7043_ (.A1(_1495_),
    .A2(_3342_),
    .B1(_3356_),
    .C1(_3282_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3357_));
 sky130_fd_sc_hd__o211a_1 _7044_ (.A1(net209),
    .A2(_3282_),
    .B1(_3357_),
    .C1(_1753_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0519_));
 sky130_fd_sc_hd__nor2_1 _7045_ (.A(_1400_),
    .B(_3295_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3358_));
 sky130_fd_sc_hd__buf_2 _7046_ (.A(_3358_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3359_));
 sky130_fd_sc_hd__clkbuf_4 _7047_ (.A(_3359_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3360_));
 sky130_fd_sc_hd__nand2_1 _7048_ (.A(\i_tinyqv.cpu.i_core.i_cycles.rstn ),
    .B(_3281_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3361_));
 sky130_fd_sc_hd__buf_2 _7049_ (.A(_3361_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3362_));
 sky130_fd_sc_hd__nor2_1 _7050_ (.A(_2140_),
    .B(_3329_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3363_));
 sky130_fd_sc_hd__buf_2 _7051_ (.A(_3363_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3364_));
 sky130_fd_sc_hd__nand2_1 _7052_ (.A(_1504_),
    .B(_1461_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3365_));
 sky130_fd_sc_hd__clkbuf_4 _7053_ (.A(_3365_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3366_));
 sky130_fd_sc_hd__nand2_1 _7054_ (.A(_1422_),
    .B(_1432_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3367_));
 sky130_fd_sc_hd__clkbuf_4 _7055_ (.A(_3367_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3368_));
 sky130_fd_sc_hd__clkbuf_4 _7056_ (.A(_1504_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3369_));
 sky130_fd_sc_hd__clkbuf_4 _7057_ (.A(_1461_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3370_));
 sky130_fd_sc_hd__nand2_1 _7058_ (.A(_3365_),
    .B(_3367_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3371_));
 sky130_fd_sc_hd__clkbuf_4 _7059_ (.A(_3371_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3372_));
 sky130_fd_sc_hd__a221o_1 _7060_ (.A1(\i_tinyqv.cpu.instr_data[3][4] ),
    .A2(_3369_),
    .B1(_3370_),
    .B2(\i_tinyqv.cpu.instr_data[2][4] ),
    .C1(_3372_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3373_));
 sky130_fd_sc_hd__o221a_2 _7061_ (.A1(\i_tinyqv.cpu.instr_data[0][4] ),
    .A2(_3366_),
    .B1(_3368_),
    .B2(\i_tinyqv.cpu.instr_data[1][4] ),
    .C1(_3373_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3374_));
 sky130_fd_sc_hd__a32o_1 _7062_ (.A1(_1467_),
    .A2(_3319_),
    .A3(_3374_),
    .B1(_3320_),
    .B2(_1510_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3375_));
 sky130_fd_sc_hd__and2_1 _7063_ (.A(_3364_),
    .B(_3375_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3376_));
 sky130_fd_sc_hd__and3b_1 _7064_ (.A_N(_3300_),
    .B(_3299_),
    .C(_2121_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3377_));
 sky130_fd_sc_hd__or3_1 _7065_ (.A(_3334_),
    .B(_2165_),
    .C(_3283_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3378_));
 sky130_fd_sc_hd__o221a_1 _7066_ (.A1(_1490_),
    .A2(_3342_),
    .B1(_3346_),
    .B2(_3313_),
    .C1(_3378_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3379_));
 sky130_fd_sc_hd__or4b_2 _7067_ (.A(_3362_),
    .B(_3376_),
    .C(_3377_),
    .D_N(_3379_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3380_));
 sky130_fd_sc_hd__o21a_1 _7068_ (.A1(net221),
    .A2(_3360_),
    .B1(_3380_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0520_));
 sky130_fd_sc_hd__a22o_1 _7069_ (.A1(_1452_),
    .A2(_3284_),
    .B1(_3348_),
    .B2(_2155_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3381_));
 sky130_fd_sc_hd__or3b_1 _7070_ (.A(_3381_),
    .B(_3377_),
    .C_N(_3355_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3382_));
 sky130_fd_sc_hd__a221o_1 _7071_ (.A1(\i_tinyqv.cpu.instr_data[3][5] ),
    .A2(_3369_),
    .B1(_3370_),
    .B2(\i_tinyqv.cpu.instr_data[2][5] ),
    .C1(_3372_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3383_));
 sky130_fd_sc_hd__o221a_2 _7072_ (.A1(\i_tinyqv.cpu.instr_data[0][5] ),
    .A2(_3366_),
    .B1(_3368_),
    .B2(\i_tinyqv.cpu.instr_data[1][5] ),
    .C1(_3383_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3384_));
 sky130_fd_sc_hd__mux2_1 _7073_ (.A0(_1514_),
    .A1(_3384_),
    .S(_3319_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3385_));
 sky130_fd_sc_hd__a22o_1 _7074_ (.A1(_2140_),
    .A2(_3382_),
    .B1(_3385_),
    .B2(_3364_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3386_));
 sky130_fd_sc_hd__mux2_1 _7075_ (.A0(\i_tinyqv.cpu.i_core.imm_lo[1] ),
    .A1(_3386_),
    .S(_3359_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3387_));
 sky130_fd_sc_hd__clkbuf_1 _7076_ (.A(_3387_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0521_));
 sky130_fd_sc_hd__o21a_1 _7077_ (.A1(_1491_),
    .A2(_3377_),
    .B1(_3348_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3388_));
 sky130_fd_sc_hd__a221o_1 _7078_ (.A1(\i_tinyqv.cpu.instr_data[3][6] ),
    .A2(_1504_),
    .B1(_1461_),
    .B2(\i_tinyqv.cpu.instr_data[2][6] ),
    .C1(_3371_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3389_));
 sky130_fd_sc_hd__o221a_2 _7079_ (.A1(\i_tinyqv.cpu.instr_data[0][6] ),
    .A2(_3365_),
    .B1(_3367_),
    .B2(\i_tinyqv.cpu.instr_data[1][6] ),
    .C1(_3389_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3390_));
 sky130_fd_sc_hd__mux2_1 _7080_ (.A0(_1501_),
    .A1(_3390_),
    .S(_3319_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3391_));
 sky130_fd_sc_hd__o21a_1 _7081_ (.A1(_3292_),
    .A2(_3349_),
    .B1(_3305_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3392_));
 sky130_fd_sc_hd__a221o_1 _7082_ (.A1(_1501_),
    .A2(_3350_),
    .B1(_3363_),
    .B2(_3391_),
    .C1(_3392_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3393_));
 sky130_fd_sc_hd__a211o_1 _7083_ (.A1(_1491_),
    .A2(_2133_),
    .B1(_3388_),
    .C1(_3393_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3394_));
 sky130_fd_sc_hd__buf_4 _7084_ (.A(_3358_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3395_));
 sky130_fd_sc_hd__clkbuf_4 _7085_ (.A(_3395_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3396_));
 sky130_fd_sc_hd__mux2_1 _7086_ (.A0(\i_tinyqv.cpu.i_core.imm_lo[2] ),
    .A1(_3394_),
    .S(_3396_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3397_));
 sky130_fd_sc_hd__clkbuf_1 _7087_ (.A(_3397_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0522_));
 sky130_fd_sc_hd__or2_1 _7088_ (.A(_1478_),
    .B(_3349_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3398_));
 sky130_fd_sc_hd__or3_1 _7089_ (.A(_2121_),
    .B(_2130_),
    .C(_2133_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3399_));
 sky130_fd_sc_hd__o21a_1 _7090_ (.A1(_3398_),
    .A2(_3399_),
    .B1(_3304_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3400_));
 sky130_fd_sc_hd__a221o_1 _7091_ (.A1(\i_tinyqv.cpu.instr_data[3][7] ),
    .A2(_3369_),
    .B1(_3370_),
    .B2(\i_tinyqv.cpu.instr_data[2][7] ),
    .C1(_3372_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3401_));
 sky130_fd_sc_hd__o221a_1 _7092_ (.A1(\i_tinyqv.cpu.instr_data[0][7] ),
    .A2(_3366_),
    .B1(_3368_),
    .B2(\i_tinyqv.cpu.instr_data[1][7] ),
    .C1(_3401_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3402_));
 sky130_fd_sc_hd__mux2_1 _7093_ (.A0(_2165_),
    .A1(_3402_),
    .S(_3319_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3403_));
 sky130_fd_sc_hd__or3_1 _7094_ (.A(_3292_),
    .B(_3337_),
    .C(_3350_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3404_));
 sky130_fd_sc_hd__a22o_1 _7095_ (.A1(_3364_),
    .A2(_3403_),
    .B1(_3404_),
    .B2(_2165_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3405_));
 sky130_fd_sc_hd__or4_1 _7096_ (.A(_3362_),
    .B(_3377_),
    .C(_3400_),
    .D(_3405_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3406_));
 sky130_fd_sc_hd__o21a_1 _7097_ (.A1(\i_tinyqv.cpu.i_core.imm_lo[3] ),
    .A2(_3360_),
    .B1(_3406_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0523_));
 sky130_fd_sc_hd__a221o_1 _7098_ (.A1(\i_tinyqv.cpu.instr_data[3][8] ),
    .A2(_3369_),
    .B1(_3370_),
    .B2(\i_tinyqv.cpu.instr_data[2][8] ),
    .C1(_3372_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3407_));
 sky130_fd_sc_hd__o221a_1 _7099_ (.A1(\i_tinyqv.cpu.instr_data[0][8] ),
    .A2(_3366_),
    .B1(_3368_),
    .B2(\i_tinyqv.cpu.instr_data[1][8] ),
    .C1(_3407_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3408_));
 sky130_fd_sc_hd__mux2_1 _7100_ (.A0(_3287_),
    .A1(_3408_),
    .S(_3319_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3409_));
 sky130_fd_sc_hd__o41a_1 _7101_ (.A1(_1478_),
    .A2(_3292_),
    .A3(_3337_),
    .A4(_3352_),
    .B1(_3287_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3410_));
 sky130_fd_sc_hd__a32o_1 _7102_ (.A1(_3305_),
    .A2(_2126_),
    .A3(_3308_),
    .B1(_2132_),
    .B2(_1483_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3411_));
 sky130_fd_sc_hd__o32a_1 _7103_ (.A1(_2121_),
    .A2(_2130_),
    .A3(_3411_),
    .B1(_3377_),
    .B2(_3305_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3412_));
 sky130_fd_sc_hd__a211o_1 _7104_ (.A1(_3364_),
    .A2(_3409_),
    .B1(_3410_),
    .C1(_3412_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3413_));
 sky130_fd_sc_hd__mux2_1 _7105_ (.A0(\i_tinyqv.cpu.i_core.imm_lo[4] ),
    .A1(_3413_),
    .S(_3396_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3414_));
 sky130_fd_sc_hd__clkbuf_1 _7106_ (.A(_3414_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0524_));
 sky130_fd_sc_hd__a21oi_1 _7107_ (.A1(_2126_),
    .A2(_3308_),
    .B1(_2143_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3415_));
 sky130_fd_sc_hd__nand2_1 _7108_ (.A(_3347_),
    .B(_3415_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3416_));
 sky130_fd_sc_hd__a221o_1 _7109_ (.A1(\i_tinyqv.cpu.instr_data[3][9] ),
    .A2(_3369_),
    .B1(_3370_),
    .B2(\i_tinyqv.cpu.instr_data[2][9] ),
    .C1(_3372_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3417_));
 sky130_fd_sc_hd__o221a_1 _7110_ (.A1(\i_tinyqv.cpu.instr_data[0][9] ),
    .A2(_3366_),
    .B1(_3368_),
    .B2(\i_tinyqv.cpu.instr_data[1][9] ),
    .C1(_3417_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3418_));
 sky130_fd_sc_hd__a22o_1 _7111_ (.A1(_2165_),
    .A2(_3351_),
    .B1(_3363_),
    .B2(_3418_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3419_));
 sky130_fd_sc_hd__o41a_1 _7112_ (.A1(_3292_),
    .A2(_3349_),
    .A3(_3350_),
    .A4(_3399_),
    .B1(_3299_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3420_));
 sky130_fd_sc_hd__a211o_1 _7113_ (.A1(_1460_),
    .A2(_3416_),
    .B1(_3419_),
    .C1(_3420_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3421_));
 sky130_fd_sc_hd__mux2_1 _7114_ (.A0(\i_tinyqv.cpu.i_core.imm_lo[5] ),
    .A1(_3421_),
    .S(_3396_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3422_));
 sky130_fd_sc_hd__clkbuf_1 _7115_ (.A(_3422_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0525_));
 sky130_fd_sc_hd__inv_2 _7116_ (.A(_3415_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3423_));
 sky130_fd_sc_hd__o31a_1 _7117_ (.A1(_3292_),
    .A2(_3337_),
    .A3(_3423_),
    .B1(_3304_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3424_));
 sky130_fd_sc_hd__nor2_1 _7118_ (.A(_1507_),
    .B(_3346_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3425_));
 sky130_fd_sc_hd__a221o_1 _7119_ (.A1(\i_tinyqv.cpu.instr_data[3][10] ),
    .A2(_1504_),
    .B1(_1461_),
    .B2(\i_tinyqv.cpu.instr_data[2][10] ),
    .C1(_3371_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3426_));
 sky130_fd_sc_hd__o221a_1 _7120_ (.A1(\i_tinyqv.cpu.instr_data[0][10] ),
    .A2(_3365_),
    .B1(_3367_),
    .B2(\i_tinyqv.cpu.instr_data[1][10] ),
    .C1(_3426_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3427_));
 sky130_fd_sc_hd__nand2_1 _7121_ (.A(_3289_),
    .B(_3427_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3428_));
 sky130_fd_sc_hd__a2bb2o_1 _7122_ (.A1_N(_3428_),
    .A2_N(_3329_),
    .B1(_2133_),
    .B2(_1460_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3429_));
 sky130_fd_sc_hd__o21a_1 _7123_ (.A1(_1478_),
    .A2(_3352_),
    .B1(_1510_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3430_));
 sky130_fd_sc_hd__or4_1 _7124_ (.A(_3424_),
    .B(_3425_),
    .C(_3429_),
    .D(_3430_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3431_));
 sky130_fd_sc_hd__mux2_1 _7125_ (.A0(\i_tinyqv.cpu.i_core.imm_lo[6] ),
    .A1(_3431_),
    .S(_3396_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3432_));
 sky130_fd_sc_hd__clkbuf_1 _7126_ (.A(_3432_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0526_));
 sky130_fd_sc_hd__a221o_1 _7127_ (.A1(\i_tinyqv.cpu.instr_data[3][11] ),
    .A2(_3369_),
    .B1(_3370_),
    .B2(\i_tinyqv.cpu.instr_data[2][11] ),
    .C1(_3372_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3433_));
 sky130_fd_sc_hd__o221a_1 _7128_ (.A1(\i_tinyqv.cpu.instr_data[0][11] ),
    .A2(_3366_),
    .B1(_3368_),
    .B2(\i_tinyqv.cpu.instr_data[1][11] ),
    .C1(_3433_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3434_));
 sky130_fd_sc_hd__a22o_1 _7129_ (.A1(_1483_),
    .A2(_2132_),
    .B1(_3308_),
    .B2(_2126_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3435_));
 sky130_fd_sc_hd__o22ai_1 _7130_ (.A1(_1507_),
    .A2(_3346_),
    .B1(_3347_),
    .B2(_3334_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3436_));
 sky130_fd_sc_hd__a221o_1 _7131_ (.A1(_1514_),
    .A2(_3352_),
    .B1(_3435_),
    .B2(_2155_),
    .C1(_3436_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3437_));
 sky130_fd_sc_hd__clkbuf_4 _7132_ (.A(_3361_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3438_));
 sky130_fd_sc_hd__a211o_1 _7133_ (.A1(_3364_),
    .A2(_3434_),
    .B1(_3437_),
    .C1(_3438_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3439_));
 sky130_fd_sc_hd__o21a_1 _7134_ (.A1(net295),
    .A2(_3360_),
    .B1(_3439_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0527_));
 sky130_fd_sc_hd__a221o_1 _7135_ (.A1(\i_tinyqv.cpu.instr_data[3][12] ),
    .A2(_3369_),
    .B1(_3370_),
    .B2(\i_tinyqv.cpu.instr_data[2][12] ),
    .C1(_3372_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3440_));
 sky130_fd_sc_hd__o221a_1 _7136_ (.A1(\i_tinyqv.cpu.instr_data[0][12] ),
    .A2(_3366_),
    .B1(_3368_),
    .B2(\i_tinyqv.cpu.instr_data[1][12] ),
    .C1(_3440_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3441_));
 sky130_fd_sc_hd__o21a_1 _7137_ (.A1(_3351_),
    .A2(_3398_),
    .B1(_1501_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3442_));
 sky130_fd_sc_hd__a221o_1 _7138_ (.A1(_1491_),
    .A2(_3423_),
    .B1(_3441_),
    .B2(_3364_),
    .C1(_3442_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3443_));
 sky130_fd_sc_hd__inv_2 _7139_ (.A(_3314_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3444_));
 sky130_fd_sc_hd__o211a_1 _7140_ (.A1(_3300_),
    .A2(_3444_),
    .B1(_3298_),
    .C1(_2120_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3445_));
 sky130_fd_sc_hd__and3_1 _7141_ (.A(_2155_),
    .B(_3299_),
    .C(_2120_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3446_));
 sky130_fd_sc_hd__o21ai_1 _7142_ (.A1(_2130_),
    .A2(_3337_),
    .B1(_3298_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3447_));
 sky130_fd_sc_hd__or3b_1 _7143_ (.A(_3445_),
    .B(_3446_),
    .C_N(_3447_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3448_));
 sky130_fd_sc_hd__or3_1 _7144_ (.A(_3362_),
    .B(_3443_),
    .C(_3448_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3449_));
 sky130_fd_sc_hd__o21a_1 _7145_ (.A1(\i_tinyqv.cpu.i_core.imm_lo[8] ),
    .A2(_3360_),
    .B1(_3449_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0528_));
 sky130_fd_sc_hd__a221o_1 _7146_ (.A1(\i_tinyqv.cpu.instr_data[3][13] ),
    .A2(_3369_),
    .B1(_3370_),
    .B2(\i_tinyqv.cpu.instr_data[2][13] ),
    .C1(_3372_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3450_));
 sky130_fd_sc_hd__o221a_1 _7147_ (.A1(\i_tinyqv.cpu.instr_data[0][13] ),
    .A2(_3366_),
    .B1(_3368_),
    .B2(\i_tinyqv.cpu.instr_data[1][13] ),
    .C1(_3450_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3451_));
 sky130_fd_sc_hd__nand2_1 _7148_ (.A(_3290_),
    .B(_3451_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3452_));
 sky130_fd_sc_hd__inv_2 _7149_ (.A(_3452_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3453_));
 sky130_fd_sc_hd__or3_2 _7150_ (.A(_1468_),
    .B(_1487_),
    .C(_2125_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3454_));
 sky130_fd_sc_hd__a21oi_1 _7151_ (.A1(_3309_),
    .A2(_3454_),
    .B1(_1507_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3455_));
 sky130_fd_sc_hd__a211o_1 _7152_ (.A1(_3299_),
    .A2(_2143_),
    .B1(_3448_),
    .C1(_3455_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3456_));
 sky130_fd_sc_hd__a221o_1 _7153_ (.A1(_2165_),
    .A2(_3398_),
    .B1(_3453_),
    .B2(_3315_),
    .C1(_3456_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3457_));
 sky130_fd_sc_hd__mux2_1 _7154_ (.A0(\i_tinyqv.cpu.i_core.imm_lo[9] ),
    .A1(_3457_),
    .S(_3396_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3458_));
 sky130_fd_sc_hd__clkbuf_1 _7155_ (.A(_3458_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0529_));
 sky130_fd_sc_hd__a221o_1 _7156_ (.A1(\i_tinyqv.cpu.instr_data[3][14] ),
    .A2(_3369_),
    .B1(_3370_),
    .B2(\i_tinyqv.cpu.instr_data[2][14] ),
    .C1(_3372_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3459_));
 sky130_fd_sc_hd__o221a_2 _7157_ (.A1(\i_tinyqv.cpu.instr_data[0][14] ),
    .A2(_3366_),
    .B1(_3368_),
    .B2(\i_tinyqv.cpu.instr_data[1][14] ),
    .C1(_3459_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3460_));
 sky130_fd_sc_hd__a221o_1 _7158_ (.A1(_1478_),
    .A2(_1514_),
    .B1(_3364_),
    .B2(_3460_),
    .C1(_3456_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3461_));
 sky130_fd_sc_hd__mux2_1 _7159_ (.A0(\i_tinyqv.cpu.i_core.imm_lo[10] ),
    .A1(_3461_),
    .S(_3396_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3462_));
 sky130_fd_sc_hd__clkbuf_1 _7160_ (.A(_3462_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0530_));
 sky130_fd_sc_hd__a221o_1 _7161_ (.A1(\i_tinyqv.cpu.instr_data[3][15] ),
    .A2(_3369_),
    .B1(_3370_),
    .B2(\i_tinyqv.cpu.instr_data[2][15] ),
    .C1(_3372_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3463_));
 sky130_fd_sc_hd__o221a_2 _7162_ (.A1(\i_tinyqv.cpu.instr_data[0][15] ),
    .A2(_3366_),
    .B1(_3368_),
    .B2(\i_tinyqv.cpu.instr_data[1][15] ),
    .C1(_3463_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3464_));
 sky130_fd_sc_hd__and2_1 _7163_ (.A(_1467_),
    .B(_3464_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3465_));
 sky130_fd_sc_hd__a31o_1 _7164_ (.A1(_2155_),
    .A2(_1466_),
    .A3(_3374_),
    .B1(_3465_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3466_));
 sky130_fd_sc_hd__or2_1 _7165_ (.A(_3334_),
    .B(_3319_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3467_));
 sky130_fd_sc_hd__mux2_1 _7166_ (.A0(_1510_),
    .A1(_3466_),
    .S(_3467_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3468_));
 sky130_fd_sc_hd__o21a_1 _7167_ (.A1(_1478_),
    .A2(_2143_),
    .B1(_3298_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3469_));
 sky130_fd_sc_hd__or3b_1 _7168_ (.A(_3445_),
    .B(_3469_),
    .C_N(_3447_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3470_));
 sky130_fd_sc_hd__or2_1 _7169_ (.A(_3446_),
    .B(_3470_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3471_));
 sky130_fd_sc_hd__or2_1 _7170_ (.A(_3455_),
    .B(_3471_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3472_));
 sky130_fd_sc_hd__a211o_1 _7171_ (.A1(_3364_),
    .A2(_3468_),
    .B1(_3472_),
    .C1(_3438_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3473_));
 sky130_fd_sc_hd__o21a_1 _7172_ (.A1(net296),
    .A2(_3360_),
    .B1(_3473_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0531_));
 sky130_fd_sc_hd__clkbuf_4 _7173_ (.A(_3359_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3474_));
 sky130_fd_sc_hd__a211o_1 _7174_ (.A1(_3364_),
    .A2(_3465_),
    .B1(_3472_),
    .C1(_3362_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3475_));
 sky130_fd_sc_hd__nand2_2 _7175_ (.A(_1467_),
    .B(_3315_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3476_));
 sky130_fd_sc_hd__a32o_1 _7176_ (.A1(_3328_),
    .A2(_3299_),
    .A3(_3476_),
    .B1(_3331_),
    .B2(_1460_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3477_));
 sky130_fd_sc_hd__o22a_1 _7177_ (.A1(net259),
    .A2(_3474_),
    .B1(_3475_),
    .B2(_3477_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0532_));
 sky130_fd_sc_hd__a32o_1 _7178_ (.A1(_3328_),
    .A2(_2123_),
    .A3(_3476_),
    .B1(_3331_),
    .B2(_2155_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3478_));
 sky130_fd_sc_hd__o22a_1 _7179_ (.A1(net257),
    .A2(_3474_),
    .B1(_3475_),
    .B2(_3478_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0533_));
 sky130_fd_sc_hd__a21o_1 _7180_ (.A1(_3315_),
    .A2(_3465_),
    .B1(_2140_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3479_));
 sky130_fd_sc_hd__a21o_1 _7181_ (.A1(_2124_),
    .A2(_3476_),
    .B1(_3479_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3480_));
 sky130_fd_sc_hd__or2_1 _7182_ (.A(_3290_),
    .B(_3455_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3481_));
 sky130_fd_sc_hd__a211o_1 _7183_ (.A1(_1491_),
    .A2(_3331_),
    .B1(_3471_),
    .C1(_3481_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3482_));
 sky130_fd_sc_hd__and3_1 _7184_ (.A(_3359_),
    .B(_3480_),
    .C(_3482_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3483_));
 sky130_fd_sc_hd__a21o_1 _7185_ (.A1(net231),
    .A2(_3438_),
    .B1(_3483_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0534_));
 sky130_fd_sc_hd__a21o_1 _7186_ (.A1(_1486_),
    .A2(_3476_),
    .B1(_3479_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3484_));
 sky130_fd_sc_hd__a211o_1 _7187_ (.A1(_3304_),
    .A2(_3331_),
    .B1(_3471_),
    .C1(_3481_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3485_));
 sky130_fd_sc_hd__and3_1 _7188_ (.A(_3359_),
    .B(_3484_),
    .C(_3485_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3486_));
 sky130_fd_sc_hd__a21o_1 _7189_ (.A1(net227),
    .A2(_3438_),
    .B1(_3486_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0535_));
 sky130_fd_sc_hd__nor2_1 _7190_ (.A(_1422_),
    .B(_1432_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3487_));
 sky130_fd_sc_hd__nor2_2 _7191_ (.A(_1504_),
    .B(_1461_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3488_));
 sky130_fd_sc_hd__nor2_1 _7192_ (.A(_3487_),
    .B(_3488_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3489_));
 sky130_fd_sc_hd__o211a_1 _7193_ (.A1(\i_tinyqv.cpu.instr_data[2][0] ),
    .A2(_1432_),
    .B1(_1418_),
    .C1(_3489_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3490_));
 sky130_fd_sc_hd__a221o_1 _7194_ (.A1(\i_tinyqv.cpu.instr_data[0][0] ),
    .A2(_3487_),
    .B1(_3488_),
    .B2(\i_tinyqv.cpu.instr_data[1][0] ),
    .C1(_3490_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3491_));
 sky130_fd_sc_hd__a21o_1 _7195_ (.A1(_3476_),
    .A2(_3491_),
    .B1(_3479_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3492_));
 sky130_fd_sc_hd__a211o_1 _7196_ (.A1(_3305_),
    .A2(_3331_),
    .B1(_3470_),
    .C1(_3481_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3493_));
 sky130_fd_sc_hd__and3_1 _7197_ (.A(_3359_),
    .B(_3492_),
    .C(_3493_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3494_));
 sky130_fd_sc_hd__a21o_1 _7198_ (.A1(net213),
    .A2(_3438_),
    .B1(_3494_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0536_));
 sky130_fd_sc_hd__o211a_1 _7199_ (.A1(\i_tinyqv.cpu.instr_data[2][1] ),
    .A2(_1432_),
    .B1(_1423_),
    .C1(_3489_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3495_));
 sky130_fd_sc_hd__a221o_1 _7200_ (.A1(\i_tinyqv.cpu.instr_data[0][1] ),
    .A2(_3487_),
    .B1(_3488_),
    .B2(\i_tinyqv.cpu.instr_data[1][1] ),
    .C1(_3495_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3496_));
 sky130_fd_sc_hd__and2_1 _7201_ (.A(_3290_),
    .B(_3496_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3497_));
 sky130_fd_sc_hd__o21a_1 _7202_ (.A1(_2126_),
    .A2(_3351_),
    .B1(_3298_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3498_));
 sky130_fd_sc_hd__or2_1 _7203_ (.A(_3470_),
    .B(_3498_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3499_));
 sky130_fd_sc_hd__a21o_1 _7204_ (.A1(_3364_),
    .A2(_3465_),
    .B1(_3499_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3500_));
 sky130_fd_sc_hd__a211o_1 _7205_ (.A1(_3476_),
    .A2(_3497_),
    .B1(_3500_),
    .C1(_3438_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3501_));
 sky130_fd_sc_hd__o21a_1 _7206_ (.A1(\i_tinyqv.cpu.imm[17] ),
    .A2(_3360_),
    .B1(_3501_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0537_));
 sky130_fd_sc_hd__o211a_1 _7207_ (.A1(\i_tinyqv.cpu.instr_data[2][2] ),
    .A2(_1432_),
    .B1(_1457_),
    .C1(_3489_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3502_));
 sky130_fd_sc_hd__a221o_1 _7208_ (.A1(\i_tinyqv.cpu.instr_data[0][2] ),
    .A2(_3487_),
    .B1(_3488_),
    .B2(\i_tinyqv.cpu.instr_data[1][2] ),
    .C1(_3502_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3503_));
 sky130_fd_sc_hd__and2_1 _7209_ (.A(_3290_),
    .B(_3503_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3504_));
 sky130_fd_sc_hd__a211o_1 _7210_ (.A1(_3476_),
    .A2(_3504_),
    .B1(_3500_),
    .C1(_3438_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3505_));
 sky130_fd_sc_hd__o21a_1 _7211_ (.A1(\i_tinyqv.cpu.imm[18] ),
    .A2(_3360_),
    .B1(_3505_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0538_));
 sky130_fd_sc_hd__o211a_1 _7212_ (.A1(\i_tinyqv.cpu.instr_data[2][3] ),
    .A2(_1432_),
    .B1(_1445_),
    .C1(_3489_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3506_));
 sky130_fd_sc_hd__a221o_1 _7213_ (.A1(\i_tinyqv.cpu.instr_data[0][3] ),
    .A2(_3487_),
    .B1(_3488_),
    .B2(\i_tinyqv.cpu.instr_data[1][3] ),
    .C1(_3506_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3507_));
 sky130_fd_sc_hd__a31o_1 _7214_ (.A1(_3328_),
    .A2(_3476_),
    .A3(_3507_),
    .B1(_3362_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3508_));
 sky130_fd_sc_hd__o22a_1 _7215_ (.A1(\i_tinyqv.cpu.imm[19] ),
    .A2(_3474_),
    .B1(_3500_),
    .B2(_3508_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0539_));
 sky130_fd_sc_hd__a21o_1 _7216_ (.A1(_3363_),
    .A2(_3464_),
    .B1(_3499_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3509_));
 sky130_fd_sc_hd__buf_2 _7217_ (.A(_3509_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3510_));
 sky130_fd_sc_hd__a31o_1 _7218_ (.A1(_3328_),
    .A2(_3330_),
    .A3(_3374_),
    .B1(_3362_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3511_));
 sky130_fd_sc_hd__o22a_1 _7219_ (.A1(\i_tinyqv.cpu.imm[20] ),
    .A2(_3474_),
    .B1(_3510_),
    .B2(_3511_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0540_));
 sky130_fd_sc_hd__a31o_1 _7220_ (.A1(_3328_),
    .A2(_3330_),
    .A3(_3384_),
    .B1(_3362_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3512_));
 sky130_fd_sc_hd__o22a_1 _7221_ (.A1(\i_tinyqv.cpu.imm[21] ),
    .A2(_3474_),
    .B1(_3510_),
    .B2(_3512_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0541_));
 sky130_fd_sc_hd__a311o_1 _7222_ (.A1(_3328_),
    .A2(_3330_),
    .A3(_3390_),
    .B1(_3510_),
    .C1(_3362_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3513_));
 sky130_fd_sc_hd__o21a_1 _7223_ (.A1(\i_tinyqv.cpu.imm[22] ),
    .A2(_3360_),
    .B1(_3513_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0542_));
 sky130_fd_sc_hd__nand2_1 _7224_ (.A(_3289_),
    .B(_3402_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3514_));
 sky130_fd_sc_hd__o21ba_1 _7225_ (.A1(_3315_),
    .A2(_3514_),
    .B1_N(_3510_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3515_));
 sky130_fd_sc_hd__nor2_1 _7226_ (.A(\i_tinyqv.cpu.imm[23] ),
    .B(_3359_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3516_));
 sky130_fd_sc_hd__a21oi_1 _7227_ (.A1(_3474_),
    .A2(_3515_),
    .B1(_3516_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0543_));
 sky130_fd_sc_hd__a31o_1 _7228_ (.A1(_3328_),
    .A2(_3330_),
    .A3(_3408_),
    .B1(_3510_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3517_));
 sky130_fd_sc_hd__mux2_1 _7229_ (.A0(\i_tinyqv.cpu.imm[24] ),
    .A1(_3517_),
    .S(_3396_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3518_));
 sky130_fd_sc_hd__clkbuf_1 _7230_ (.A(_3518_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0544_));
 sky130_fd_sc_hd__a31o_1 _7231_ (.A1(_3291_),
    .A2(_3330_),
    .A3(_3418_),
    .B1(_3510_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3519_));
 sky130_fd_sc_hd__mux2_1 _7232_ (.A0(\i_tinyqv.cpu.imm[25] ),
    .A1(_3519_),
    .S(_3396_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3520_));
 sky130_fd_sc_hd__clkbuf_1 _7233_ (.A(_3520_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0545_));
 sky130_fd_sc_hd__o21ai_1 _7234_ (.A1(_3315_),
    .A2(_3428_),
    .B1(_3359_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3521_));
 sky130_fd_sc_hd__o22a_1 _7235_ (.A1(net190),
    .A2(_3474_),
    .B1(_3510_),
    .B2(_3521_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0546_));
 sky130_fd_sc_hd__a31o_1 _7236_ (.A1(_3291_),
    .A2(_3330_),
    .A3(_3434_),
    .B1(_3510_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3522_));
 sky130_fd_sc_hd__mux2_1 _7237_ (.A0(\i_tinyqv.cpu.imm[27] ),
    .A1(_3522_),
    .S(_3396_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3523_));
 sky130_fd_sc_hd__clkbuf_1 _7238_ (.A(_3523_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0547_));
 sky130_fd_sc_hd__a31o_1 _7239_ (.A1(_3291_),
    .A2(_3330_),
    .A3(_3441_),
    .B1(_3510_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3524_));
 sky130_fd_sc_hd__mux2_1 _7240_ (.A0(\i_tinyqv.cpu.imm[28] ),
    .A1(_3524_),
    .S(_3396_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3525_));
 sky130_fd_sc_hd__clkbuf_1 _7241_ (.A(_3525_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0548_));
 sky130_fd_sc_hd__a211o_1 _7242_ (.A1(_3330_),
    .A2(_3453_),
    .B1(_3510_),
    .C1(_3438_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3526_));
 sky130_fd_sc_hd__o21a_1 _7243_ (.A1(net146),
    .A2(_3360_),
    .B1(_3526_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0549_));
 sky130_fd_sc_hd__a31o_1 _7244_ (.A1(_3291_),
    .A2(_3330_),
    .A3(_3460_),
    .B1(_3509_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3527_));
 sky130_fd_sc_hd__mux2_1 _7245_ (.A0(net284),
    .A1(_3527_),
    .S(_3395_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3528_));
 sky130_fd_sc_hd__clkbuf_1 _7246_ (.A(_3528_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0550_));
 sky130_fd_sc_hd__a211o_1 _7247_ (.A1(_3328_),
    .A2(_3464_),
    .B1(_3499_),
    .C1(_3438_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3529_));
 sky130_fd_sc_hd__o21a_1 _7248_ (.A1(net135),
    .A2(_3360_),
    .B1(_3529_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0551_));
 sky130_fd_sc_hd__nor2_1 _7249_ (.A(_2140_),
    .B(_1466_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3530_));
 sky130_fd_sc_hd__o211a_1 _7250_ (.A1(_3304_),
    .A2(_3315_),
    .B1(_3530_),
    .C1(_1493_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3531_));
 sky130_fd_sc_hd__and2_1 _7251_ (.A(_3325_),
    .B(_3427_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3532_));
 sky130_fd_sc_hd__nor2_1 _7252_ (.A(_3335_),
    .B(_3532_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3533_));
 sky130_fd_sc_hd__a22o_1 _7253_ (.A1(_2123_),
    .A2(_3335_),
    .B1(_3533_),
    .B2(_3299_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3534_));
 sky130_fd_sc_hd__o31a_1 _7254_ (.A1(_1507_),
    .A2(_3300_),
    .A3(_3314_),
    .B1(_2121_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3535_));
 sky130_fd_sc_hd__a21boi_1 _7255_ (.A1(_1456_),
    .A2(_3301_),
    .B1_N(_3535_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3536_));
 sky130_fd_sc_hd__a211o_1 _7256_ (.A1(_3531_),
    .A2(_3534_),
    .B1(_3536_),
    .C1(_2129_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3537_));
 sky130_fd_sc_hd__mux2_1 _7257_ (.A0(net69),
    .A1(_3537_),
    .S(_3395_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3538_));
 sky130_fd_sc_hd__clkbuf_1 _7258_ (.A(_3538_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0552_));
 sky130_fd_sc_hd__nand2_1 _7259_ (.A(_3334_),
    .B(_3301_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3539_));
 sky130_fd_sc_hd__or2_1 _7260_ (.A(_2124_),
    .B(_3467_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3540_));
 sky130_fd_sc_hd__o311a_1 _7261_ (.A1(_2123_),
    .A2(_3335_),
    .A3(_3532_),
    .B1(_3540_),
    .C1(_3531_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3541_));
 sky130_fd_sc_hd__a311o_2 _7262_ (.A1(_3287_),
    .A2(_3535_),
    .A3(_3539_),
    .B1(_3541_),
    .C1(_2131_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3542_));
 sky130_fd_sc_hd__mux2_1 _7263_ (.A0(_0656_),
    .A1(_3542_),
    .S(_3395_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3543_));
 sky130_fd_sc_hd__clkbuf_1 _7264_ (.A(_3543_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0553_));
 sky130_fd_sc_hd__a21bo_1 _7265_ (.A1(_2124_),
    .A2(_3533_),
    .B1_N(_3540_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3544_));
 sky130_fd_sc_hd__or2_1 _7266_ (.A(_3304_),
    .B(_3539_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3545_));
 sky130_fd_sc_hd__a221o_2 _7267_ (.A1(_3531_),
    .A2(_3544_),
    .B1(_3545_),
    .B2(_2121_),
    .C1(_3337_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3546_));
 sky130_fd_sc_hd__mux2_1 _7268_ (.A0(_1030_),
    .A1(_3546_),
    .S(_3395_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3547_));
 sky130_fd_sc_hd__clkbuf_1 _7269_ (.A(_3547_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0554_));
 sky130_fd_sc_hd__a21o_1 _7270_ (.A1(_1473_),
    .A2(_3299_),
    .B1(_3304_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3548_));
 sky130_fd_sc_hd__a21o_1 _7271_ (.A1(_3460_),
    .A2(_3548_),
    .B1(_3532_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3549_));
 sky130_fd_sc_hd__a21bo_1 _7272_ (.A1(_2165_),
    .A2(_3288_),
    .B1_N(_3545_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3550_));
 sky130_fd_sc_hd__a32o_1 _7273_ (.A1(_3467_),
    .A2(_3531_),
    .A3(_3549_),
    .B1(_3550_),
    .B2(_2121_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3551_));
 sky130_fd_sc_hd__or3_1 _7274_ (.A(_2131_),
    .B(_3362_),
    .C(_3551_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3552_));
 sky130_fd_sc_hd__o21a_1 _7275_ (.A1(net243),
    .A2(_3474_),
    .B1(_3552_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0555_));
 sky130_fd_sc_hd__nor2_1 _7276_ (.A(_1473_),
    .B(_1493_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3553_));
 sky130_fd_sc_hd__inv_2 _7277_ (.A(_3553_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3554_));
 sky130_fd_sc_hd__nor2_1 _7278_ (.A(_3293_),
    .B(_3322_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3555_));
 sky130_fd_sc_hd__nor2_2 _7279_ (.A(_3289_),
    .B(_3337_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3556_));
 sky130_fd_sc_hd__a32o_1 _7280_ (.A1(_2165_),
    .A2(_3555_),
    .A3(_3556_),
    .B1(_3337_),
    .B2(_2123_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3557_));
 sky130_fd_sc_hd__a31o_1 _7281_ (.A1(_3291_),
    .A2(_3299_),
    .A3(_3554_),
    .B1(_3557_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3558_));
 sky130_fd_sc_hd__mux2_1 _7282_ (.A0(\i_tinyqv.cpu.i_core.mem_op[0] ),
    .A1(_3558_),
    .S(_3395_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3559_));
 sky130_fd_sc_hd__clkbuf_1 _7283_ (.A(_3559_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0556_));
 sky130_fd_sc_hd__o21ai_1 _7284_ (.A1(_2140_),
    .A2(_1473_),
    .B1(_3555_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3560_));
 sky130_fd_sc_hd__mux2_1 _7285_ (.A0(\i_tinyqv.cpu.i_core.mem_op[1] ),
    .A1(_3560_),
    .S(_3395_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3561_));
 sky130_fd_sc_hd__clkbuf_1 _7286_ (.A(_3561_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0557_));
 sky130_fd_sc_hd__and4_1 _7287_ (.A(_2123_),
    .B(_2124_),
    .C(_1507_),
    .D(_3320_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3562_));
 sky130_fd_sc_hd__a21o_1 _7288_ (.A1(_3299_),
    .A2(_3553_),
    .B1(_3562_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3563_));
 sky130_fd_sc_hd__inv_2 _7289_ (.A(_3563_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3564_));
 sky130_fd_sc_hd__a21oi_1 _7290_ (.A1(_3305_),
    .A2(_2165_),
    .B1(_3287_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3565_));
 sky130_fd_sc_hd__and3_1 _7291_ (.A(_3555_),
    .B(_3556_),
    .C(_3565_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3566_));
 sky130_fd_sc_hd__a31o_1 _7292_ (.A1(_3291_),
    .A2(_2124_),
    .A3(_3564_),
    .B1(_3566_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3567_));
 sky130_fd_sc_hd__mux2_1 _7293_ (.A0(\i_tinyqv.cpu.i_core.mem_op[2] ),
    .A1(_3567_),
    .S(_3395_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3568_));
 sky130_fd_sc_hd__clkbuf_1 _7294_ (.A(_3568_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0558_));
 sky130_fd_sc_hd__nor2_1 _7295_ (.A(_1483_),
    .B(_2122_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3569_));
 sky130_fd_sc_hd__or4_1 _7296_ (.A(_2129_),
    .B(_2131_),
    .C(_2142_),
    .D(_3569_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3570_));
 sky130_fd_sc_hd__or3_1 _7297_ (.A(_2121_),
    .B(_3337_),
    .C(_3353_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3571_));
 sky130_fd_sc_hd__or3_2 _7298_ (.A(_3341_),
    .B(_3570_),
    .C(_3571_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3572_));
 sky130_fd_sc_hd__or2_1 _7299_ (.A(_2143_),
    .B(_3351_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3573_));
 sky130_fd_sc_hd__a221o_1 _7300_ (.A1(_3291_),
    .A2(_1486_),
    .B1(_1510_),
    .B2(_3572_),
    .C1(_3573_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3574_));
 sky130_fd_sc_hd__mux2_1 _7301_ (.A0(_0627_),
    .A1(_3574_),
    .S(_3395_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3575_));
 sky130_fd_sc_hd__clkbuf_1 _7302_ (.A(_3575_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0559_));
 sky130_fd_sc_hd__or3_1 _7303_ (.A(_1426_),
    .B(_2123_),
    .C(_3321_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3576_));
 sky130_fd_sc_hd__or4b_1 _7304_ (.A(_3289_),
    .B(_2126_),
    .C(_3349_),
    .D_N(_3576_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3577_));
 sky130_fd_sc_hd__a211o_1 _7305_ (.A1(_1514_),
    .A2(_3572_),
    .B1(_3573_),
    .C1(_3577_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3578_));
 sky130_fd_sc_hd__o211a_1 _7306_ (.A1(_2140_),
    .A2(_3491_),
    .B1(_3578_),
    .C1(_3359_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3579_));
 sky130_fd_sc_hd__a21o_1 _7307_ (.A1(_0624_),
    .A2(_3438_),
    .B1(_3579_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0560_));
 sky130_fd_sc_hd__nor2_1 _7308_ (.A(_1473_),
    .B(_3321_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3580_));
 sky130_fd_sc_hd__a221o_1 _7309_ (.A1(_1468_),
    .A2(_3580_),
    .B1(_3572_),
    .B2(_1501_),
    .C1(_3497_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3581_));
 sky130_fd_sc_hd__mux2_1 _7310_ (.A0(_0625_),
    .A1(_3581_),
    .S(_3395_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3582_));
 sky130_fd_sc_hd__clkbuf_1 _7311_ (.A(_3582_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0561_));
 sky130_fd_sc_hd__o21a_1 _7312_ (.A1(_2165_),
    .A2(_3571_),
    .B1(_3572_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3583_));
 sky130_fd_sc_hd__or3_1 _7313_ (.A(_3362_),
    .B(_3504_),
    .C(_3583_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3584_));
 sky130_fd_sc_hd__o21a_1 _7314_ (.A1(net324),
    .A2(_3474_),
    .B1(_3584_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0562_));
 sky130_fd_sc_hd__xor2_1 _7315_ (.A(_0662_),
    .B(\i_tinyqv.cpu.mem_op_increment_reg ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3585_));
 sky130_fd_sc_hd__nand2_1 _7316_ (.A(_3313_),
    .B(_3454_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3586_));
 sky130_fd_sc_hd__a221o_1 _7317_ (.A1(_3290_),
    .A2(_3374_),
    .B1(_3556_),
    .B2(_3586_),
    .C1(_2149_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3587_));
 sky130_fd_sc_hd__o21a_1 _7318_ (.A1(_2147_),
    .A2(_3585_),
    .B1(_3587_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3588_));
 sky130_fd_sc_hd__mux2_1 _7319_ (.A0(_3588_),
    .A1(_0662_),
    .S(_2153_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3589_));
 sky130_fd_sc_hd__clkbuf_1 _7320_ (.A(_3589_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0563_));
 sky130_fd_sc_hd__a32o_1 _7321_ (.A1(_2155_),
    .A2(_3454_),
    .A3(_3556_),
    .B1(_3384_),
    .B2(_3290_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3590_));
 sky130_fd_sc_hd__a21oi_1 _7322_ (.A1(_0662_),
    .A2(\i_tinyqv.cpu.mem_op_increment_reg ),
    .B1(_0663_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3591_));
 sky130_fd_sc_hd__a21oi_1 _7323_ (.A1(\i_tinyqv.cpu.mem_op_increment_reg ),
    .A2(_0711_),
    .B1(_3591_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3592_));
 sky130_fd_sc_hd__mux2_1 _7324_ (.A0(_3590_),
    .A1(_3592_),
    .S(_2149_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3593_));
 sky130_fd_sc_hd__mux2_1 _7325_ (.A0(_3593_),
    .A1(_0663_),
    .S(_2153_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3594_));
 sky130_fd_sc_hd__clkbuf_1 _7326_ (.A(_3594_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0564_));
 sky130_fd_sc_hd__and3_1 _7327_ (.A(_0660_),
    .B(\i_tinyqv.cpu.mem_op_increment_reg ),
    .C(_0711_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3595_));
 sky130_fd_sc_hd__a21oi_1 _7328_ (.A1(\i_tinyqv.cpu.mem_op_increment_reg ),
    .A2(_0711_),
    .B1(_0660_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3596_));
 sky130_fd_sc_hd__nor2_1 _7329_ (.A(_3595_),
    .B(_3596_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3597_));
 sky130_fd_sc_hd__a32o_1 _7330_ (.A1(_1491_),
    .A2(_3454_),
    .A3(_3556_),
    .B1(_3390_),
    .B2(_3290_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3598_));
 sky130_fd_sc_hd__mux2_1 _7331_ (.A0(_3597_),
    .A1(_3598_),
    .S(_2147_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3599_));
 sky130_fd_sc_hd__mux2_1 _7332_ (.A0(_3599_),
    .A1(_0660_),
    .S(_2153_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3600_));
 sky130_fd_sc_hd__clkbuf_1 _7333_ (.A(_3600_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0565_));
 sky130_fd_sc_hd__xor2_1 _7334_ (.A(_0661_),
    .B(_3595_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3601_));
 sky130_fd_sc_hd__a211o_1 _7335_ (.A1(_1426_),
    .A2(_2125_),
    .B1(_1487_),
    .C1(_3304_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3602_));
 sky130_fd_sc_hd__a21bo_1 _7336_ (.A1(_3556_),
    .A2(_3602_),
    .B1_N(_3514_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3603_));
 sky130_fd_sc_hd__mux2_1 _7337_ (.A0(_3601_),
    .A1(_3603_),
    .S(_2147_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3604_));
 sky130_fd_sc_hd__mux2_1 _7338_ (.A0(_3604_),
    .A1(_0661_),
    .S(_2153_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3605_));
 sky130_fd_sc_hd__clkbuf_1 _7339_ (.A(_3605_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0566_));
 sky130_fd_sc_hd__o211a_1 _7340_ (.A1(\i_tinyqv.cpu.instr_len[1] ),
    .A2(_3282_),
    .B1(_3312_),
    .C1(_1753_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0567_));
 sky130_fd_sc_hd__a211o_1 _7341_ (.A1(net196),
    .A2(_3295_),
    .B1(_3333_),
    .C1(_2067_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0568_));
 sky130_fd_sc_hd__a221o_1 _7342_ (.A1(_1510_),
    .A2(_2143_),
    .B1(_3351_),
    .B2(_1460_),
    .C1(_3328_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3606_));
 sky130_fd_sc_hd__o211ai_1 _7343_ (.A1(_2140_),
    .A2(_3563_),
    .B1(_3606_),
    .C1(_3282_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3607_));
 sky130_fd_sc_hd__mux2_1 _7344_ (.A0(_2147_),
    .A1(_2152_),
    .S(\i_tinyqv.cpu.additional_mem_ops[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3608_));
 sky130_fd_sc_hd__a21oi_1 _7345_ (.A1(_3607_),
    .A2(_3608_),
    .B1(_2067_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0569_));
 sky130_fd_sc_hd__a221o_1 _7346_ (.A1(_1514_),
    .A2(_2143_),
    .B1(_3351_),
    .B2(_2155_),
    .C1(_2149_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3609_));
 sky130_fd_sc_hd__a31o_1 _7347_ (.A1(_3291_),
    .A2(_2124_),
    .A3(_3563_),
    .B1(_3609_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3610_));
 sky130_fd_sc_hd__nor2_1 _7348_ (.A(\i_tinyqv.cpu.additional_mem_ops[1] ),
    .B(\i_tinyqv.cpu.additional_mem_ops[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3611_));
 sky130_fd_sc_hd__and2_1 _7349_ (.A(\i_tinyqv.cpu.additional_mem_ops[1] ),
    .B(\i_tinyqv.cpu.additional_mem_ops[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3612_));
 sky130_fd_sc_hd__or3_1 _7350_ (.A(_1439_),
    .B(_3611_),
    .C(_3612_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3613_));
 sky130_fd_sc_hd__a21bo_1 _7351_ (.A1(_3610_),
    .A2(_3613_),
    .B1_N(_2152_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3614_));
 sky130_fd_sc_hd__o211a_1 _7352_ (.A1(net242),
    .A2(_2152_),
    .B1(_3614_),
    .C1(_1753_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0570_));
 sky130_fd_sc_hd__o21ai_1 _7353_ (.A1(_1439_),
    .A2(_3611_),
    .B1(_2152_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3615_));
 sky130_fd_sc_hd__a22o_1 _7354_ (.A1(_1501_),
    .A2(_2143_),
    .B1(_3351_),
    .B2(_1491_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3616_));
 sky130_fd_sc_hd__a32o_1 _7355_ (.A1(net154),
    .A2(_2049_),
    .A3(_3615_),
    .B1(_3616_),
    .B2(_3359_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0571_));
 sky130_fd_sc_hd__nand2_1 _7356_ (.A(_2079_),
    .B(_3562_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3617_));
 sky130_fd_sc_hd__o22a_1 _7357_ (.A1(\i_tinyqv.cpu.mem_op_increment_reg ),
    .A2(_3474_),
    .B1(_3617_),
    .B2(_3312_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0572_));
 sky130_fd_sc_hd__nand2_1 _7358_ (.A(_1405_),
    .B(_2147_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3618_));
 sky130_fd_sc_hd__o21ai_1 _7359_ (.A1(_2993_),
    .A2(_1443_),
    .B1(_2147_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3619_));
 sky130_fd_sc_hd__nand2_1 _7360_ (.A(net127),
    .B(_3619_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3620_));
 sky130_fd_sc_hd__a21oi_1 _7361_ (.A1(_3618_),
    .A2(_3620_),
    .B1(_2067_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0573_));
 sky130_fd_sc_hd__nand2_1 _7362_ (.A(_2150_),
    .B(_1515_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3621_));
 sky130_fd_sc_hd__o2bb2a_1 _7363_ (.A1_N(_3619_),
    .A2_N(_3618_),
    .B1(_3621_),
    .B2(_2993_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3622_));
 sky130_fd_sc_hd__a311oi_1 _7364_ (.A1(_1410_),
    .A2(_3619_),
    .A3(_3618_),
    .B1(_3622_),
    .C1(_2066_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0574_));
 sky130_fd_sc_hd__and3_1 _7365_ (.A(_2079_),
    .B(_1528_),
    .C(_2995_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3623_));
 sky130_fd_sc_hd__clkbuf_1 _7366_ (.A(_3623_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0575_));
 sky130_fd_sc_hd__nand2_8 _7367_ (.A(net155),
    .B(_1709_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3624_));
 sky130_fd_sc_hd__nand2_4 _7368_ (.A(_2732_),
    .B(_3624_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3625_));
 sky130_fd_sc_hd__a21oi_1 _7369_ (.A1(_0884_),
    .A2(\i_tinyqv.cpu.instr_write_offset[3] ),
    .B1(\i_tinyqv.cpu.instr_data_start[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3626_));
 sky130_fd_sc_hd__a31o_1 _7370_ (.A1(\i_tinyqv.cpu.instr_data_start[4] ),
    .A2(_0884_),
    .A3(\i_tinyqv.cpu.instr_write_offset[3] ),
    .B1(_3010_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3627_));
 sky130_fd_sc_hd__o221a_1 _7371_ (.A1(_3239_),
    .A2(_3045_),
    .B1(_3626_),
    .B2(_3627_),
    .C1(_2681_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3628_));
 sky130_fd_sc_hd__o21ai_1 _7372_ (.A1(\i_tinyqv.cpu.data_addr[4] ),
    .A2(_2682_),
    .B1(_3005_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3629_));
 sky130_fd_sc_hd__nor2_1 _7373_ (.A(_3628_),
    .B(_3629_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3630_));
 sky130_fd_sc_hd__o21a_1 _7374_ (.A1(net310),
    .A2(_3624_),
    .B1(_2733_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3631_));
 sky130_fd_sc_hd__o22a_1 _7375_ (.A1(net151),
    .A2(_3625_),
    .B1(_3630_),
    .B2(_3631_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0576_));
 sky130_fd_sc_hd__clkbuf_4 _7376_ (.A(\i_tinyqv.cpu.was_early_branch ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3632_));
 sky130_fd_sc_hd__a31o_1 _7377_ (.A1(\i_tinyqv.cpu.instr_data_start[4] ),
    .A2(_0884_),
    .A3(\i_tinyqv.cpu.instr_write_offset[3] ),
    .B1(\i_tinyqv.cpu.instr_data_start[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3633_));
 sky130_fd_sc_hd__and4_2 _7378_ (.A(\i_tinyqv.cpu.instr_data_start[5] ),
    .B(\i_tinyqv.cpu.instr_data_start[4] ),
    .C(_0884_),
    .D(\i_tinyqv.cpu.instr_write_offset[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3634_));
 sky130_fd_sc_hd__nor2_1 _7379_ (.A(_3010_),
    .B(_3634_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3635_));
 sky130_fd_sc_hd__a221o_1 _7380_ (.A1(_3632_),
    .A2(_3056_),
    .B1(_3633_),
    .B2(_3635_),
    .C1(_2877_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3636_));
 sky130_fd_sc_hd__o211a_1 _7381_ (.A1(net299),
    .A2(_2682_),
    .B1(_3004_),
    .C1(_3636_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3637_));
 sky130_fd_sc_hd__o21a_1 _7382_ (.A1(net93),
    .A2(_3624_),
    .B1(_2733_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3638_));
 sky130_fd_sc_hd__o22a_1 _7383_ (.A1(net305),
    .A2(_3625_),
    .B1(_3637_),
    .B2(_3638_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0577_));
 sky130_fd_sc_hd__nor2_1 _7384_ (.A(_0883_),
    .B(_3634_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3639_));
 sky130_fd_sc_hd__a21o_1 _7385_ (.A1(_0883_),
    .A2(_3634_),
    .B1(\i_tinyqv.cpu.was_early_branch ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3640_));
 sky130_fd_sc_hd__o22a_1 _7386_ (.A1(_3239_),
    .A2(_3067_),
    .B1(_3639_),
    .B2(_3640_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3641_));
 sky130_fd_sc_hd__a21oi_1 _7387_ (.A1(_3012_),
    .A2(_3641_),
    .B1(_2732_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3642_));
 sky130_fd_sc_hd__o21a_1 _7388_ (.A1(\i_tinyqv.cpu.data_addr[6] ),
    .A2(_2682_),
    .B1(_3642_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3643_));
 sky130_fd_sc_hd__o21a_1 _7389_ (.A1(net126),
    .A2(_3624_),
    .B1(_2733_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3644_));
 sky130_fd_sc_hd__o22a_1 _7390_ (.A1(net89),
    .A2(_3625_),
    .B1(_3643_),
    .B2(_3644_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0578_));
 sky130_fd_sc_hd__and3_1 _7391_ (.A(\i_tinyqv.cpu.instr_data_start[7] ),
    .B(_0883_),
    .C(_3634_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3645_));
 sky130_fd_sc_hd__a21oi_1 _7392_ (.A1(_0883_),
    .A2(_3634_),
    .B1(\i_tinyqv.cpu.instr_data_start[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3646_));
 sky130_fd_sc_hd__o21a_1 _7393_ (.A1(_3645_),
    .A2(_3646_),
    .B1(_3239_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3647_));
 sky130_fd_sc_hd__a211oi_1 _7394_ (.A1(_3017_),
    .A2(_3080_),
    .B1(_3647_),
    .C1(_2877_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3648_));
 sky130_fd_sc_hd__a211o_1 _7395_ (.A1(net297),
    .A2(_2878_),
    .B1(_2733_),
    .C1(_3648_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3649_));
 sky130_fd_sc_hd__o221a_1 _7396_ (.A1(net95),
    .A2(_3624_),
    .B1(_3625_),
    .B2(net302),
    .C1(_3649_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0579_));
 sky130_fd_sc_hd__or2_1 _7397_ (.A(\i_tinyqv.cpu.instr_data_start[8] ),
    .B(_3645_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3650_));
 sky130_fd_sc_hd__and2_1 _7398_ (.A(\i_tinyqv.cpu.instr_data_start[8] ),
    .B(_3645_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3651_));
 sky130_fd_sc_hd__nor2_1 _7399_ (.A(_3017_),
    .B(_3651_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3652_));
 sky130_fd_sc_hd__a221o_1 _7400_ (.A1(_3017_),
    .A2(_3088_),
    .B1(_3650_),
    .B2(_3652_),
    .C1(_2878_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3653_));
 sky130_fd_sc_hd__o21a_1 _7401_ (.A1(\i_tinyqv.cpu.data_addr[8] ),
    .A2(_2682_),
    .B1(_3005_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3654_));
 sky130_fd_sc_hd__mux2_1 _7402_ (.A0(\i_tinyqv.mem.q_ctrl.addr[4] ),
    .A1(net312),
    .S(_3624_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3655_));
 sky130_fd_sc_hd__a22o_1 _7403_ (.A1(_3653_),
    .A2(_3654_),
    .B1(_3655_),
    .B2(_2733_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0580_));
 sky130_fd_sc_hd__or2_1 _7404_ (.A(_0882_),
    .B(_3651_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3656_));
 sky130_fd_sc_hd__a21oi_1 _7405_ (.A1(_0882_),
    .A2(_3651_),
    .B1(_3010_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3657_));
 sky130_fd_sc_hd__a221o_1 _7406_ (.A1(_3632_),
    .A2(_3099_),
    .B1(_3656_),
    .B2(_3657_),
    .C1(_2877_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3658_));
 sky130_fd_sc_hd__o211a_1 _7407_ (.A1(\i_tinyqv.cpu.data_addr[9] ),
    .A2(_3012_),
    .B1(_3004_),
    .C1(_3658_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3659_));
 sky130_fd_sc_hd__a221o_1 _7408_ (.A1(net305),
    .A2(_3007_),
    .B1(_3009_),
    .B2(net187),
    .C1(_3659_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0581_));
 sky130_fd_sc_hd__nor2_1 _7409_ (.A(_3239_),
    .B(_3108_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3660_));
 sky130_fd_sc_hd__and3_1 _7410_ (.A(\i_tinyqv.cpu.instr_data_start[10] ),
    .B(_0882_),
    .C(_3651_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3661_));
 sky130_fd_sc_hd__a21oi_1 _7411_ (.A1(_0882_),
    .A2(_3651_),
    .B1(\i_tinyqv.cpu.instr_data_start[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3662_));
 sky130_fd_sc_hd__nor3_1 _7412_ (.A(_3010_),
    .B(_3661_),
    .C(_3662_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3663_));
 sky130_fd_sc_hd__o31a_1 _7413_ (.A1(_2877_),
    .A2(_3660_),
    .A3(_3663_),
    .B1(_3004_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3664_));
 sky130_fd_sc_hd__o21a_1 _7414_ (.A1(net298),
    .A2(_2682_),
    .B1(_3664_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3665_));
 sky130_fd_sc_hd__a221o_1 _7415_ (.A1(net89),
    .A2(_3007_),
    .B1(_3009_),
    .B2(net317),
    .C1(_3665_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0582_));
 sky130_fd_sc_hd__or2_1 _7416_ (.A(\i_tinyqv.cpu.instr_data_start[11] ),
    .B(_3661_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3666_));
 sky130_fd_sc_hd__and2_1 _7417_ (.A(\i_tinyqv.cpu.instr_data_start[11] ),
    .B(_3661_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3667_));
 sky130_fd_sc_hd__nor2_1 _7418_ (.A(_3010_),
    .B(_3667_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3668_));
 sky130_fd_sc_hd__a221o_1 _7419_ (.A1(_3632_),
    .A2(_3119_),
    .B1(_3666_),
    .B2(_3668_),
    .C1(_2877_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3669_));
 sky130_fd_sc_hd__o211a_1 _7420_ (.A1(net96),
    .A2(_3012_),
    .B1(_3004_),
    .C1(_3669_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3670_));
 sky130_fd_sc_hd__a221o_1 _7421_ (.A1(net302),
    .A2(_3007_),
    .B1(_3009_),
    .B2(net303),
    .C1(_3670_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0583_));
 sky130_fd_sc_hd__xor2_1 _7422_ (.A(_0726_),
    .B(_3667_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3671_));
 sky130_fd_sc_hd__nand2_1 _7423_ (.A(_3632_),
    .B(_3129_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3672_));
 sky130_fd_sc_hd__o211a_1 _7424_ (.A1(_3632_),
    .A2(_3671_),
    .B1(_3672_),
    .C1(_2681_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3673_));
 sky130_fd_sc_hd__a211o_1 _7425_ (.A1(\i_tinyqv.cpu.data_addr[12] ),
    .A2(_2878_),
    .B1(_2732_),
    .C1(_3673_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3674_));
 sky130_fd_sc_hd__o221a_1 _7426_ (.A1(net153),
    .A2(_3624_),
    .B1(_3625_),
    .B2(net147),
    .C1(_3674_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0584_));
 sky130_fd_sc_hd__a31o_1 _7427_ (.A1(_0726_),
    .A2(\i_tinyqv.cpu.instr_data_start[11] ),
    .A3(_3661_),
    .B1(\i_tinyqv.cpu.instr_data_start[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3675_));
 sky130_fd_sc_hd__and3_1 _7428_ (.A(\i_tinyqv.cpu.instr_data_start[13] ),
    .B(_0726_),
    .C(_3667_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3676_));
 sky130_fd_sc_hd__nor2_1 _7429_ (.A(\i_tinyqv.cpu.was_early_branch ),
    .B(_3676_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3677_));
 sky130_fd_sc_hd__a221o_1 _7430_ (.A1(_3632_),
    .A2(_3141_),
    .B1(_3675_),
    .B2(_3677_),
    .C1(_2877_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3678_));
 sky130_fd_sc_hd__o211a_1 _7431_ (.A1(net181),
    .A2(_3012_),
    .B1(_3004_),
    .C1(_3678_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3679_));
 sky130_fd_sc_hd__a221o_1 _7432_ (.A1(net187),
    .A2(_3007_),
    .B1(_3009_),
    .B2(net304),
    .C1(_3679_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0585_));
 sky130_fd_sc_hd__or2_1 _7433_ (.A(\i_tinyqv.cpu.instr_data_start[14] ),
    .B(_3676_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3680_));
 sky130_fd_sc_hd__and2_1 _7434_ (.A(\i_tinyqv.cpu.instr_data_start[14] ),
    .B(_3676_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3681_));
 sky130_fd_sc_hd__nor2_1 _7435_ (.A(_3010_),
    .B(_3681_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3682_));
 sky130_fd_sc_hd__a22o_1 _7436_ (.A1(_3632_),
    .A2(_3150_),
    .B1(_3680_),
    .B2(_3682_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3683_));
 sky130_fd_sc_hd__mux2_1 _7437_ (.A0(net111),
    .A1(_3683_),
    .S(_3012_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3684_));
 sky130_fd_sc_hd__a22o_1 _7438_ (.A1(\i_tinyqv.mem.q_ctrl.addr[10] ),
    .A2(_3007_),
    .B1(_3008_),
    .B2(net315),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3685_));
 sky130_fd_sc_hd__a21o_1 _7439_ (.A1(_3005_),
    .A2(_3684_),
    .B1(_3685_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0586_));
 sky130_fd_sc_hd__or2_1 _7440_ (.A(_0881_),
    .B(_3681_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3686_));
 sky130_fd_sc_hd__a21oi_1 _7441_ (.A1(_0881_),
    .A2(_3681_),
    .B1(_3010_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3687_));
 sky130_fd_sc_hd__a221o_1 _7442_ (.A1(_3632_),
    .A2(_3158_),
    .B1(_3686_),
    .B2(_3687_),
    .C1(_2877_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3688_));
 sky130_fd_sc_hd__o211a_1 _7443_ (.A1(net173),
    .A2(_3012_),
    .B1(_3004_),
    .C1(_3688_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3689_));
 sky130_fd_sc_hd__a221o_1 _7444_ (.A1(net303),
    .A2(_3007_),
    .B1(_3009_),
    .B2(net318),
    .C1(_3689_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0587_));
 sky130_fd_sc_hd__and3_1 _7445_ (.A(\i_tinyqv.cpu.instr_data_start[16] ),
    .B(_0881_),
    .C(_3681_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3690_));
 sky130_fd_sc_hd__a21oi_1 _7446_ (.A1(_0881_),
    .A2(_3681_),
    .B1(\i_tinyqv.cpu.instr_data_start[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3691_));
 sky130_fd_sc_hd__or3_1 _7447_ (.A(\i_tinyqv.cpu.was_early_branch ),
    .B(_3690_),
    .C(_3691_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3692_));
 sky130_fd_sc_hd__o21ai_1 _7448_ (.A1(_1437_),
    .A2(_3169_),
    .B1(_3692_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3693_));
 sky130_fd_sc_hd__mux2_1 _7449_ (.A0(\i_tinyqv.cpu.data_addr[16] ),
    .A1(_3693_),
    .S(_2681_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3694_));
 sky130_fd_sc_hd__mux2_1 _7450_ (.A0(net147),
    .A1(_3694_),
    .S(_3004_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3695_));
 sky130_fd_sc_hd__mux2_1 _7451_ (.A0(\i_tinyqv.mem.q_ctrl.addr[16] ),
    .A1(_3695_),
    .S(_3625_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3696_));
 sky130_fd_sc_hd__clkbuf_1 _7452_ (.A(_3696_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0588_));
 sky130_fd_sc_hd__and2_1 _7453_ (.A(\i_tinyqv.cpu.instr_data_start[17] ),
    .B(_3690_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3697_));
 sky130_fd_sc_hd__nor2_1 _7454_ (.A(\i_tinyqv.cpu.instr_data_start[17] ),
    .B(_3690_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3698_));
 sky130_fd_sc_hd__o21a_1 _7455_ (.A1(_3697_),
    .A2(_3698_),
    .B1(_3239_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3699_));
 sky130_fd_sc_hd__a211oi_1 _7456_ (.A1(_3017_),
    .A2(_3180_),
    .B1(_3699_),
    .C1(_2877_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3700_));
 sky130_fd_sc_hd__a211o_1 _7457_ (.A1(net161),
    .A2(_2878_),
    .B1(_2732_),
    .C1(_3700_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3701_));
 sky130_fd_sc_hd__o221a_1 _7458_ (.A1(net304),
    .A2(_3624_),
    .B1(_3625_),
    .B2(net301),
    .C1(_3701_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0589_));
 sky130_fd_sc_hd__xnor2_1 _7459_ (.A(_0784_),
    .B(_3697_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3702_));
 sky130_fd_sc_hd__mux2_1 _7460_ (.A0(_3190_),
    .A1(_3702_),
    .S(_3239_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3703_));
 sky130_fd_sc_hd__nand2_1 _7461_ (.A(_3012_),
    .B(_3703_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3704_));
 sky130_fd_sc_hd__o21a_1 _7462_ (.A1(\i_tinyqv.cpu.data_addr[18] ),
    .A2(_2681_),
    .B1(_3004_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3705_));
 sky130_fd_sc_hd__a221o_1 _7463_ (.A1(\i_tinyqv.mem.q_ctrl.addr[14] ),
    .A2(_2732_),
    .B1(_3704_),
    .B2(_3705_),
    .C1(_3008_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3706_));
 sky130_fd_sc_hd__o21a_1 _7464_ (.A1(net189),
    .A2(_3625_),
    .B1(_3706_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0590_));
 sky130_fd_sc_hd__and3_1 _7465_ (.A(\i_tinyqv.cpu.instr_data_start[19] ),
    .B(_0784_),
    .C(_3697_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3707_));
 sky130_fd_sc_hd__a21oi_1 _7466_ (.A1(_0784_),
    .A2(_3697_),
    .B1(\i_tinyqv.cpu.instr_data_start[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3708_));
 sky130_fd_sc_hd__or3_1 _7467_ (.A(_3632_),
    .B(_3707_),
    .C(_3708_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3709_));
 sky130_fd_sc_hd__o211a_1 _7468_ (.A1(_3239_),
    .A2(_3199_),
    .B1(_3709_),
    .C1(_2682_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3710_));
 sky130_fd_sc_hd__o21ai_1 _7469_ (.A1(net288),
    .A2(_2682_),
    .B1(_3005_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3711_));
 sky130_fd_sc_hd__mux2_1 _7470_ (.A0(\i_tinyqv.mem.q_ctrl.addr[15] ),
    .A1(\i_tinyqv.mem.q_ctrl.addr[19] ),
    .S(_3624_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3712_));
 sky130_fd_sc_hd__a2bb2o_1 _7471_ (.A1_N(_3710_),
    .A2_N(_3711_),
    .B1(_2733_),
    .B2(_3712_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0591_));
 sky130_fd_sc_hd__mux2_1 _7472_ (.A0(\i_tinyqv.mem.q_ctrl.addr[20] ),
    .A1(\i_tinyqv.mem.q_ctrl.addr[16] ),
    .S(_3007_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3713_));
 sky130_fd_sc_hd__or2_1 _7473_ (.A(\i_tinyqv.cpu.instr_data_start[20] ),
    .B(_3707_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3714_));
 sky130_fd_sc_hd__and2_1 _7474_ (.A(\i_tinyqv.cpu.instr_data_start[20] ),
    .B(_3707_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3715_));
 sky130_fd_sc_hd__nor2_1 _7475_ (.A(_3017_),
    .B(_3715_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3716_));
 sky130_fd_sc_hd__a221o_1 _7476_ (.A1(_3017_),
    .A2(_3211_),
    .B1(_3714_),
    .B2(_3716_),
    .C1(_2878_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3717_));
 sky130_fd_sc_hd__o21a_1 _7477_ (.A1(\i_tinyqv.cpu.data_addr[20] ),
    .A2(_2682_),
    .B1(_3005_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3718_));
 sky130_fd_sc_hd__a22o_1 _7478_ (.A1(_2733_),
    .A2(_3713_),
    .B1(_3717_),
    .B2(_3718_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0592_));
 sky130_fd_sc_hd__or2_1 _7479_ (.A(\i_tinyqv.cpu.instr_data_start[21] ),
    .B(_3715_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3719_));
 sky130_fd_sc_hd__and3_1 _7480_ (.A(\i_tinyqv.cpu.instr_data_start[21] ),
    .B(\i_tinyqv.cpu.instr_data_start[20] ),
    .C(_3707_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3720_));
 sky130_fd_sc_hd__nor2_1 _7481_ (.A(_3010_),
    .B(_3720_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3721_));
 sky130_fd_sc_hd__a221o_1 _7482_ (.A1(_3632_),
    .A2(_3219_),
    .B1(_3719_),
    .B2(_3721_),
    .C1(_2877_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3722_));
 sky130_fd_sc_hd__o21a_1 _7483_ (.A1(\i_tinyqv.cpu.data_addr[21] ),
    .A2(_2682_),
    .B1(_3722_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3723_));
 sky130_fd_sc_hd__or2_1 _7484_ (.A(\i_tinyqv.mem.q_ctrl.addr[17] ),
    .B(_3624_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3724_));
 sky130_fd_sc_hd__o221a_1 _7485_ (.A1(\i_tinyqv.mem.q_ctrl.addr[21] ),
    .A2(_3625_),
    .B1(_3723_),
    .B2(_2733_),
    .C1(_3724_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0593_));
 sky130_fd_sc_hd__nor2_1 _7486_ (.A(_3239_),
    .B(_3228_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3725_));
 sky130_fd_sc_hd__nand2_1 _7487_ (.A(\i_tinyqv.cpu.instr_data_start[22] ),
    .B(_3720_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3726_));
 sky130_fd_sc_hd__or2_1 _7488_ (.A(\i_tinyqv.cpu.instr_data_start[22] ),
    .B(_3720_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3727_));
 sky130_fd_sc_hd__a21oi_1 _7489_ (.A1(_3726_),
    .A2(_3727_),
    .B1(_3017_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3728_));
 sky130_fd_sc_hd__a21oi_1 _7490_ (.A1(net177),
    .A2(_2878_),
    .B1(_2732_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3729_));
 sky130_fd_sc_hd__o31ai_1 _7491_ (.A1(_2878_),
    .A2(_3725_),
    .A3(_3728_),
    .B1(_3729_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3730_));
 sky130_fd_sc_hd__a21o_1 _7492_ (.A1(\i_tinyqv.mem.q_ctrl.addr[18] ),
    .A2(_3007_),
    .B1(_3005_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3731_));
 sky130_fd_sc_hd__a22o_1 _7493_ (.A1(\i_tinyqv.mem.q_ctrl.addr[22] ),
    .A2(_3009_),
    .B1(_3730_),
    .B2(_3731_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0594_));
 sky130_fd_sc_hd__nor2_1 _7494_ (.A(\i_tinyqv.cpu.instr_data_start[23] ),
    .B(_3726_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3732_));
 sky130_fd_sc_hd__a21o_1 _7495_ (.A1(\i_tinyqv.cpu.instr_data_start[23] ),
    .A2(_3726_),
    .B1(\i_tinyqv.cpu.was_early_branch ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3733_));
 sky130_fd_sc_hd__o22a_1 _7496_ (.A1(_3239_),
    .A2(_3234_),
    .B1(_3732_),
    .B2(_3733_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3734_));
 sky130_fd_sc_hd__mux2_1 _7497_ (.A0(\i_tinyqv.cpu.data_addr[23] ),
    .A1(_3734_),
    .S(_2681_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3735_));
 sky130_fd_sc_hd__mux2_1 _7498_ (.A0(\i_tinyqv.mem.q_ctrl.addr[23] ),
    .A1(\i_tinyqv.mem.q_ctrl.addr[19] ),
    .S(_3007_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3736_));
 sky130_fd_sc_hd__mux2_1 _7499_ (.A0(_3735_),
    .A1(_3736_),
    .S(_2732_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3737_));
 sky130_fd_sc_hd__clkbuf_1 _7500_ (.A(_3737_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0595_));
 sky130_fd_sc_hd__nor2_1 _7501_ (.A(_2066_),
    .B(_2071_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3738_));
 sky130_fd_sc_hd__o31a_1 _7502_ (.A1(net248),
    .A2(\i_tinyqv.cpu.i_core.cycle_count[0] ),
    .A3(_0744_),
    .B1(_3738_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0596_));
 sky130_fd_sc_hd__and2_1 _7503_ (.A(net121),
    .B(_2071_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3739_));
 sky130_fd_sc_hd__o21ai_1 _7504_ (.A1(net121),
    .A2(_2071_),
    .B1(_2049_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3740_));
 sky130_fd_sc_hd__nor2_1 _7505_ (.A(_3739_),
    .B(_3740_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0597_));
 sky130_fd_sc_hd__o21ai_1 _7506_ (.A1(\i_tinyqv.cpu.i_core.cycle_count[2] ),
    .A2(_3739_),
    .B1(_2049_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3741_));
 sky130_fd_sc_hd__nor2_1 _7507_ (.A(_2072_),
    .B(_3741_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0598_));
 sky130_fd_sc_hd__or2_1 _7508_ (.A(\i_tinyqv.cpu.i_core.cycle_count[3] ),
    .B(_2072_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3742_));
 sky130_fd_sc_hd__and3_1 _7509_ (.A(_2079_),
    .B(_2073_),
    .C(_3742_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3743_));
 sky130_fd_sc_hd__clkbuf_1 _7510_ (.A(_3743_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0599_));
 sky130_fd_sc_hd__mux2_1 _7511_ (.A0(\i_tinyqv.cpu.i_core.i_instrret.add ),
    .A1(\i_tinyqv.cpu.i_core.i_instrret.cy ),
    .S(_1026_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3744_));
 sky130_fd_sc_hd__and3_1 _7512_ (.A(net92),
    .B(\i_tinyqv.cpu.i_core.i_instrret.data[1] ),
    .C(_3744_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3745_));
 sky130_fd_sc_hd__and2_1 _7513_ (.A(\i_tinyqv.cpu.i_core.i_instrret.data[2] ),
    .B(_3745_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3746_));
 sky130_fd_sc_hd__and3_1 _7514_ (.A(_1752_),
    .B(net90),
    .C(_3746_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3747_));
 sky130_fd_sc_hd__clkbuf_1 _7515_ (.A(_3747_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0600_));
 sky130_fd_sc_hd__nor2_1 _7516_ (.A(_0939_),
    .B(_1755_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3748_));
 sky130_fd_sc_hd__mux2_1 _7517_ (.A0(\i_tinyqv.cpu.i_core.i_shift.b[4] ),
    .A1(_2644_),
    .S(_3748_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3749_));
 sky130_fd_sc_hd__clkbuf_1 _7518_ (.A(_3749_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0601_));
 sky130_fd_sc_hd__nor2_1 _7519_ (.A(_2067_),
    .B(_2073_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0602_));
 sky130_fd_sc_hd__and2_1 _7520_ (.A(net92),
    .B(_3744_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_3750_));
 sky130_fd_sc_hd__o21ai_1 _7521_ (.A1(net92),
    .A2(_3744_),
    .B1(_2049_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3751_));
 sky130_fd_sc_hd__nor2_1 _7522_ (.A(_3750_),
    .B(_3751_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0603_));
 sky130_fd_sc_hd__o21ai_1 _7523_ (.A1(net176),
    .A2(_3750_),
    .B1(_2049_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3752_));
 sky130_fd_sc_hd__nor2_1 _7524_ (.A(_3745_),
    .B(_3752_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0604_));
 sky130_fd_sc_hd__o21ai_1 _7525_ (.A1(net217),
    .A2(_3745_),
    .B1(_2049_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3753_));
 sky130_fd_sc_hd__nor2_1 _7526_ (.A(_3746_),
    .B(_3753_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0605_));
 sky130_fd_sc_hd__o21ai_1 _7527_ (.A1(net90),
    .A2(_3746_),
    .B1(_2079_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_3754_));
 sky130_fd_sc_hd__a21oi_1 _7528_ (.A1(net90),
    .A2(_3746_),
    .B1(_3754_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0606_));
 sky130_fd_sc_hd__dfxtp_1 _7529_ (.CLK(clknet_leaf_45_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.reg_buf[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[15][0] ));
 sky130_fd_sc_hd__dfxtp_1 _7530_ (.CLK(clknet_leaf_46_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.reg_buf[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[15][1] ));
 sky130_fd_sc_hd__dfxtp_1 _7531_ (.CLK(clknet_leaf_44_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.reg_buf[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[15][2] ));
 sky130_fd_sc_hd__dfxtp_1 _7532_ (.CLK(clknet_leaf_45_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.reg_buf[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[15][3] ));
 sky130_fd_sc_hd__dfxtp_1 _7533_ (.CLK(clknet_leaf_46_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.reg_buf[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[15][8] ));
 sky130_fd_sc_hd__dfxtp_1 _7534_ (.CLK(clknet_leaf_47_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.reg_buf[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[15][9] ));
 sky130_fd_sc_hd__dfxtp_1 _7535_ (.CLK(clknet_leaf_45_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.reg_buf[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[15][10] ));
 sky130_fd_sc_hd__dfxtp_1 _7536_ (.CLK(clknet_leaf_45_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.reg_buf[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[15][11] ));
 sky130_fd_sc_hd__dfxtp_1 _7537_ (.CLK(clknet_leaf_47_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.reg_buf[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[15][12] ));
 sky130_fd_sc_hd__dfxtp_1 _7538_ (.CLK(clknet_leaf_47_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.reg_buf[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[15][13] ));
 sky130_fd_sc_hd__dfxtp_1 _7539_ (.CLK(clknet_leaf_45_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.reg_buf[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[15][14] ));
 sky130_fd_sc_hd__dfxtp_1 _7540_ (.CLK(clknet_leaf_46_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.reg_buf[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[15][15] ));
 sky130_fd_sc_hd__dfxtp_1 _7541_ (.CLK(clknet_leaf_47_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.reg_buf[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[15][16] ));
 sky130_fd_sc_hd__dfxtp_1 _7542_ (.CLK(clknet_leaf_54_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.reg_buf[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[15][17] ));
 sky130_fd_sc_hd__dfxtp_1 _7543_ (.CLK(clknet_leaf_46_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.reg_buf[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[15][18] ));
 sky130_fd_sc_hd__dfxtp_1 _7544_ (.CLK(clknet_leaf_46_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.reg_buf[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[15][19] ));
 sky130_fd_sc_hd__dfxtp_1 _7545_ (.CLK(clknet_leaf_47_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.reg_buf[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[15][20] ));
 sky130_fd_sc_hd__dfxtp_1 _7546_ (.CLK(clknet_leaf_54_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.reg_buf[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[15][21] ));
 sky130_fd_sc_hd__dfxtp_1 _7547_ (.CLK(clknet_leaf_46_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.reg_buf[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[15][22] ));
 sky130_fd_sc_hd__dfxtp_1 _7548_ (.CLK(clknet_leaf_46_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.reg_buf[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[15][23] ));
 sky130_fd_sc_hd__dfxtp_1 _7549_ (.CLK(clknet_leaf_47_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.reg_buf[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[15][24] ));
 sky130_fd_sc_hd__dfxtp_1 _7550_ (.CLK(clknet_leaf_54_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.reg_buf[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[15][25] ));
 sky130_fd_sc_hd__dfxtp_1 _7551_ (.CLK(clknet_leaf_46_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.reg_buf[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[15][26] ));
 sky130_fd_sc_hd__dfxtp_1 _7552_ (.CLK(clknet_leaf_46_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.reg_buf[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[15][27] ));
 sky130_fd_sc_hd__dfxtp_1 _7553_ (.CLK(clknet_leaf_47_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.reg_buf[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[15][28] ));
 sky130_fd_sc_hd__dfxtp_1 _7554_ (.CLK(clknet_leaf_54_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.reg_buf[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[15][29] ));
 sky130_fd_sc_hd__dfxtp_1 _7555_ (.CLK(clknet_leaf_46_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.reg_buf[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[15][30] ));
 sky130_fd_sc_hd__dfxtp_1 _7556_ (.CLK(clknet_leaf_46_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.reg_buf[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[15][31] ));
 sky130_fd_sc_hd__dfxtp_1 _7557_ (.CLK(clknet_leaf_53_clk),
    .D(_0050_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[15][0] ));
 sky130_fd_sc_hd__dfxtp_1 _7558_ (.CLK(clknet_leaf_55_clk),
    .D(_0051_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[15][1] ));
 sky130_fd_sc_hd__dfxtp_1 _7559_ (.CLK(clknet_leaf_47_clk),
    .D(_0052_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[15][2] ));
 sky130_fd_sc_hd__dfxtp_1 _7560_ (.CLK(clknet_leaf_47_clk),
    .D(_0053_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[15][3] ));
 sky130_fd_sc_hd__dfxtp_1 _7561_ (.CLK(clknet_leaf_57_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.reg_buf[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[14][0] ));
 sky130_fd_sc_hd__dfxtp_1 _7562_ (.CLK(clknet_leaf_57_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.reg_buf[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[14][1] ));
 sky130_fd_sc_hd__dfxtp_1 _7563_ (.CLK(clknet_leaf_53_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.reg_buf[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[14][2] ));
 sky130_fd_sc_hd__dfxtp_1 _7564_ (.CLK(clknet_leaf_57_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.reg_buf[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[14][3] ));
 sky130_fd_sc_hd__dfxtp_1 _7565_ (.CLK(clknet_leaf_57_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.reg_buf[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[14][8] ));
 sky130_fd_sc_hd__dfxtp_1 _7566_ (.CLK(clknet_leaf_58_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.reg_buf[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[14][9] ));
 sky130_fd_sc_hd__dfxtp_1 _7567_ (.CLK(clknet_leaf_54_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.reg_buf[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[14][10] ));
 sky130_fd_sc_hd__dfxtp_1 _7568_ (.CLK(clknet_leaf_58_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.reg_buf[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[14][11] ));
 sky130_fd_sc_hd__dfxtp_1 _7569_ (.CLK(clknet_leaf_58_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.reg_buf[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[14][12] ));
 sky130_fd_sc_hd__dfxtp_1 _7570_ (.CLK(clknet_leaf_58_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.reg_buf[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[14][13] ));
 sky130_fd_sc_hd__dfxtp_1 _7571_ (.CLK(clknet_leaf_54_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.reg_buf[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[14][14] ));
 sky130_fd_sc_hd__dfxtp_1 _7572_ (.CLK(clknet_leaf_58_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.reg_buf[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[14][15] ));
 sky130_fd_sc_hd__dfxtp_1 _7573_ (.CLK(clknet_leaf_59_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.reg_buf[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[14][16] ));
 sky130_fd_sc_hd__dfxtp_1 _7574_ (.CLK(clknet_leaf_58_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.reg_buf[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[14][17] ));
 sky130_fd_sc_hd__dfxtp_1 _7575_ (.CLK(clknet_leaf_54_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.reg_buf[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[14][18] ));
 sky130_fd_sc_hd__dfxtp_1 _7576_ (.CLK(clknet_leaf_58_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.reg_buf[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[14][19] ));
 sky130_fd_sc_hd__dfxtp_1 _7577_ (.CLK(clknet_leaf_59_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.reg_buf[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[14][20] ));
 sky130_fd_sc_hd__dfxtp_1 _7578_ (.CLK(clknet_leaf_58_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.reg_buf[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[14][21] ));
 sky130_fd_sc_hd__dfxtp_1 _7579_ (.CLK(clknet_leaf_55_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.reg_buf[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[14][22] ));
 sky130_fd_sc_hd__dfxtp_1 _7580_ (.CLK(clknet_leaf_59_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.reg_buf[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[14][23] ));
 sky130_fd_sc_hd__dfxtp_1 _7581_ (.CLK(clknet_leaf_59_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.reg_buf[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[14][24] ));
 sky130_fd_sc_hd__dfxtp_1 _7582_ (.CLK(clknet_leaf_58_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.reg_buf[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[14][25] ));
 sky130_fd_sc_hd__dfxtp_1 _7583_ (.CLK(clknet_leaf_55_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.reg_buf[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[14][26] ));
 sky130_fd_sc_hd__dfxtp_1 _7584_ (.CLK(clknet_leaf_59_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.reg_buf[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[14][27] ));
 sky130_fd_sc_hd__dfxtp_1 _7585_ (.CLK(clknet_leaf_59_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.reg_buf[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[14][28] ));
 sky130_fd_sc_hd__dfxtp_1 _7586_ (.CLK(clknet_leaf_58_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.reg_buf[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[14][29] ));
 sky130_fd_sc_hd__dfxtp_1 _7587_ (.CLK(clknet_leaf_55_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.reg_buf[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[14][30] ));
 sky130_fd_sc_hd__dfxtp_1 _7588_ (.CLK(clknet_leaf_59_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.reg_buf[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[14][31] ));
 sky130_fd_sc_hd__dfxtp_1 _7589_ (.CLK(clknet_leaf_57_clk),
    .D(_0046_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[14][0] ));
 sky130_fd_sc_hd__dfxtp_1 _7590_ (.CLK(clknet_leaf_55_clk),
    .D(_0047_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[14][1] ));
 sky130_fd_sc_hd__dfxtp_1 _7591_ (.CLK(clknet_leaf_55_clk),
    .D(_0048_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[14][2] ));
 sky130_fd_sc_hd__dfxtp_1 _7592_ (.CLK(clknet_leaf_57_clk),
    .D(_0049_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[14][3] ));
 sky130_fd_sc_hd__dfxtp_1 _7593_ (.CLK(clknet_leaf_1_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.reg_buf[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[13][0] ));
 sky130_fd_sc_hd__dfxtp_1 _7594_ (.CLK(clknet_leaf_53_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.reg_buf[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[13][1] ));
 sky130_fd_sc_hd__dfxtp_1 _7595_ (.CLK(clknet_leaf_2_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.reg_buf[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[13][2] ));
 sky130_fd_sc_hd__dfxtp_1 _7596_ (.CLK(clknet_leaf_1_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.reg_buf[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[13][3] ));
 sky130_fd_sc_hd__dfxtp_1 _7597_ (.CLK(clknet_leaf_0_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.reg_buf[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[13][8] ));
 sky130_fd_sc_hd__dfxtp_1 _7598_ (.CLK(clknet_leaf_53_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.reg_buf[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[13][9] ));
 sky130_fd_sc_hd__dfxtp_1 _7599_ (.CLK(clknet_leaf_2_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.reg_buf[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[13][10] ));
 sky130_fd_sc_hd__dfxtp_1 _7600_ (.CLK(clknet_leaf_1_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.reg_buf[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[13][11] ));
 sky130_fd_sc_hd__dfxtp_1 _7601_ (.CLK(clknet_leaf_0_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.reg_buf[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[13][12] ));
 sky130_fd_sc_hd__dfxtp_1 _7602_ (.CLK(clknet_leaf_53_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.reg_buf[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[13][13] ));
 sky130_fd_sc_hd__dfxtp_1 _7603_ (.CLK(clknet_leaf_2_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.reg_buf[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[13][14] ));
 sky130_fd_sc_hd__dfxtp_1 _7604_ (.CLK(clknet_leaf_1_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.reg_buf[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[13][15] ));
 sky130_fd_sc_hd__dfxtp_1 _7605_ (.CLK(clknet_leaf_0_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.reg_buf[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[13][16] ));
 sky130_fd_sc_hd__dfxtp_1 _7606_ (.CLK(clknet_leaf_52_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.reg_buf[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[13][17] ));
 sky130_fd_sc_hd__dfxtp_1 _7607_ (.CLK(clknet_leaf_2_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.reg_buf[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[13][18] ));
 sky130_fd_sc_hd__dfxtp_1 _7608_ (.CLK(clknet_leaf_2_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.reg_buf[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[13][19] ));
 sky130_fd_sc_hd__dfxtp_1 _7609_ (.CLK(clknet_leaf_0_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.reg_buf[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[13][20] ));
 sky130_fd_sc_hd__dfxtp_1 _7610_ (.CLK(clknet_leaf_52_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.reg_buf[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[13][21] ));
 sky130_fd_sc_hd__dfxtp_1 _7611_ (.CLK(clknet_leaf_2_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.reg_buf[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[13][22] ));
 sky130_fd_sc_hd__dfxtp_1 _7612_ (.CLK(clknet_leaf_2_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.reg_buf[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[13][23] ));
 sky130_fd_sc_hd__dfxtp_1 _7613_ (.CLK(clknet_leaf_0_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.reg_buf[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[13][24] ));
 sky130_fd_sc_hd__dfxtp_1 _7614_ (.CLK(clknet_leaf_52_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.reg_buf[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[13][25] ));
 sky130_fd_sc_hd__dfxtp_1 _7615_ (.CLK(clknet_leaf_2_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.reg_buf[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[13][26] ));
 sky130_fd_sc_hd__dfxtp_1 _7616_ (.CLK(clknet_leaf_2_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.reg_buf[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[13][27] ));
 sky130_fd_sc_hd__dfxtp_1 _7617_ (.CLK(clknet_leaf_0_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.reg_buf[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[13][28] ));
 sky130_fd_sc_hd__dfxtp_1 _7618_ (.CLK(clknet_leaf_52_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.reg_buf[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[13][29] ));
 sky130_fd_sc_hd__dfxtp_1 _7619_ (.CLK(clknet_leaf_2_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.reg_buf[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[13][30] ));
 sky130_fd_sc_hd__dfxtp_1 _7620_ (.CLK(clknet_leaf_2_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.reg_buf[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[13][31] ));
 sky130_fd_sc_hd__dfxtp_1 _7621_ (.CLK(clknet_leaf_1_clk),
    .D(_0042_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[13][0] ));
 sky130_fd_sc_hd__dfxtp_1 _7622_ (.CLK(clknet_leaf_56_clk),
    .D(_0043_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[13][1] ));
 sky130_fd_sc_hd__dfxtp_1 _7623_ (.CLK(clknet_leaf_1_clk),
    .D(_0044_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[13][2] ));
 sky130_fd_sc_hd__dfxtp_1 _7624_ (.CLK(clknet_leaf_1_clk),
    .D(_0045_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[13][3] ));
 sky130_fd_sc_hd__dfxtp_1 _7625_ (.CLK(clknet_leaf_52_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.reg_buf[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[12][0] ));
 sky130_fd_sc_hd__dfxtp_1 _7626_ (.CLK(clknet_leaf_55_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.reg_buf[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[12][1] ));
 sky130_fd_sc_hd__dfxtp_1 _7627_ (.CLK(clknet_leaf_44_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.reg_buf[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[12][2] ));
 sky130_fd_sc_hd__dfxtp_1 _7628_ (.CLK(clknet_leaf_44_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.reg_buf[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[12][3] ));
 sky130_fd_sc_hd__dfxtp_1 _7629_ (.CLK(clknet_leaf_56_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.reg_buf[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[12][8] ));
 sky130_fd_sc_hd__dfxtp_1 _7630_ (.CLK(clknet_leaf_55_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.reg_buf[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[12][9] ));
 sky130_fd_sc_hd__dfxtp_1 _7631_ (.CLK(clknet_leaf_45_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.reg_buf[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[12][10] ));
 sky130_fd_sc_hd__dfxtp_1 _7632_ (.CLK(clknet_leaf_44_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.reg_buf[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[12][11] ));
 sky130_fd_sc_hd__dfxtp_1 _7633_ (.CLK(clknet_leaf_56_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.reg_buf[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[12][12] ));
 sky130_fd_sc_hd__dfxtp_1 _7634_ (.CLK(clknet_leaf_55_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.reg_buf[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[12][13] ));
 sky130_fd_sc_hd__dfxtp_1 _7635_ (.CLK(clknet_leaf_45_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.reg_buf[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[12][14] ));
 sky130_fd_sc_hd__dfxtp_1 _7636_ (.CLK(clknet_leaf_45_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.reg_buf[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[12][15] ));
 sky130_fd_sc_hd__dfxtp_1 _7637_ (.CLK(clknet_leaf_56_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.reg_buf[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[12][16] ));
 sky130_fd_sc_hd__dfxtp_1 _7638_ (.CLK(clknet_leaf_55_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.reg_buf[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[12][17] ));
 sky130_fd_sc_hd__dfxtp_1 _7639_ (.CLK(clknet_leaf_46_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.reg_buf[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[12][18] ));
 sky130_fd_sc_hd__dfxtp_1 _7640_ (.CLK(clknet_leaf_46_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.reg_buf[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[12][19] ));
 sky130_fd_sc_hd__dfxtp_1 _7641_ (.CLK(clknet_leaf_56_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.reg_buf[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[12][20] ));
 sky130_fd_sc_hd__dfxtp_1 _7642_ (.CLK(clknet_leaf_55_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.reg_buf[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[12][21] ));
 sky130_fd_sc_hd__dfxtp_1 _7643_ (.CLK(clknet_leaf_46_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.reg_buf[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[12][22] ));
 sky130_fd_sc_hd__dfxtp_1 _7644_ (.CLK(clknet_leaf_46_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.reg_buf[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[12][23] ));
 sky130_fd_sc_hd__dfxtp_1 _7645_ (.CLK(clknet_leaf_57_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.reg_buf[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[12][24] ));
 sky130_fd_sc_hd__dfxtp_1 _7646_ (.CLK(clknet_leaf_57_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.reg_buf[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[12][25] ));
 sky130_fd_sc_hd__dfxtp_1 _7647_ (.CLK(clknet_leaf_46_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.reg_buf[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[12][26] ));
 sky130_fd_sc_hd__dfxtp_1 _7648_ (.CLK(clknet_leaf_46_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.reg_buf[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[12][27] ));
 sky130_fd_sc_hd__dfxtp_1 _7649_ (.CLK(clknet_leaf_57_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.reg_buf[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[12][28] ));
 sky130_fd_sc_hd__dfxtp_1 _7650_ (.CLK(clknet_leaf_58_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.reg_buf[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[12][29] ));
 sky130_fd_sc_hd__dfxtp_1 _7651_ (.CLK(clknet_leaf_47_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.reg_buf[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[12][30] ));
 sky130_fd_sc_hd__dfxtp_1 _7652_ (.CLK(clknet_leaf_46_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.reg_buf[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[12][31] ));
 sky130_fd_sc_hd__dfxtp_1 _7653_ (.CLK(clknet_leaf_56_clk),
    .D(_0038_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[12][0] ));
 sky130_fd_sc_hd__dfxtp_1 _7654_ (.CLK(clknet_leaf_55_clk),
    .D(_0039_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[12][1] ));
 sky130_fd_sc_hd__dfxtp_1 _7655_ (.CLK(clknet_leaf_47_clk),
    .D(_0040_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[12][2] ));
 sky130_fd_sc_hd__dfxtp_1 _7656_ (.CLK(clknet_leaf_47_clk),
    .D(_0041_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[12][3] ));
 sky130_fd_sc_hd__dfxtp_1 _7657_ (.CLK(clknet_leaf_1_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.reg_buf[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[11][0] ));
 sky130_fd_sc_hd__dfxtp_1 _7658_ (.CLK(clknet_leaf_55_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.reg_buf[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[11][1] ));
 sky130_fd_sc_hd__dfxtp_1 _7659_ (.CLK(clknet_leaf_58_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.reg_buf[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[11][2] ));
 sky130_fd_sc_hd__dfxtp_1 _7660_ (.CLK(clknet_leaf_45_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.reg_buf[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[11][3] ));
 sky130_fd_sc_hd__dfxtp_1 _7661_ (.CLK(clknet_leaf_0_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.reg_buf[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[11][8] ));
 sky130_fd_sc_hd__dfxtp_1 _7662_ (.CLK(clknet_leaf_55_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.reg_buf[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[11][9] ));
 sky130_fd_sc_hd__dfxtp_1 _7663_ (.CLK(clknet_leaf_58_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.reg_buf[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[11][10] ));
 sky130_fd_sc_hd__dfxtp_1 _7664_ (.CLK(clknet_leaf_45_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.reg_buf[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[11][11] ));
 sky130_fd_sc_hd__dfxtp_1 _7665_ (.CLK(clknet_leaf_0_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.reg_buf[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[11][12] ));
 sky130_fd_sc_hd__dfxtp_1 _7666_ (.CLK(clknet_leaf_56_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.reg_buf[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[11][13] ));
 sky130_fd_sc_hd__dfxtp_1 _7667_ (.CLK(clknet_leaf_58_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.reg_buf[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[11][14] ));
 sky130_fd_sc_hd__dfxtp_1 _7668_ (.CLK(clknet_leaf_46_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.reg_buf[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[11][15] ));
 sky130_fd_sc_hd__dfxtp_1 _7669_ (.CLK(clknet_leaf_59_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.reg_buf[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[11][16] ));
 sky130_fd_sc_hd__dfxtp_1 _7670_ (.CLK(clknet_leaf_55_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.reg_buf[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[11][17] ));
 sky130_fd_sc_hd__dfxtp_1 _7671_ (.CLK(clknet_leaf_58_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.reg_buf[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[11][18] ));
 sky130_fd_sc_hd__dfxtp_1 _7672_ (.CLK(clknet_leaf_46_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.reg_buf[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[11][19] ));
 sky130_fd_sc_hd__dfxtp_1 _7673_ (.CLK(clknet_leaf_59_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.reg_buf[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[11][20] ));
 sky130_fd_sc_hd__dfxtp_1 _7674_ (.CLK(clknet_leaf_55_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.reg_buf[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[11][21] ));
 sky130_fd_sc_hd__dfxtp_1 _7675_ (.CLK(clknet_leaf_58_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.reg_buf[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[11][22] ));
 sky130_fd_sc_hd__dfxtp_1 _7676_ (.CLK(clknet_leaf_46_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.reg_buf[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[11][23] ));
 sky130_fd_sc_hd__dfxtp_1 _7677_ (.CLK(clknet_leaf_59_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.reg_buf[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[11][24] ));
 sky130_fd_sc_hd__dfxtp_1 _7678_ (.CLK(clknet_leaf_55_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.reg_buf[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[11][25] ));
 sky130_fd_sc_hd__dfxtp_1 _7679_ (.CLK(clknet_leaf_58_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.reg_buf[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[11][26] ));
 sky130_fd_sc_hd__dfxtp_1 _7680_ (.CLK(clknet_leaf_46_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.reg_buf[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[11][27] ));
 sky130_fd_sc_hd__dfxtp_1 _7681_ (.CLK(clknet_leaf_59_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.reg_buf[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[11][28] ));
 sky130_fd_sc_hd__dfxtp_1 _7682_ (.CLK(clknet_leaf_57_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.reg_buf[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[11][29] ));
 sky130_fd_sc_hd__dfxtp_1 _7683_ (.CLK(clknet_leaf_58_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.reg_buf[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[11][30] ));
 sky130_fd_sc_hd__dfxtp_1 _7684_ (.CLK(clknet_leaf_47_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.reg_buf[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[11][31] ));
 sky130_fd_sc_hd__dfxtp_1 _7685_ (.CLK(clknet_leaf_57_clk),
    .D(_0034_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[11][0] ));
 sky130_fd_sc_hd__dfxtp_1 _7686_ (.CLK(clknet_leaf_56_clk),
    .D(_0035_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[11][1] ));
 sky130_fd_sc_hd__dfxtp_1 _7687_ (.CLK(clknet_leaf_57_clk),
    .D(_0036_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[11][2] ));
 sky130_fd_sc_hd__dfxtp_1 _7688_ (.CLK(clknet_leaf_54_clk),
    .D(_0037_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[11][3] ));
 sky130_fd_sc_hd__dfxtp_1 _7689_ (.CLK(clknet_leaf_1_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.reg_buf[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[10][0] ));
 sky130_fd_sc_hd__dfxtp_1 _7690_ (.CLK(clknet_leaf_53_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.reg_buf[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[10][1] ));
 sky130_fd_sc_hd__dfxtp_1 _7691_ (.CLK(clknet_leaf_53_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.reg_buf[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[10][2] ));
 sky130_fd_sc_hd__dfxtp_1 _7692_ (.CLK(clknet_leaf_57_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.reg_buf[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[10][3] ));
 sky130_fd_sc_hd__dfxtp_1 _7693_ (.CLK(clknet_leaf_2_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.reg_buf[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[10][8] ));
 sky130_fd_sc_hd__dfxtp_1 _7694_ (.CLK(clknet_leaf_53_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.reg_buf[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[10][9] ));
 sky130_fd_sc_hd__dfxtp_1 _7695_ (.CLK(clknet_leaf_53_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.reg_buf[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[10][10] ));
 sky130_fd_sc_hd__dfxtp_1 _7696_ (.CLK(clknet_leaf_57_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.reg_buf[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[10][11] ));
 sky130_fd_sc_hd__dfxtp_1 _7697_ (.CLK(clknet_leaf_2_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.reg_buf[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[10][12] ));
 sky130_fd_sc_hd__dfxtp_1 _7698_ (.CLK(clknet_leaf_56_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.reg_buf[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[10][13] ));
 sky130_fd_sc_hd__dfxtp_1 _7699_ (.CLK(clknet_leaf_53_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.reg_buf[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[10][14] ));
 sky130_fd_sc_hd__dfxtp_1 _7700_ (.CLK(clknet_leaf_58_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.reg_buf[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[10][15] ));
 sky130_fd_sc_hd__dfxtp_1 _7701_ (.CLK(clknet_leaf_2_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.reg_buf[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[10][16] ));
 sky130_fd_sc_hd__dfxtp_1 _7702_ (.CLK(clknet_leaf_56_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.reg_buf[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[10][17] ));
 sky130_fd_sc_hd__dfxtp_1 _7703_ (.CLK(clknet_leaf_53_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.reg_buf[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[10][18] ));
 sky130_fd_sc_hd__dfxtp_1 _7704_ (.CLK(clknet_leaf_58_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.reg_buf[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[10][19] ));
 sky130_fd_sc_hd__dfxtp_1 _7705_ (.CLK(clknet_leaf_0_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.reg_buf[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[10][20] ));
 sky130_fd_sc_hd__dfxtp_1 _7706_ (.CLK(clknet_leaf_56_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.reg_buf[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[10][21] ));
 sky130_fd_sc_hd__dfxtp_1 _7707_ (.CLK(clknet_leaf_52_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.reg_buf[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[10][22] ));
 sky130_fd_sc_hd__dfxtp_1 _7708_ (.CLK(clknet_leaf_59_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.reg_buf[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[10][23] ));
 sky130_fd_sc_hd__dfxtp_1 _7709_ (.CLK(clknet_leaf_2_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.reg_buf[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[10][24] ));
 sky130_fd_sc_hd__dfxtp_1 _7710_ (.CLK(clknet_leaf_56_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.reg_buf[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[10][25] ));
 sky130_fd_sc_hd__dfxtp_1 _7711_ (.CLK(clknet_leaf_52_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.reg_buf[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[10][26] ));
 sky130_fd_sc_hd__dfxtp_1 _7712_ (.CLK(clknet_leaf_59_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.reg_buf[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[10][27] ));
 sky130_fd_sc_hd__dfxtp_1 _7713_ (.CLK(clknet_leaf_0_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.reg_buf[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[10][28] ));
 sky130_fd_sc_hd__dfxtp_1 _7714_ (.CLK(clknet_leaf_56_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.reg_buf[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[10][29] ));
 sky130_fd_sc_hd__dfxtp_1 _7715_ (.CLK(clknet_leaf_56_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.reg_buf[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[10][30] ));
 sky130_fd_sc_hd__dfxtp_1 _7716_ (.CLK(clknet_leaf_59_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.reg_buf[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[10][31] ));
 sky130_fd_sc_hd__dfxtp_1 _7717_ (.CLK(clknet_leaf_1_clk),
    .D(_0030_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[10][0] ));
 sky130_fd_sc_hd__dfxtp_1 _7718_ (.CLK(clknet_leaf_56_clk),
    .D(_0031_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[10][1] ));
 sky130_fd_sc_hd__dfxtp_1 _7719_ (.CLK(clknet_leaf_56_clk),
    .D(_0032_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[10][2] ));
 sky130_fd_sc_hd__dfxtp_1 _7720_ (.CLK(clknet_leaf_57_clk),
    .D(_0033_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[10][3] ));
 sky130_fd_sc_hd__dfxtp_1 _7721_ (.CLK(clknet_leaf_1_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.reg_buf[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[9][0] ));
 sky130_fd_sc_hd__dfxtp_1 _7722_ (.CLK(clknet_leaf_54_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.reg_buf[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[9][1] ));
 sky130_fd_sc_hd__dfxtp_1 _7723_ (.CLK(clknet_leaf_1_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.reg_buf[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[9][2] ));
 sky130_fd_sc_hd__dfxtp_1 _7724_ (.CLK(clknet_leaf_53_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.reg_buf[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[9][3] ));
 sky130_fd_sc_hd__dfxtp_1 _7725_ (.CLK(clknet_leaf_0_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.reg_buf[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[9][8] ));
 sky130_fd_sc_hd__dfxtp_1 _7726_ (.CLK(clknet_leaf_54_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.reg_buf[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[9][9] ));
 sky130_fd_sc_hd__dfxtp_1 _7727_ (.CLK(clknet_leaf_0_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.reg_buf[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[9][10] ));
 sky130_fd_sc_hd__dfxtp_1 _7728_ (.CLK(clknet_leaf_53_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.reg_buf[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[9][11] ));
 sky130_fd_sc_hd__dfxtp_1 _7729_ (.CLK(clknet_leaf_59_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.reg_buf[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[9][12] ));
 sky130_fd_sc_hd__dfxtp_1 _7730_ (.CLK(clknet_leaf_54_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.reg_buf[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[9][13] ));
 sky130_fd_sc_hd__dfxtp_1 _7731_ (.CLK(clknet_leaf_0_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.reg_buf[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[9][14] ));
 sky130_fd_sc_hd__dfxtp_1 _7732_ (.CLK(clknet_leaf_53_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.reg_buf[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[9][15] ));
 sky130_fd_sc_hd__dfxtp_1 _7733_ (.CLK(clknet_leaf_59_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.reg_buf[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[9][16] ));
 sky130_fd_sc_hd__dfxtp_1 _7734_ (.CLK(clknet_leaf_55_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.reg_buf[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[9][17] ));
 sky130_fd_sc_hd__dfxtp_1 _7735_ (.CLK(clknet_leaf_59_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.reg_buf[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[9][18] ));
 sky130_fd_sc_hd__dfxtp_1 _7736_ (.CLK(clknet_leaf_53_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.reg_buf[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[9][19] ));
 sky130_fd_sc_hd__dfxtp_1 _7737_ (.CLK(clknet_leaf_59_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.reg_buf[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[9][20] ));
 sky130_fd_sc_hd__dfxtp_1 _7738_ (.CLK(clknet_leaf_55_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.reg_buf[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[9][21] ));
 sky130_fd_sc_hd__dfxtp_1 _7739_ (.CLK(clknet_leaf_0_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.reg_buf[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[9][22] ));
 sky130_fd_sc_hd__dfxtp_1 _7740_ (.CLK(clknet_leaf_53_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.reg_buf[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[9][23] ));
 sky130_fd_sc_hd__dfxtp_1 _7741_ (.CLK(clknet_leaf_59_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.reg_buf[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[9][24] ));
 sky130_fd_sc_hd__dfxtp_1 _7742_ (.CLK(clknet_leaf_55_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.reg_buf[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[9][25] ));
 sky130_fd_sc_hd__dfxtp_1 _7743_ (.CLK(clknet_leaf_0_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.reg_buf[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[9][26] ));
 sky130_fd_sc_hd__dfxtp_1 _7744_ (.CLK(clknet_leaf_54_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.reg_buf[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[9][27] ));
 sky130_fd_sc_hd__dfxtp_1 _7745_ (.CLK(clknet_leaf_0_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.reg_buf[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[9][28] ));
 sky130_fd_sc_hd__dfxtp_1 _7746_ (.CLK(clknet_leaf_55_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.reg_buf[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[9][29] ));
 sky130_fd_sc_hd__dfxtp_1 _7747_ (.CLK(clknet_leaf_0_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.reg_buf[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[9][30] ));
 sky130_fd_sc_hd__dfxtp_1 _7748_ (.CLK(clknet_leaf_55_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.reg_buf[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[9][31] ));
 sky130_fd_sc_hd__dfxtp_1 _7749_ (.CLK(clknet_leaf_57_clk),
    .D(_0078_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[9][0] ));
 sky130_fd_sc_hd__dfxtp_1 _7750_ (.CLK(clknet_leaf_55_clk),
    .D(_0079_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[9][1] ));
 sky130_fd_sc_hd__dfxtp_1 _7751_ (.CLK(clknet_leaf_1_clk),
    .D(_0080_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[9][2] ));
 sky130_fd_sc_hd__dfxtp_1 _7752_ (.CLK(clknet_leaf_56_clk),
    .D(_0081_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[9][3] ));
 sky130_fd_sc_hd__dfxtp_1 _7753_ (.CLK(clknet_leaf_57_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.reg_buf[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[8][0] ));
 sky130_fd_sc_hd__dfxtp_1 _7754_ (.CLK(clknet_leaf_46_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.reg_buf[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[8][1] ));
 sky130_fd_sc_hd__dfxtp_1 _7755_ (.CLK(clknet_leaf_47_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.reg_buf[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[8][2] ));
 sky130_fd_sc_hd__dfxtp_1 _7756_ (.CLK(clknet_leaf_55_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.reg_buf[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[8][3] ));
 sky130_fd_sc_hd__dfxtp_1 _7757_ (.CLK(clknet_leaf_1_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.reg_buf[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[8][8] ));
 sky130_fd_sc_hd__dfxtp_1 _7758_ (.CLK(clknet_leaf_47_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.reg_buf[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[8][9] ));
 sky130_fd_sc_hd__dfxtp_1 _7759_ (.CLK(clknet_leaf_53_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.reg_buf[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[8][10] ));
 sky130_fd_sc_hd__dfxtp_1 _7760_ (.CLK(clknet_leaf_57_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.reg_buf[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[8][11] ));
 sky130_fd_sc_hd__dfxtp_1 _7761_ (.CLK(clknet_leaf_1_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.reg_buf[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[8][12] ));
 sky130_fd_sc_hd__dfxtp_1 _7762_ (.CLK(clknet_leaf_54_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.reg_buf[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[8][13] ));
 sky130_fd_sc_hd__dfxtp_1 _7763_ (.CLK(clknet_leaf_53_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.reg_buf[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[8][14] ));
 sky130_fd_sc_hd__dfxtp_1 _7764_ (.CLK(clknet_leaf_58_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.reg_buf[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[8][15] ));
 sky130_fd_sc_hd__dfxtp_1 _7765_ (.CLK(clknet_leaf_1_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.reg_buf[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[8][16] ));
 sky130_fd_sc_hd__dfxtp_1 _7766_ (.CLK(clknet_leaf_54_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.reg_buf[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[8][17] ));
 sky130_fd_sc_hd__dfxtp_1 _7767_ (.CLK(clknet_leaf_54_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.reg_buf[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[8][18] ));
 sky130_fd_sc_hd__dfxtp_1 _7768_ (.CLK(clknet_leaf_58_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.reg_buf[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[8][19] ));
 sky130_fd_sc_hd__dfxtp_1 _7769_ (.CLK(clknet_leaf_0_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.reg_buf[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[8][20] ));
 sky130_fd_sc_hd__dfxtp_1 _7770_ (.CLK(clknet_leaf_54_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.reg_buf[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[8][21] ));
 sky130_fd_sc_hd__dfxtp_1 _7771_ (.CLK(clknet_leaf_53_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.reg_buf[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[8][22] ));
 sky130_fd_sc_hd__dfxtp_1 _7772_ (.CLK(clknet_leaf_58_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.reg_buf[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[8][23] ));
 sky130_fd_sc_hd__dfxtp_1 _7773_ (.CLK(clknet_leaf_0_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.reg_buf[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[8][24] ));
 sky130_fd_sc_hd__dfxtp_1 _7774_ (.CLK(clknet_leaf_54_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.reg_buf[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[8][25] ));
 sky130_fd_sc_hd__dfxtp_1 _7775_ (.CLK(clknet_leaf_53_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.reg_buf[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[8][26] ));
 sky130_fd_sc_hd__dfxtp_1 _7776_ (.CLK(clknet_leaf_58_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.reg_buf[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[8][27] ));
 sky130_fd_sc_hd__dfxtp_1 _7777_ (.CLK(clknet_leaf_0_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.reg_buf[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[8][28] ));
 sky130_fd_sc_hd__dfxtp_1 _7778_ (.CLK(clknet_leaf_54_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.reg_buf[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[8][29] ));
 sky130_fd_sc_hd__dfxtp_1 _7779_ (.CLK(clknet_leaf_54_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.reg_buf[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[8][30] ));
 sky130_fd_sc_hd__dfxtp_1 _7780_ (.CLK(clknet_leaf_58_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.reg_buf[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[8][31] ));
 sky130_fd_sc_hd__dfxtp_1 _7781_ (.CLK(clknet_leaf_56_clk),
    .D(_0074_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[8][0] ));
 sky130_fd_sc_hd__dfxtp_1 _7782_ (.CLK(clknet_leaf_55_clk),
    .D(_0075_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[8][1] ));
 sky130_fd_sc_hd__dfxtp_1 _7783_ (.CLK(clknet_leaf_54_clk),
    .D(_0076_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[8][2] ));
 sky130_fd_sc_hd__dfxtp_1 _7784_ (.CLK(clknet_leaf_57_clk),
    .D(_0077_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[8][3] ));
 sky130_fd_sc_hd__dfxtp_1 _7785_ (.CLK(clknet_leaf_1_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.reg_buf[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[7][0] ));
 sky130_fd_sc_hd__dfxtp_1 _7786_ (.CLK(clknet_leaf_52_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.reg_buf[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[7][1] ));
 sky130_fd_sc_hd__dfxtp_1 _7787_ (.CLK(clknet_leaf_52_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.reg_buf[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[7][2] ));
 sky130_fd_sc_hd__dfxtp_1 _7788_ (.CLK(clknet_leaf_1_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.reg_buf[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[7][3] ));
 sky130_fd_sc_hd__dfxtp_1 _7789_ (.CLK(clknet_leaf_2_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.reg_buf[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[7][8] ));
 sky130_fd_sc_hd__dfxtp_1 _7790_ (.CLK(clknet_leaf_56_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.reg_buf[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[7][9] ));
 sky130_fd_sc_hd__dfxtp_1 _7791_ (.CLK(clknet_leaf_56_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.reg_buf[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[7][10] ));
 sky130_fd_sc_hd__dfxtp_1 _7792_ (.CLK(clknet_leaf_1_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.reg_buf[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[7][11] ));
 sky130_fd_sc_hd__dfxtp_1 _7793_ (.CLK(clknet_leaf_2_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.reg_buf[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[7][12] ));
 sky130_fd_sc_hd__dfxtp_1 _7794_ (.CLK(clknet_leaf_57_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.reg_buf[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[7][13] ));
 sky130_fd_sc_hd__dfxtp_1 _7795_ (.CLK(clknet_leaf_56_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.reg_buf[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[7][14] ));
 sky130_fd_sc_hd__dfxtp_1 _7796_ (.CLK(clknet_leaf_0_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.reg_buf[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[7][15] ));
 sky130_fd_sc_hd__dfxtp_1 _7797_ (.CLK(clknet_leaf_3_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.reg_buf[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[7][16] ));
 sky130_fd_sc_hd__dfxtp_1 _7798_ (.CLK(clknet_leaf_1_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.reg_buf[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[7][17] ));
 sky130_fd_sc_hd__dfxtp_1 _7799_ (.CLK(clknet_leaf_57_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.reg_buf[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[7][18] ));
 sky130_fd_sc_hd__dfxtp_1 _7800_ (.CLK(clknet_leaf_0_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.reg_buf[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[7][19] ));
 sky130_fd_sc_hd__dfxtp_1 _7801_ (.CLK(clknet_leaf_3_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.reg_buf[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[7][20] ));
 sky130_fd_sc_hd__dfxtp_1 _7802_ (.CLK(clknet_leaf_1_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.reg_buf[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[7][21] ));
 sky130_fd_sc_hd__dfxtp_1 _7803_ (.CLK(clknet_leaf_57_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.reg_buf[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[7][22] ));
 sky130_fd_sc_hd__dfxtp_1 _7804_ (.CLK(clknet_leaf_0_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.reg_buf[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[7][23] ));
 sky130_fd_sc_hd__dfxtp_1 _7805_ (.CLK(clknet_leaf_2_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.reg_buf[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[7][24] ));
 sky130_fd_sc_hd__dfxtp_1 _7806_ (.CLK(clknet_leaf_1_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.reg_buf[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[7][25] ));
 sky130_fd_sc_hd__dfxtp_1 _7807_ (.CLK(clknet_leaf_57_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.reg_buf[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[7][26] ));
 sky130_fd_sc_hd__dfxtp_1 _7808_ (.CLK(clknet_leaf_0_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.reg_buf[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[7][27] ));
 sky130_fd_sc_hd__dfxtp_1 _7809_ (.CLK(clknet_leaf_2_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.reg_buf[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[7][28] ));
 sky130_fd_sc_hd__dfxtp_1 _7810_ (.CLK(clknet_leaf_57_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.reg_buf[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[7][29] ));
 sky130_fd_sc_hd__dfxtp_1 _7811_ (.CLK(clknet_leaf_56_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.reg_buf[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[7][30] ));
 sky130_fd_sc_hd__dfxtp_1 _7812_ (.CLK(clknet_leaf_0_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.reg_buf[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[7][31] ));
 sky130_fd_sc_hd__dfxtp_1 _7813_ (.CLK(clknet_leaf_5_clk),
    .D(_0070_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[7][0] ));
 sky130_fd_sc_hd__dfxtp_1 _7814_ (.CLK(clknet_leaf_56_clk),
    .D(_0071_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[7][1] ));
 sky130_fd_sc_hd__dfxtp_1 _7815_ (.CLK(clknet_leaf_57_clk),
    .D(_0072_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[7][2] ));
 sky130_fd_sc_hd__dfxtp_1 _7816_ (.CLK(clknet_leaf_1_clk),
    .D(_0073_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[7][3] ));
 sky130_fd_sc_hd__dfxtp_1 _7817_ (.CLK(clknet_leaf_49_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.reg_buf[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[6][0] ));
 sky130_fd_sc_hd__dfxtp_1 _7818_ (.CLK(clknet_leaf_5_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.reg_buf[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[6][1] ));
 sky130_fd_sc_hd__dfxtp_1 _7819_ (.CLK(clknet_leaf_5_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.reg_buf[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[6][2] ));
 sky130_fd_sc_hd__dfxtp_1 _7820_ (.CLK(clknet_leaf_52_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.reg_buf[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[6][3] ));
 sky130_fd_sc_hd__dfxtp_1 _7821_ (.CLK(clknet_leaf_49_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.reg_buf[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[6][8] ));
 sky130_fd_sc_hd__dfxtp_1 _7822_ (.CLK(clknet_leaf_5_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.reg_buf[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[6][9] ));
 sky130_fd_sc_hd__dfxtp_1 _7823_ (.CLK(clknet_leaf_5_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.reg_buf[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[6][10] ));
 sky130_fd_sc_hd__dfxtp_1 _7824_ (.CLK(clknet_leaf_52_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.reg_buf[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[6][11] ));
 sky130_fd_sc_hd__dfxtp_1 _7825_ (.CLK(clknet_leaf_49_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.reg_buf[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[6][12] ));
 sky130_fd_sc_hd__dfxtp_1 _7826_ (.CLK(clknet_leaf_4_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.reg_buf[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[6][13] ));
 sky130_fd_sc_hd__dfxtp_1 _7827_ (.CLK(clknet_leaf_4_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.reg_buf[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[6][14] ));
 sky130_fd_sc_hd__dfxtp_1 _7828_ (.CLK(clknet_leaf_52_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.reg_buf[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[6][15] ));
 sky130_fd_sc_hd__dfxtp_1 _7829_ (.CLK(clknet_leaf_49_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.reg_buf[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[6][16] ));
 sky130_fd_sc_hd__dfxtp_1 _7830_ (.CLK(clknet_leaf_3_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.reg_buf[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[6][17] ));
 sky130_fd_sc_hd__dfxtp_1 _7831_ (.CLK(clknet_leaf_3_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.reg_buf[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[6][18] ));
 sky130_fd_sc_hd__dfxtp_1 _7832_ (.CLK(clknet_leaf_52_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.reg_buf[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[6][19] ));
 sky130_fd_sc_hd__dfxtp_1 _7833_ (.CLK(clknet_leaf_48_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.reg_buf[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[6][20] ));
 sky130_fd_sc_hd__dfxtp_1 _7834_ (.CLK(clknet_leaf_3_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.reg_buf[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[6][21] ));
 sky130_fd_sc_hd__dfxtp_1 _7835_ (.CLK(clknet_leaf_3_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.reg_buf[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[6][22] ));
 sky130_fd_sc_hd__dfxtp_1 _7836_ (.CLK(clknet_leaf_1_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.reg_buf[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[6][23] ));
 sky130_fd_sc_hd__dfxtp_1 _7837_ (.CLK(clknet_leaf_48_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.reg_buf[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[6][24] ));
 sky130_fd_sc_hd__dfxtp_1 _7838_ (.CLK(clknet_leaf_3_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.reg_buf[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[6][25] ));
 sky130_fd_sc_hd__dfxtp_1 _7839_ (.CLK(clknet_leaf_3_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.reg_buf[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[6][26] ));
 sky130_fd_sc_hd__dfxtp_1 _7840_ (.CLK(clknet_leaf_5_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.reg_buf[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[6][27] ));
 sky130_fd_sc_hd__dfxtp_1 _7841_ (.CLK(clknet_leaf_48_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.reg_buf[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[6][28] ));
 sky130_fd_sc_hd__dfxtp_1 _7842_ (.CLK(clknet_leaf_3_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.reg_buf[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[6][29] ));
 sky130_fd_sc_hd__dfxtp_1 _7843_ (.CLK(clknet_leaf_3_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.reg_buf[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[6][30] ));
 sky130_fd_sc_hd__dfxtp_1 _7844_ (.CLK(clknet_leaf_1_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.reg_buf[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[6][31] ));
 sky130_fd_sc_hd__dfxtp_1 _7845_ (.CLK(clknet_leaf_48_clk),
    .D(_0066_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[6][0] ));
 sky130_fd_sc_hd__dfxtp_1 _7846_ (.CLK(clknet_leaf_5_clk),
    .D(_0067_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[6][1] ));
 sky130_fd_sc_hd__dfxtp_1 _7847_ (.CLK(clknet_leaf_5_clk),
    .D(_0068_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[6][2] ));
 sky130_fd_sc_hd__dfxtp_1 _7848_ (.CLK(clknet_leaf_50_clk),
    .D(_0069_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[6][3] ));
 sky130_fd_sc_hd__dfxtp_1 _7849_ (.CLK(clknet_leaf_45_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.reg_buf[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[5][0] ));
 sky130_fd_sc_hd__dfxtp_1 _7850_ (.CLK(clknet_leaf_47_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.reg_buf[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[5][1] ));
 sky130_fd_sc_hd__dfxtp_1 _7851_ (.CLK(clknet_leaf_5_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.reg_buf[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[5][2] ));
 sky130_fd_sc_hd__dfxtp_1 _7852_ (.CLK(clknet_leaf_45_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.reg_buf[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[5][3] ));
 sky130_fd_sc_hd__dfxtp_1 _7853_ (.CLK(clknet_leaf_49_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.reg_buf[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[5][8] ));
 sky130_fd_sc_hd__dfxtp_1 _7854_ (.CLK(clknet_leaf_47_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.reg_buf[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[5][9] ));
 sky130_fd_sc_hd__dfxtp_1 _7855_ (.CLK(clknet_leaf_5_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.reg_buf[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[5][10] ));
 sky130_fd_sc_hd__dfxtp_1 _7856_ (.CLK(clknet_leaf_45_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.reg_buf[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[5][11] ));
 sky130_fd_sc_hd__dfxtp_1 _7857_ (.CLK(clknet_leaf_49_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.reg_buf[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[5][12] ));
 sky130_fd_sc_hd__dfxtp_1 _7858_ (.CLK(clknet_leaf_47_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.reg_buf[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[5][13] ));
 sky130_fd_sc_hd__dfxtp_1 _7859_ (.CLK(clknet_leaf_2_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.reg_buf[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[5][14] ));
 sky130_fd_sc_hd__dfxtp_1 _7860_ (.CLK(clknet_leaf_45_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.reg_buf[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[5][15] ));
 sky130_fd_sc_hd__dfxtp_1 _7861_ (.CLK(clknet_leaf_49_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.reg_buf[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[5][16] ));
 sky130_fd_sc_hd__dfxtp_1 _7862_ (.CLK(clknet_leaf_47_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.reg_buf[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[5][17] ));
 sky130_fd_sc_hd__dfxtp_1 _7863_ (.CLK(clknet_leaf_3_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.reg_buf[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[5][18] ));
 sky130_fd_sc_hd__dfxtp_1 _7864_ (.CLK(clknet_leaf_48_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.reg_buf[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[5][19] ));
 sky130_fd_sc_hd__dfxtp_1 _7865_ (.CLK(clknet_leaf_48_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.reg_buf[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[5][20] ));
 sky130_fd_sc_hd__dfxtp_1 _7866_ (.CLK(clknet_leaf_53_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.reg_buf[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[5][21] ));
 sky130_fd_sc_hd__dfxtp_1 _7867_ (.CLK(clknet_leaf_3_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.reg_buf[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[5][22] ));
 sky130_fd_sc_hd__dfxtp_1 _7868_ (.CLK(clknet_leaf_47_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.reg_buf[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[5][23] ));
 sky130_fd_sc_hd__dfxtp_1 _7869_ (.CLK(clknet_leaf_48_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.reg_buf[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[5][24] ));
 sky130_fd_sc_hd__dfxtp_1 _7870_ (.CLK(clknet_leaf_53_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.reg_buf[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[5][25] ));
 sky130_fd_sc_hd__dfxtp_1 _7871_ (.CLK(clknet_leaf_3_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.reg_buf[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[5][26] ));
 sky130_fd_sc_hd__dfxtp_1 _7872_ (.CLK(clknet_leaf_48_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.reg_buf[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[5][27] ));
 sky130_fd_sc_hd__dfxtp_1 _7873_ (.CLK(clknet_leaf_48_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.reg_buf[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[5][28] ));
 sky130_fd_sc_hd__dfxtp_1 _7874_ (.CLK(clknet_leaf_47_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.reg_buf[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[5][29] ));
 sky130_fd_sc_hd__dfxtp_1 _7875_ (.CLK(clknet_leaf_3_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.reg_buf[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[5][30] ));
 sky130_fd_sc_hd__dfxtp_1 _7876_ (.CLK(clknet_leaf_47_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.reg_buf[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[5][31] ));
 sky130_fd_sc_hd__dfxtp_1 _7877_ (.CLK(clknet_leaf_48_clk),
    .D(_0062_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[5][0] ));
 sky130_fd_sc_hd__dfxtp_1 _7878_ (.CLK(clknet_leaf_53_clk),
    .D(_0063_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[5][1] ));
 sky130_fd_sc_hd__dfxtp_1 _7879_ (.CLK(clknet_leaf_5_clk),
    .D(_0064_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[5][2] ));
 sky130_fd_sc_hd__dfxtp_1 _7880_ (.CLK(clknet_leaf_48_clk),
    .D(_0065_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[5][3] ));
 sky130_fd_sc_hd__dfxtp_1 _7881_ (.CLK(clknet_leaf_49_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.reg_buf[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[2][0] ));
 sky130_fd_sc_hd__dfxtp_1 _7882_ (.CLK(clknet_leaf_5_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.reg_buf[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[2][1] ));
 sky130_fd_sc_hd__dfxtp_1 _7883_ (.CLK(clknet_leaf_5_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.reg_buf[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[2][2] ));
 sky130_fd_sc_hd__dfxtp_1 _7884_ (.CLK(clknet_leaf_48_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.reg_buf[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[2][3] ));
 sky130_fd_sc_hd__dfxtp_1 _7885_ (.CLK(clknet_leaf_49_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.reg_buf[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[2][8] ));
 sky130_fd_sc_hd__dfxtp_1 _7886_ (.CLK(clknet_leaf_5_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.reg_buf[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[2][9] ));
 sky130_fd_sc_hd__dfxtp_1 _7887_ (.CLK(clknet_leaf_5_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.reg_buf[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[2][10] ));
 sky130_fd_sc_hd__dfxtp_1 _7888_ (.CLK(clknet_leaf_48_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.reg_buf[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[2][11] ));
 sky130_fd_sc_hd__dfxtp_1 _7889_ (.CLK(clknet_leaf_49_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.reg_buf[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[2][12] ));
 sky130_fd_sc_hd__dfxtp_1 _7890_ (.CLK(clknet_leaf_5_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.reg_buf[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[2][13] ));
 sky130_fd_sc_hd__dfxtp_1 _7891_ (.CLK(clknet_leaf_2_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.reg_buf[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[2][14] ));
 sky130_fd_sc_hd__dfxtp_1 _7892_ (.CLK(clknet_leaf_48_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.reg_buf[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[2][15] ));
 sky130_fd_sc_hd__dfxtp_1 _7893_ (.CLK(clknet_leaf_49_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.reg_buf[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[2][16] ));
 sky130_fd_sc_hd__dfxtp_1 _7894_ (.CLK(clknet_leaf_2_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.reg_buf[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[2][17] ));
 sky130_fd_sc_hd__dfxtp_1 _7895_ (.CLK(clknet_leaf_3_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.reg_buf[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[2][18] ));
 sky130_fd_sc_hd__dfxtp_1 _7896_ (.CLK(clknet_leaf_48_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.reg_buf[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[2][19] ));
 sky130_fd_sc_hd__dfxtp_1 _7897_ (.CLK(clknet_leaf_48_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.reg_buf[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[2][20] ));
 sky130_fd_sc_hd__dfxtp_1 _7898_ (.CLK(clknet_leaf_5_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.reg_buf[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[2][21] ));
 sky130_fd_sc_hd__dfxtp_1 _7899_ (.CLK(clknet_leaf_3_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.reg_buf[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[2][22] ));
 sky130_fd_sc_hd__dfxtp_1 _7900_ (.CLK(clknet_leaf_47_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.reg_buf[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[2][23] ));
 sky130_fd_sc_hd__dfxtp_1 _7901_ (.CLK(clknet_leaf_48_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.reg_buf[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[2][24] ));
 sky130_fd_sc_hd__dfxtp_1 _7902_ (.CLK(clknet_leaf_2_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.reg_buf[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[2][25] ));
 sky130_fd_sc_hd__dfxtp_1 _7903_ (.CLK(clknet_leaf_3_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.reg_buf[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[2][26] ));
 sky130_fd_sc_hd__dfxtp_1 _7904_ (.CLK(clknet_leaf_53_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.reg_buf[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[2][27] ));
 sky130_fd_sc_hd__dfxtp_1 _7905_ (.CLK(clknet_leaf_48_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.reg_buf[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[2][28] ));
 sky130_fd_sc_hd__dfxtp_1 _7906_ (.CLK(clknet_leaf_2_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.reg_buf[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[2][29] ));
 sky130_fd_sc_hd__dfxtp_1 _7907_ (.CLK(clknet_leaf_2_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.reg_buf[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[2][30] ));
 sky130_fd_sc_hd__dfxtp_1 _7908_ (.CLK(clknet_leaf_48_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.reg_buf[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[2][31] ));
 sky130_fd_sc_hd__dfxtp_1 _7909_ (.CLK(clknet_leaf_48_clk),
    .D(_0058_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[2][0] ));
 sky130_fd_sc_hd__dfxtp_1 _7910_ (.CLK(clknet_leaf_5_clk),
    .D(_0059_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[2][1] ));
 sky130_fd_sc_hd__dfxtp_1 _7911_ (.CLK(clknet_leaf_5_clk),
    .D(_0060_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[2][2] ));
 sky130_fd_sc_hd__dfxtp_1 _7912_ (.CLK(clknet_leaf_48_clk),
    .D(_0061_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[2][3] ));
 sky130_fd_sc_hd__dfxtp_1 _7913_ (.CLK(clknet_leaf_39_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.reg_buf[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 _7914_ (.CLK(clknet_leaf_51_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.reg_buf[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _7915_ (.CLK(clknet_leaf_50_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.reg_buf[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 _7916_ (.CLK(clknet_leaf_50_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.reg_buf[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 _7917_ (.CLK(clknet_leaf_39_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.reg_buf[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[1][8] ));
 sky130_fd_sc_hd__dfxtp_1 _7918_ (.CLK(clknet_leaf_24_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.reg_buf[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[1][9] ));
 sky130_fd_sc_hd__dfxtp_1 _7919_ (.CLK(clknet_leaf_26_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.reg_buf[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[1][10] ));
 sky130_fd_sc_hd__dfxtp_1 _7920_ (.CLK(clknet_leaf_24_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.reg_buf[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[1][11] ));
 sky130_fd_sc_hd__dfxtp_1 _7921_ (.CLK(clknet_leaf_36_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.reg_buf[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[1][12] ));
 sky130_fd_sc_hd__dfxtp_1 _7922_ (.CLK(clknet_leaf_25_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.reg_buf[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[1][13] ));
 sky130_fd_sc_hd__dfxtp_1 _7923_ (.CLK(clknet_leaf_25_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.reg_buf[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[1][14] ));
 sky130_fd_sc_hd__dfxtp_1 _7924_ (.CLK(clknet_leaf_24_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.reg_buf[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[1][15] ));
 sky130_fd_sc_hd__dfxtp_1 _7925_ (.CLK(clknet_leaf_36_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.reg_buf[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[1][16] ));
 sky130_fd_sc_hd__dfxtp_1 _7926_ (.CLK(clknet_leaf_25_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.reg_buf[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[1][17] ));
 sky130_fd_sc_hd__dfxtp_1 _7927_ (.CLK(clknet_leaf_25_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.reg_buf[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[1][18] ));
 sky130_fd_sc_hd__dfxtp_1 _7928_ (.CLK(clknet_leaf_36_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.reg_buf[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[1][19] ));
 sky130_fd_sc_hd__dfxtp_1 _7929_ (.CLK(clknet_leaf_36_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.reg_buf[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[1][20] ));
 sky130_fd_sc_hd__dfxtp_1 _7930_ (.CLK(clknet_leaf_24_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.reg_buf[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[1][21] ));
 sky130_fd_sc_hd__dfxtp_1 _7931_ (.CLK(clknet_leaf_36_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.reg_buf[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[1][22] ));
 sky130_fd_sc_hd__dfxtp_1 _7932_ (.CLK(clknet_leaf_36_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.reg_buf[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[1][23] ));
 sky130_fd_sc_hd__dfxtp_1 _7933_ (.CLK(clknet_leaf_37_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.reg_buf[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[1][24] ));
 sky130_fd_sc_hd__dfxtp_1 _7934_ (.CLK(clknet_leaf_24_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.reg_buf[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[1][25] ));
 sky130_fd_sc_hd__dfxtp_1 _7935_ (.CLK(clknet_leaf_36_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.reg_buf[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[1][26] ));
 sky130_fd_sc_hd__dfxtp_1 _7936_ (.CLK(clknet_leaf_36_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.reg_buf[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[1][27] ));
 sky130_fd_sc_hd__dfxtp_1 _7937_ (.CLK(clknet_leaf_49_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.reg_buf[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[1][28] ));
 sky130_fd_sc_hd__dfxtp_1 _7938_ (.CLK(clknet_leaf_50_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.reg_buf[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[1][29] ));
 sky130_fd_sc_hd__dfxtp_1 _7939_ (.CLK(clknet_leaf_49_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.reg_buf[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[1][30] ));
 sky130_fd_sc_hd__dfxtp_1 _7940_ (.CLK(clknet_leaf_49_clk),
    .D(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.reg_buf[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[1][31] ));
 sky130_fd_sc_hd__dfxtp_1 _7941_ (.CLK(clknet_leaf_50_clk),
    .D(_0054_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 _7942_ (.CLK(clknet_leaf_50_clk),
    .D(_0055_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _7943_ (.CLK(clknet_leaf_50_clk),
    .D(_0056_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 _7944_ (.CLK(clknet_leaf_50_clk),
    .D(_0057_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.registers[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 _7945_ (.CLK(clknet_leaf_50_clk),
    .D(\i_tinyqv.cpu.i_core.cy_out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.cy ));
 sky130_fd_sc_hd__dfxtp_1 _7946_ (.CLK(clknet_leaf_51_clk),
    .D(net139),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.load_done ));
 sky130_fd_sc_hd__dfxtp_2 _7947_ (.CLK(clknet_leaf_51_clk),
    .D(_0085_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.cycle[0] ));
 sky130_fd_sc_hd__dfxtp_1 _7948_ (.CLK(clknet_leaf_51_clk),
    .D(_0086_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.cycle[1] ));
 sky130_fd_sc_hd__dfxtp_1 _7949_ (.CLK(clknet_leaf_37_clk),
    .D(_0087_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.mcause[0] ));
 sky130_fd_sc_hd__dfxtp_1 _7950_ (.CLK(clknet_leaf_38_clk),
    .D(_0088_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.mcause[1] ));
 sky130_fd_sc_hd__dfxtp_1 _7951_ (.CLK(clknet_leaf_38_clk),
    .D(_0089_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.mcause[3] ));
 sky130_fd_sc_hd__dfxtp_1 _7952_ (.CLK(clknet_leaf_23_clk),
    .D(_0090_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.mcause[4] ));
 sky130_fd_sc_hd__dfxtp_1 _7953_ (.CLK(clknet_leaf_37_clk),
    .D(_0091_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.is_double_fault_r ));
 sky130_fd_sc_hd__dfxtp_1 _7954_ (.CLK(clknet_leaf_51_clk),
    .D(_0092_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.time_hi[0] ));
 sky130_fd_sc_hd__dfxtp_1 _7955_ (.CLK(clknet_leaf_51_clk),
    .D(_0093_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.time_hi[1] ));
 sky130_fd_sc_hd__dfxtp_1 _7956_ (.CLK(clknet_leaf_51_clk),
    .D(_0094_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.time_hi[2] ));
 sky130_fd_sc_hd__dfxtp_1 _7957_ (.CLK(clknet_leaf_50_clk),
    .D(net128),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.add ));
 sky130_fd_sc_hd__dfxtp_1 _7958_ (.CLK(clknet_leaf_26_clk),
    .D(_0095_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.last_interrupt_req[0] ));
 sky130_fd_sc_hd__dfxtp_1 _7959_ (.CLK(clknet_leaf_26_clk),
    .D(_0096_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.last_interrupt_req[1] ));
 sky130_fd_sc_hd__dfxtp_1 _7960_ (.CLK(clknet_leaf_36_clk),
    .D(_0097_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.mepc[20] ));
 sky130_fd_sc_hd__dfxtp_1 _7961_ (.CLK(clknet_leaf_35_clk),
    .D(_0098_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.mepc[21] ));
 sky130_fd_sc_hd__dfxtp_1 _7962_ (.CLK(clknet_leaf_35_clk),
    .D(_0099_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.mepc[22] ));
 sky130_fd_sc_hd__dfxtp_1 _7963_ (.CLK(clknet_leaf_35_clk),
    .D(_0100_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.mepc[23] ));
 sky130_fd_sc_hd__dfxtp_1 _7964_ (.CLK(clknet_leaf_38_clk),
    .D(_0101_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.mstatus_mpie ));
 sky130_fd_sc_hd__dfxtp_1 _7965_ (.CLK(clknet_leaf_37_clk),
    .D(_0102_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.mstatus_mie ));
 sky130_fd_sc_hd__dfxtp_1 _7966_ (.CLK(clknet_leaf_37_clk),
    .D(_0103_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.mstatus_mte ));
 sky130_fd_sc_hd__dfxtp_1 _7967_ (.CLK(clknet_leaf_5_clk),
    .D(_0104_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.rd[0] ));
 sky130_fd_sc_hd__dfxtp_2 _7968_ (.CLK(clknet_leaf_5_clk),
    .D(_0105_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.rd[1] ));
 sky130_fd_sc_hd__dfxtp_2 _7969_ (.CLK(clknet_leaf_6_clk),
    .D(_0106_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.rd[2] ));
 sky130_fd_sc_hd__dfxtp_2 _7970_ (.CLK(clknet_leaf_6_clk),
    .D(_0107_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.rd[3] ));
 sky130_fd_sc_hd__dfxtp_1 _7971_ (.CLK(clknet_leaf_50_clk),
    .D(\i_tinyqv.cpu.i_core.cmp_out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.cmp ));
 sky130_fd_sc_hd__dfxtp_2 _7972_ (.CLK(clknet_leaf_17_clk),
    .D(\i_debug_uart_tx.resetn ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.rstn ));
 sky130_fd_sc_hd__dfxtp_1 _7973_ (.CLK(clknet_leaf_29_clk),
    .D(_0108_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_uart_tx.data_to_send[0] ));
 sky130_fd_sc_hd__dfxtp_1 _7974_ (.CLK(clknet_leaf_29_clk),
    .D(_0109_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_uart_tx.data_to_send[1] ));
 sky130_fd_sc_hd__dfxtp_1 _7975_ (.CLK(clknet_leaf_29_clk),
    .D(_0110_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_uart_tx.data_to_send[2] ));
 sky130_fd_sc_hd__dfxtp_1 _7976_ (.CLK(clknet_leaf_28_clk),
    .D(_0111_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_uart_tx.data_to_send[3] ));
 sky130_fd_sc_hd__dfxtp_1 _7977_ (.CLK(clknet_leaf_28_clk),
    .D(_0112_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_uart_tx.data_to_send[4] ));
 sky130_fd_sc_hd__dfxtp_1 _7978_ (.CLK(clknet_leaf_28_clk),
    .D(_0113_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_uart_tx.data_to_send[5] ));
 sky130_fd_sc_hd__dfxtp_1 _7979_ (.CLK(clknet_leaf_28_clk),
    .D(_0114_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_uart_tx.data_to_send[6] ));
 sky130_fd_sc_hd__dfxtp_1 _7980_ (.CLK(clknet_leaf_28_clk),
    .D(_0115_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_uart_tx.data_to_send[7] ));
 sky130_fd_sc_hd__dfxtp_1 _7981_ (.CLK(clknet_leaf_32_clk),
    .D(_0116_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_uart_tx.cycle_counter[0] ));
 sky130_fd_sc_hd__dfxtp_1 _7982_ (.CLK(clknet_leaf_31_clk),
    .D(_0117_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_uart_tx.cycle_counter[1] ));
 sky130_fd_sc_hd__dfxtp_1 _7983_ (.CLK(clknet_leaf_32_clk),
    .D(_0118_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_uart_tx.cycle_counter[2] ));
 sky130_fd_sc_hd__dfxtp_1 _7984_ (.CLK(clknet_leaf_32_clk),
    .D(_0119_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_uart_tx.cycle_counter[3] ));
 sky130_fd_sc_hd__dfxtp_1 _7985_ (.CLK(clknet_leaf_32_clk),
    .D(_0120_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_uart_tx.cycle_counter[4] ));
 sky130_fd_sc_hd__dfxtp_1 _7986_ (.CLK(clknet_leaf_31_clk),
    .D(_0121_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_uart_tx.cycle_counter[5] ));
 sky130_fd_sc_hd__dfxtp_1 _7987_ (.CLK(clknet_leaf_31_clk),
    .D(_0122_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_uart_tx.cycle_counter[6] ));
 sky130_fd_sc_hd__dfxtp_1 _7988_ (.CLK(clknet_leaf_31_clk),
    .D(_0123_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_uart_tx.cycle_counter[7] ));
 sky130_fd_sc_hd__dfxtp_1 _7989_ (.CLK(clknet_leaf_31_clk),
    .D(_0124_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_uart_tx.cycle_counter[8] ));
 sky130_fd_sc_hd__dfxtp_1 _7990_ (.CLK(clknet_leaf_30_clk),
    .D(_0125_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_uart_tx.cycle_counter[9] ));
 sky130_fd_sc_hd__dfxtp_1 _7991_ (.CLK(clknet_leaf_31_clk),
    .D(_0126_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_uart_tx.cycle_counter[10] ));
 sky130_fd_sc_hd__dfxtp_2 _7992_ (.CLK(clknet_leaf_32_clk),
    .D(_0127_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_uart_tx.fsm_state[0] ));
 sky130_fd_sc_hd__dfxtp_1 _7993_ (.CLK(clknet_leaf_29_clk),
    .D(_0128_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_uart_tx.fsm_state[1] ));
 sky130_fd_sc_hd__dfxtp_2 _7994_ (.CLK(clknet_leaf_29_clk),
    .D(_0129_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_uart_tx.fsm_state[2] ));
 sky130_fd_sc_hd__dfxtp_1 _7995_ (.CLK(clknet_leaf_30_clk),
    .D(net166),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_uart_tx.fsm_state[3] ));
 sky130_fd_sc_hd__dfxtp_1 _7996_ (.CLK(clknet_leaf_31_clk),
    .D(_0131_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_uart_rx.cycle_counter[0] ));
 sky130_fd_sc_hd__dfxtp_1 _7997_ (.CLK(clknet_leaf_30_clk),
    .D(_0132_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_uart_rx.cycle_counter[1] ));
 sky130_fd_sc_hd__dfxtp_1 _7998_ (.CLK(clknet_leaf_31_clk),
    .D(_0133_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_uart_rx.cycle_counter[2] ));
 sky130_fd_sc_hd__dfxtp_1 _7999_ (.CLK(clknet_leaf_30_clk),
    .D(_0134_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_uart_rx.cycle_counter[3] ));
 sky130_fd_sc_hd__dfxtp_1 _8000_ (.CLK(clknet_leaf_31_clk),
    .D(_0135_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_uart_rx.cycle_counter[4] ));
 sky130_fd_sc_hd__dfxtp_1 _8001_ (.CLK(clknet_leaf_30_clk),
    .D(_0136_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_uart_rx.cycle_counter[5] ));
 sky130_fd_sc_hd__dfxtp_1 _8002_ (.CLK(clknet_leaf_30_clk),
    .D(_0137_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_uart_rx.cycle_counter[6] ));
 sky130_fd_sc_hd__dfxtp_1 _8003_ (.CLK(clknet_leaf_30_clk),
    .D(_0138_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_uart_rx.cycle_counter[7] ));
 sky130_fd_sc_hd__dfxtp_1 _8004_ (.CLK(clknet_leaf_30_clk),
    .D(_0139_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_uart_rx.cycle_counter[8] ));
 sky130_fd_sc_hd__dfxtp_1 _8005_ (.CLK(clknet_leaf_30_clk),
    .D(_0140_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_uart_rx.cycle_counter[9] ));
 sky130_fd_sc_hd__dfxtp_1 _8006_ (.CLK(clknet_leaf_30_clk),
    .D(_0141_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_uart_rx.cycle_counter[10] ));
 sky130_fd_sc_hd__dfxtp_1 _8007_ (.CLK(clknet_leaf_27_clk),
    .D(net202),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_uart_rx.recieved_data[0] ));
 sky130_fd_sc_hd__dfxtp_1 _8008_ (.CLK(clknet_leaf_19_clk),
    .D(_0143_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_uart_rx.recieved_data[1] ));
 sky130_fd_sc_hd__dfxtp_1 _8009_ (.CLK(clknet_leaf_19_clk),
    .D(_0144_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_uart_rx.recieved_data[2] ));
 sky130_fd_sc_hd__dfxtp_1 _8010_ (.CLK(clknet_leaf_19_clk),
    .D(_0145_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_uart_rx.recieved_data[3] ));
 sky130_fd_sc_hd__dfxtp_1 _8011_ (.CLK(clknet_leaf_18_clk),
    .D(_0146_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_uart_rx.recieved_data[4] ));
 sky130_fd_sc_hd__dfxtp_1 _8012_ (.CLK(clknet_leaf_19_clk),
    .D(_0147_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_uart_rx.recieved_data[5] ));
 sky130_fd_sc_hd__dfxtp_1 _8013_ (.CLK(clknet_leaf_19_clk),
    .D(_0148_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_uart_rx.recieved_data[6] ));
 sky130_fd_sc_hd__dfxtp_1 _8014_ (.CLK(clknet_leaf_28_clk),
    .D(_0149_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_uart_rx.recieved_data[7] ));
 sky130_fd_sc_hd__dfxtp_1 _8015_ (.CLK(clknet_leaf_27_clk),
    .D(_0150_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_uart_rx.bit_sample ));
 sky130_fd_sc_hd__dfxtp_1 _8016_ (.CLK(clknet_leaf_27_clk),
    .D(_0151_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_uart_rx.uart_rts ));
 sky130_fd_sc_hd__dfxtp_2 _8017_ (.CLK(clknet_leaf_27_clk),
    .D(_0152_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_uart_rx.fsm_state[0] ));
 sky130_fd_sc_hd__dfxtp_2 _8018_ (.CLK(clknet_leaf_28_clk),
    .D(_0153_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_uart_rx.fsm_state[1] ));
 sky130_fd_sc_hd__dfxtp_1 _8019_ (.CLK(clknet_leaf_30_clk),
    .D(_0154_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_uart_rx.fsm_state[2] ));
 sky130_fd_sc_hd__dfxtp_2 _8020_ (.CLK(clknet_leaf_30_clk),
    .D(_0155_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_uart_rx.fsm_state[3] ));
 sky130_fd_sc_hd__dfxtp_1 _8021_ (.CLK(clknet_leaf_27_clk),
    .D(_0156_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_uart_rx.rxd_reg[0] ));
 sky130_fd_sc_hd__dfxtp_1 _8022_ (.CLK(clknet_leaf_27_clk),
    .D(_0157_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_uart_rx.rxd_reg[1] ));
 sky130_fd_sc_hd__dfxtp_1 _8023_ (.CLK(clknet_leaf_16_clk),
    .D(_0158_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.mem.q_ctrl.stop_txn_reg ));
 sky130_fd_sc_hd__dfxtp_1 _8024_ (.CLK(clknet_leaf_13_clk),
    .D(_0159_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.instr_data[3][2] ));
 sky130_fd_sc_hd__dfxtp_1 _8025_ (.CLK(clknet_leaf_13_clk),
    .D(_0160_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.instr_data[3][3] ));
 sky130_fd_sc_hd__dfxtp_1 _8026_ (.CLK(clknet_leaf_10_clk),
    .D(_0161_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.instr_data[3][4] ));
 sky130_fd_sc_hd__dfxtp_1 _8027_ (.CLK(clknet_leaf_3_clk),
    .D(_0162_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.instr_data[3][5] ));
 sky130_fd_sc_hd__dfxtp_1 _8028_ (.CLK(clknet_leaf_4_clk),
    .D(_0163_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.instr_data[3][6] ));
 sky130_fd_sc_hd__dfxtp_1 _8029_ (.CLK(clknet_leaf_10_clk),
    .D(_0164_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.instr_data[3][7] ));
 sky130_fd_sc_hd__dfxtp_1 _8030_ (.CLK(clknet_leaf_11_clk),
    .D(_0165_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.instr_data[3][8] ));
 sky130_fd_sc_hd__dfxtp_1 _8031_ (.CLK(clknet_leaf_10_clk),
    .D(_0166_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.instr_data[3][9] ));
 sky130_fd_sc_hd__dfxtp_1 _8032_ (.CLK(clknet_leaf_4_clk),
    .D(_0167_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.instr_data[3][10] ));
 sky130_fd_sc_hd__dfxtp_1 _8033_ (.CLK(clknet_leaf_11_clk),
    .D(_0168_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.instr_data[3][11] ));
 sky130_fd_sc_hd__dfxtp_1 _8034_ (.CLK(clknet_leaf_11_clk),
    .D(_0169_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.instr_data[3][12] ));
 sky130_fd_sc_hd__dfxtp_1 _8035_ (.CLK(clknet_leaf_12_clk),
    .D(_0170_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.instr_data[3][13] ));
 sky130_fd_sc_hd__dfxtp_1 _8036_ (.CLK(clknet_leaf_11_clk),
    .D(_0171_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.instr_data[3][14] ));
 sky130_fd_sc_hd__dfxtp_1 _8037_ (.CLK(clknet_leaf_12_clk),
    .D(_0172_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.instr_data[3][15] ));
 sky130_fd_sc_hd__dfxtp_1 _8038_ (.CLK(clknet_leaf_29_clk),
    .D(_0173_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_debug_uart_tx.data_to_send[0] ));
 sky130_fd_sc_hd__dfxtp_1 _8039_ (.CLK(clknet_leaf_29_clk),
    .D(_0174_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_debug_uart_tx.data_to_send[1] ));
 sky130_fd_sc_hd__dfxtp_1 _8040_ (.CLK(clknet_leaf_29_clk),
    .D(_0175_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_debug_uart_tx.data_to_send[2] ));
 sky130_fd_sc_hd__dfxtp_1 _8041_ (.CLK(clknet_leaf_28_clk),
    .D(_0176_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_debug_uart_tx.data_to_send[3] ));
 sky130_fd_sc_hd__dfxtp_1 _8042_ (.CLK(clknet_leaf_28_clk),
    .D(_0177_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_debug_uart_tx.data_to_send[4] ));
 sky130_fd_sc_hd__dfxtp_1 _8043_ (.CLK(clknet_leaf_28_clk),
    .D(_0178_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_debug_uart_tx.data_to_send[5] ));
 sky130_fd_sc_hd__dfxtp_1 _8044_ (.CLK(clknet_leaf_28_clk),
    .D(_0179_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_debug_uart_tx.data_to_send[6] ));
 sky130_fd_sc_hd__dfxtp_1 _8045_ (.CLK(clknet_leaf_28_clk),
    .D(_0180_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_debug_uart_tx.data_to_send[7] ));
 sky130_fd_sc_hd__dfxtp_1 _8046_ (.CLK(clknet_leaf_30_clk),
    .D(_0181_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_debug_uart_tx.cycle_counter[0] ));
 sky130_fd_sc_hd__dfxtp_1 _8047_ (.CLK(clknet_leaf_30_clk),
    .D(_0182_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_debug_uart_tx.cycle_counter[1] ));
 sky130_fd_sc_hd__dfxtp_1 _8048_ (.CLK(clknet_leaf_30_clk),
    .D(_0183_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_debug_uart_tx.cycle_counter[2] ));
 sky130_fd_sc_hd__dfxtp_1 _8049_ (.CLK(clknet_leaf_30_clk),
    .D(_0184_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_debug_uart_tx.cycle_counter[3] ));
 sky130_fd_sc_hd__dfxtp_1 _8050_ (.CLK(clknet_leaf_30_clk),
    .D(_0185_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_debug_uart_tx.cycle_counter[4] ));
 sky130_fd_sc_hd__dfxtp_2 _8051_ (.CLK(clknet_leaf_30_clk),
    .D(_0186_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_debug_uart_tx.fsm_state[0] ));
 sky130_fd_sc_hd__dfxtp_1 _8052_ (.CLK(clknet_leaf_30_clk),
    .D(_0187_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_debug_uart_tx.fsm_state[1] ));
 sky130_fd_sc_hd__dfxtp_1 _8053_ (.CLK(clknet_leaf_30_clk),
    .D(_0188_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_debug_uart_tx.fsm_state[2] ));
 sky130_fd_sc_hd__dfxtp_1 _8054_ (.CLK(clknet_leaf_30_clk),
    .D(_0189_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_debug_uart_tx.fsm_state[3] ));
 sky130_fd_sc_hd__dfxtp_1 _8055_ (.CLK(clknet_leaf_27_clk),
    .D(_0190_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_spi.clock_count[0] ));
 sky130_fd_sc_hd__dfxtp_1 _8056_ (.CLK(clknet_leaf_27_clk),
    .D(_0191_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_spi.clock_count[1] ));
 sky130_fd_sc_hd__dfxtp_1 _8057_ (.CLK(clknet_leaf_27_clk),
    .D(_0192_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_spi.data[0] ));
 sky130_fd_sc_hd__dfxtp_1 _8058_ (.CLK(clknet_leaf_28_clk),
    .D(_0193_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_spi.bits_remaining[0] ));
 sky130_fd_sc_hd__dfxtp_1 _8059_ (.CLK(clknet_leaf_28_clk),
    .D(_0194_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_spi.bits_remaining[1] ));
 sky130_fd_sc_hd__dfxtp_1 _8060_ (.CLK(clknet_leaf_25_clk),
    .D(_0195_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_spi.bits_remaining[2] ));
 sky130_fd_sc_hd__dfxtp_1 _8061_ (.CLK(clknet_leaf_26_clk),
    .D(net195),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_spi.bits_remaining[3] ));
 sky130_fd_sc_hd__dfxtp_1 _8062_ (.CLK(clknet_leaf_27_clk),
    .D(_0197_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_spi.busy ));
 sky130_fd_sc_hd__dfxtp_1 _8063_ (.CLK(clknet_leaf_26_clk),
    .D(_0198_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_spi.spi_dc ));
 sky130_fd_sc_hd__dfxtp_1 _8064_ (.CLK(clknet_leaf_26_clk),
    .D(net185),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_spi.spi_select ));
 sky130_fd_sc_hd__dfxtp_1 _8065_ (.CLK(clknet_leaf_27_clk),
    .D(_0200_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_spi.spi_clk_out ));
 sky130_fd_sc_hd__dfxtp_1 _8066_ (.CLK(clknet_leaf_30_clk),
    .D(_0201_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_debug_uart_tx.txd_reg ));
 sky130_fd_sc_hd__dfxtp_1 _8067_ (.CLK(clknet_leaf_27_clk),
    .D(_0202_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_spi.read_latency ));
 sky130_fd_sc_hd__dfxtp_1 _8068_ (.CLK(clknet_leaf_27_clk),
    .D(net163),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_spi.clock_divider[0] ));
 sky130_fd_sc_hd__dfxtp_1 _8069_ (.CLK(clknet_leaf_27_clk),
    .D(_0204_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_spi.clock_divider[1] ));
 sky130_fd_sc_hd__dfxtp_1 _8070_ (.CLK(clknet_leaf_23_clk),
    .D(_0205_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.mip[17] ));
 sky130_fd_sc_hd__dfxtp_1 _8071_ (.CLK(clknet_leaf_23_clk),
    .D(_0206_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.mip[16] ));
 sky130_fd_sc_hd__dfxtp_1 _8072_ (.CLK(clknet_leaf_37_clk),
    .D(_0207_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.mie[19] ));
 sky130_fd_sc_hd__dfxtp_1 _8073_ (.CLK(clknet_leaf_38_clk),
    .D(_0208_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.mie[18] ));
 sky130_fd_sc_hd__dfxtp_1 _8074_ (.CLK(clknet_leaf_37_clk),
    .D(_0209_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.mie[17] ));
 sky130_fd_sc_hd__dfxtp_1 _8075_ (.CLK(clknet_leaf_37_clk),
    .D(_0210_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.mie[16] ));
 sky130_fd_sc_hd__dfxtp_1 _8076_ (.CLK(clknet_leaf_51_clk),
    .D(\i_tinyqv.cpu.debug_rd[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\debug_rd_r[0] ));
 sky130_fd_sc_hd__dfxtp_1 _8077_ (.CLK(clknet_leaf_52_clk),
    .D(\i_tinyqv.cpu.debug_rd[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\debug_rd_r[1] ));
 sky130_fd_sc_hd__dfxtp_1 _8078_ (.CLK(clknet_leaf_51_clk),
    .D(\i_tinyqv.cpu.debug_rd[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\debug_rd_r[2] ));
 sky130_fd_sc_hd__dfxtp_1 _8079_ (.CLK(clknet_leaf_53_clk),
    .D(net32),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\debug_rd_r[3] ));
 sky130_fd_sc_hd__dfxtp_1 _8080_ (.CLK(clknet_leaf_29_clk),
    .D(_0211_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_uart_tx.txd_reg ));
 sky130_fd_sc_hd__dfxtp_1 _8081_ (.CLK(clknet_leaf_19_clk),
    .D(_0008_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\gpio_out_sel[0] ));
 sky130_fd_sc_hd__dfxtp_1 _8082_ (.CLK(clknet_leaf_19_clk),
    .D(_0009_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\gpio_out_sel[1] ));
 sky130_fd_sc_hd__dfxtp_1 _8083_ (.CLK(clknet_leaf_18_clk),
    .D(_0010_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\gpio_out_sel[2] ));
 sky130_fd_sc_hd__dfxtp_1 _8084_ (.CLK(clknet_leaf_18_clk),
    .D(_0011_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\gpio_out_sel[3] ));
 sky130_fd_sc_hd__dfxtp_1 _8085_ (.CLK(clknet_leaf_18_clk),
    .D(_0012_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\gpio_out_sel[4] ));
 sky130_fd_sc_hd__dfxtp_1 _8086_ (.CLK(clknet_leaf_18_clk),
    .D(_0013_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\gpio_out_sel[5] ));
 sky130_fd_sc_hd__dfxtp_1 _8087_ (.CLK(clknet_leaf_18_clk),
    .D(_0014_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\gpio_out_sel[6] ));
 sky130_fd_sc_hd__dfxtp_1 _8088_ (.CLK(clknet_leaf_17_clk),
    .D(_0015_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\gpio_out_sel[7] ));
 sky130_fd_sc_hd__dfxtp_1 _8089_ (.CLK(clknet_leaf_27_clk),
    .D(_0000_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\gpio_out[0] ));
 sky130_fd_sc_hd__dfxtp_1 _8090_ (.CLK(clknet_leaf_27_clk),
    .D(_0001_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\gpio_out[1] ));
 sky130_fd_sc_hd__dfxtp_1 _8091_ (.CLK(clknet_leaf_19_clk),
    .D(_0002_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\gpio_out[2] ));
 sky130_fd_sc_hd__dfxtp_1 _8092_ (.CLK(clknet_leaf_18_clk),
    .D(_0003_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\gpio_out[3] ));
 sky130_fd_sc_hd__dfxtp_1 _8093_ (.CLK(clknet_leaf_18_clk),
    .D(_0004_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\gpio_out[4] ));
 sky130_fd_sc_hd__dfxtp_1 _8094_ (.CLK(clknet_leaf_17_clk),
    .D(_0005_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\gpio_out[5] ));
 sky130_fd_sc_hd__dfxtp_1 _8095_ (.CLK(clknet_leaf_18_clk),
    .D(_0006_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\gpio_out[6] ));
 sky130_fd_sc_hd__dfxtp_1 _8096_ (.CLK(clknet_leaf_17_clk),
    .D(_0007_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\gpio_out[7] ));
 sky130_fd_sc_hd__dfxtp_1 _8097_ (.CLK(clknet_leaf_26_clk),
    .D(net2),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.interrupt_req[0] ));
 sky130_fd_sc_hd__dfxtp_1 _8098_ (.CLK(clknet_leaf_18_clk),
    .D(net3),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.interrupt_req[1] ));
 sky130_fd_sc_hd__dfxtp_1 _8099_ (.CLK(net29),
    .D(net1),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_debug_uart_tx.resetn ));
 sky130_fd_sc_hd__dfxtp_1 _8100_ (.CLK(clknet_leaf_8_clk),
    .D(_0212_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.instr_data[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 _8101_ (.CLK(clknet_leaf_9_clk),
    .D(_0213_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.instr_data[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _8102_ (.CLK(clknet_leaf_11_clk),
    .D(_0214_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.instr_data[0][2] ));
 sky130_fd_sc_hd__dfxtp_1 _8103_ (.CLK(clknet_leaf_12_clk),
    .D(_0215_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.instr_data[0][3] ));
 sky130_fd_sc_hd__dfxtp_1 _8104_ (.CLK(clknet_leaf_10_clk),
    .D(_0216_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.instr_data[0][4] ));
 sky130_fd_sc_hd__dfxtp_1 _8105_ (.CLK(clknet_leaf_3_clk),
    .D(_0217_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.instr_data[0][5] ));
 sky130_fd_sc_hd__dfxtp_1 _8106_ (.CLK(clknet_leaf_4_clk),
    .D(_0218_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.instr_data[0][6] ));
 sky130_fd_sc_hd__dfxtp_1 _8107_ (.CLK(clknet_leaf_10_clk),
    .D(_0219_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.instr_data[0][7] ));
 sky130_fd_sc_hd__dfxtp_1 _8108_ (.CLK(clknet_leaf_11_clk),
    .D(_0220_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.instr_data[0][8] ));
 sky130_fd_sc_hd__dfxtp_1 _8109_ (.CLK(clknet_leaf_10_clk),
    .D(_0221_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.instr_data[0][9] ));
 sky130_fd_sc_hd__dfxtp_1 _8110_ (.CLK(clknet_leaf_4_clk),
    .D(_0222_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.instr_data[0][10] ));
 sky130_fd_sc_hd__dfxtp_1 _8111_ (.CLK(clknet_leaf_11_clk),
    .D(_0223_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.instr_data[0][11] ));
 sky130_fd_sc_hd__dfxtp_1 _8112_ (.CLK(clknet_leaf_9_clk),
    .D(_0224_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.instr_data[0][12] ));
 sky130_fd_sc_hd__dfxtp_1 _8113_ (.CLK(clknet_leaf_13_clk),
    .D(_0225_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.instr_data[0][13] ));
 sky130_fd_sc_hd__dfxtp_1 _8114_ (.CLK(clknet_leaf_12_clk),
    .D(_0226_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.instr_data[0][14] ));
 sky130_fd_sc_hd__dfxtp_1 _8115_ (.CLK(clknet_leaf_12_clk),
    .D(_0227_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.instr_data[0][15] ));
 sky130_fd_sc_hd__dfxtp_1 _8116_ (.CLK(clknet_leaf_9_clk),
    .D(_0228_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.instr_data[3][0] ));
 sky130_fd_sc_hd__dfxtp_1 _8117_ (.CLK(clknet_leaf_9_clk),
    .D(_0229_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.instr_data[3][1] ));
 sky130_fd_sc_hd__dfxtp_1 _8118_ (.CLK(clknet_leaf_27_clk),
    .D(_0230_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_spi.data[1] ));
 sky130_fd_sc_hd__dfxtp_1 _8119_ (.CLK(clknet_leaf_19_clk),
    .D(_0231_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_spi.data[2] ));
 sky130_fd_sc_hd__dfxtp_1 _8120_ (.CLK(clknet_leaf_18_clk),
    .D(_0232_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_spi.data[3] ));
 sky130_fd_sc_hd__dfxtp_1 _8121_ (.CLK(clknet_leaf_18_clk),
    .D(_0233_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_spi.data[4] ));
 sky130_fd_sc_hd__dfxtp_1 _8122_ (.CLK(clknet_leaf_18_clk),
    .D(_0234_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_spi.data[5] ));
 sky130_fd_sc_hd__dfxtp_1 _8123_ (.CLK(clknet_leaf_18_clk),
    .D(_0235_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_spi.data[6] ));
 sky130_fd_sc_hd__dfxtp_1 _8124_ (.CLK(clknet_leaf_18_clk),
    .D(_0236_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_spi.data[7] ));
 sky130_fd_sc_hd__dfxtp_1 _8125_ (.CLK(clknet_leaf_29_clk),
    .D(_0237_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.data_addr[0] ));
 sky130_fd_sc_hd__dfxtp_1 _8126_ (.CLK(clknet_leaf_33_clk),
    .D(_0238_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.data_addr[1] ));
 sky130_fd_sc_hd__dfxtp_2 _8127_ (.CLK(clknet_leaf_25_clk),
    .D(_0239_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.data_addr[2] ));
 sky130_fd_sc_hd__dfxtp_1 _8128_ (.CLK(clknet_leaf_28_clk),
    .D(_0240_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.data_addr[3] ));
 sky130_fd_sc_hd__dfxtp_1 _8129_ (.CLK(clknet_leaf_28_clk),
    .D(_0241_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.data_addr[4] ));
 sky130_fd_sc_hd__dfxtp_1 _8130_ (.CLK(clknet_leaf_25_clk),
    .D(_0242_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.data_addr[5] ));
 sky130_fd_sc_hd__dfxtp_1 _8131_ (.CLK(clknet_leaf_32_clk),
    .D(_0243_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.data_addr[6] ));
 sky130_fd_sc_hd__dfxtp_1 _8132_ (.CLK(clknet_leaf_33_clk),
    .D(_0244_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.data_addr[7] ));
 sky130_fd_sc_hd__dfxtp_1 _8133_ (.CLK(clknet_leaf_32_clk),
    .D(_0245_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.data_addr[8] ));
 sky130_fd_sc_hd__dfxtp_1 _8134_ (.CLK(clknet_leaf_32_clk),
    .D(_0246_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.data_addr[9] ));
 sky130_fd_sc_hd__dfxtp_1 _8135_ (.CLK(clknet_leaf_34_clk),
    .D(_0247_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.data_addr[10] ));
 sky130_fd_sc_hd__dfxtp_1 _8136_ (.CLK(clknet_leaf_33_clk),
    .D(_0248_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.data_addr[11] ));
 sky130_fd_sc_hd__dfxtp_1 _8137_ (.CLK(clknet_leaf_34_clk),
    .D(_0249_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.data_addr[12] ));
 sky130_fd_sc_hd__dfxtp_1 _8138_ (.CLK(clknet_leaf_34_clk),
    .D(_0250_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.data_addr[13] ));
 sky130_fd_sc_hd__dfxtp_1 _8139_ (.CLK(clknet_leaf_34_clk),
    .D(_0251_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.data_addr[14] ));
 sky130_fd_sc_hd__dfxtp_1 _8140_ (.CLK(clknet_leaf_34_clk),
    .D(_0252_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.data_addr[15] ));
 sky130_fd_sc_hd__dfxtp_1 _8141_ (.CLK(clknet_leaf_34_clk),
    .D(_0253_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.data_addr[16] ));
 sky130_fd_sc_hd__dfxtp_1 _8142_ (.CLK(clknet_leaf_34_clk),
    .D(_0254_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.data_addr[17] ));
 sky130_fd_sc_hd__dfxtp_1 _8143_ (.CLK(clknet_leaf_34_clk),
    .D(_0255_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.data_addr[18] ));
 sky130_fd_sc_hd__dfxtp_1 _8144_ (.CLK(clknet_leaf_34_clk),
    .D(_0256_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.data_addr[19] ));
 sky130_fd_sc_hd__dfxtp_1 _8145_ (.CLK(clknet_leaf_32_clk),
    .D(_0257_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.data_addr[20] ));
 sky130_fd_sc_hd__dfxtp_1 _8146_ (.CLK(clknet_leaf_35_clk),
    .D(_0258_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.data_addr[21] ));
 sky130_fd_sc_hd__dfxtp_1 _8147_ (.CLK(clknet_leaf_34_clk),
    .D(_0259_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.data_addr[22] ));
 sky130_fd_sc_hd__dfxtp_4 _8148_ (.CLK(clknet_leaf_35_clk),
    .D(_0260_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.data_addr[23] ));
 sky130_fd_sc_hd__dfxtp_4 _8149_ (.CLK(clknet_leaf_40_clk),
    .D(_0261_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.data_addr[24] ));
 sky130_fd_sc_hd__dfxtp_1 _8150_ (.CLK(clknet_leaf_40_clk),
    .D(_0262_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.data_addr[25] ));
 sky130_fd_sc_hd__dfxtp_1 _8151_ (.CLK(clknet_leaf_35_clk),
    .D(_0263_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.data_addr[26] ));
 sky130_fd_sc_hd__dfxtp_1 _8152_ (.CLK(clknet_leaf_35_clk),
    .D(_0264_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.data_addr[27] ));
 sky130_fd_sc_hd__dfxtp_1 _8153_ (.CLK(clknet_leaf_11_clk),
    .D(_0265_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.instr_data[2][2] ));
 sky130_fd_sc_hd__dfxtp_1 _8154_ (.CLK(clknet_leaf_11_clk),
    .D(_0266_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.instr_data[2][3] ));
 sky130_fd_sc_hd__dfxtp_1 _8155_ (.CLK(clknet_leaf_10_clk),
    .D(_0267_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.instr_data[2][4] ));
 sky130_fd_sc_hd__dfxtp_1 _8156_ (.CLK(clknet_leaf_3_clk),
    .D(_0268_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.instr_data[2][5] ));
 sky130_fd_sc_hd__dfxtp_1 _8157_ (.CLK(clknet_leaf_4_clk),
    .D(_0269_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.instr_data[2][6] ));
 sky130_fd_sc_hd__dfxtp_1 _8158_ (.CLK(clknet_leaf_10_clk),
    .D(_0270_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.instr_data[2][7] ));
 sky130_fd_sc_hd__dfxtp_1 _8159_ (.CLK(clknet_leaf_11_clk),
    .D(_0271_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.instr_data[2][8] ));
 sky130_fd_sc_hd__dfxtp_1 _8160_ (.CLK(clknet_leaf_10_clk),
    .D(_0272_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.instr_data[2][9] ));
 sky130_fd_sc_hd__dfxtp_1 _8161_ (.CLK(clknet_leaf_3_clk),
    .D(_0273_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.instr_data[2][10] ));
 sky130_fd_sc_hd__dfxtp_1 _8162_ (.CLK(clknet_leaf_11_clk),
    .D(_0274_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.instr_data[2][11] ));
 sky130_fd_sc_hd__dfxtp_1 _8163_ (.CLK(clknet_leaf_11_clk),
    .D(_0275_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.instr_data[2][12] ));
 sky130_fd_sc_hd__dfxtp_1 _8164_ (.CLK(clknet_leaf_12_clk),
    .D(_0276_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.instr_data[2][13] ));
 sky130_fd_sc_hd__dfxtp_1 _8165_ (.CLK(clknet_leaf_12_clk),
    .D(_0277_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.instr_data[2][14] ));
 sky130_fd_sc_hd__dfxtp_1 _8166_ (.CLK(clknet_leaf_14_clk),
    .D(_0278_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.instr_data[2][15] ));
 sky130_fd_sc_hd__dfxtp_1 _8167_ (.CLK(clknet_leaf_13_clk),
    .D(_0279_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.instr_data[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 _8168_ (.CLK(clknet_leaf_13_clk),
    .D(_0280_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.instr_data[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 _8169_ (.CLK(clknet_leaf_10_clk),
    .D(_0281_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.instr_data[1][4] ));
 sky130_fd_sc_hd__dfxtp_1 _8170_ (.CLK(clknet_leaf_10_clk),
    .D(_0282_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.instr_data[1][5] ));
 sky130_fd_sc_hd__dfxtp_1 _8171_ (.CLK(clknet_leaf_10_clk),
    .D(_0283_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.instr_data[1][6] ));
 sky130_fd_sc_hd__dfxtp_1 _8172_ (.CLK(clknet_leaf_10_clk),
    .D(_0284_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.instr_data[1][7] ));
 sky130_fd_sc_hd__dfxtp_1 _8173_ (.CLK(clknet_leaf_11_clk),
    .D(_0285_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.instr_data[1][8] ));
 sky130_fd_sc_hd__dfxtp_1 _8174_ (.CLK(clknet_leaf_10_clk),
    .D(_0286_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.instr_data[1][9] ));
 sky130_fd_sc_hd__dfxtp_1 _8175_ (.CLK(clknet_leaf_10_clk),
    .D(_0287_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.instr_data[1][10] ));
 sky130_fd_sc_hd__dfxtp_1 _8176_ (.CLK(clknet_leaf_11_clk),
    .D(_0288_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.instr_data[1][11] ));
 sky130_fd_sc_hd__dfxtp_1 _8177_ (.CLK(clknet_leaf_10_clk),
    .D(_0289_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.instr_data[1][12] ));
 sky130_fd_sc_hd__dfxtp_1 _8178_ (.CLK(clknet_leaf_13_clk),
    .D(_0290_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.instr_data[1][13] ));
 sky130_fd_sc_hd__dfxtp_1 _8179_ (.CLK(clknet_leaf_11_clk),
    .D(_0291_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.instr_data[1][14] ));
 sky130_fd_sc_hd__dfxtp_1 _8180_ (.CLK(clknet_leaf_11_clk),
    .D(_0292_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.instr_data[1][15] ));
 sky130_fd_sc_hd__dfxtp_2 _8181_ (.CLK(clknet_leaf_42_clk),
    .D(_0293_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[0] ));
 sky130_fd_sc_hd__dfxtp_2 _8182_ (.CLK(clknet_leaf_41_clk),
    .D(_0294_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[1] ));
 sky130_fd_sc_hd__dfxtp_2 _8183_ (.CLK(clknet_leaf_41_clk),
    .D(_0295_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[2] ));
 sky130_fd_sc_hd__dfxtp_2 _8184_ (.CLK(clknet_leaf_41_clk),
    .D(_0296_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[3] ));
 sky130_fd_sc_hd__dfxtp_2 _8185_ (.CLK(clknet_leaf_42_clk),
    .D(_0297_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[4] ));
 sky130_fd_sc_hd__dfxtp_2 _8186_ (.CLK(clknet_leaf_42_clk),
    .D(_0298_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[5] ));
 sky130_fd_sc_hd__dfxtp_2 _8187_ (.CLK(clknet_leaf_42_clk),
    .D(_0299_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[6] ));
 sky130_fd_sc_hd__dfxtp_1 _8188_ (.CLK(clknet_leaf_42_clk),
    .D(_0300_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[7] ));
 sky130_fd_sc_hd__dfxtp_2 _8189_ (.CLK(clknet_leaf_41_clk),
    .D(_0301_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[8] ));
 sky130_fd_sc_hd__dfxtp_2 _8190_ (.CLK(clknet_leaf_41_clk),
    .D(_0302_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[9] ));
 sky130_fd_sc_hd__dfxtp_2 _8191_ (.CLK(clknet_leaf_41_clk),
    .D(_0303_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[10] ));
 sky130_fd_sc_hd__dfxtp_2 _8192_ (.CLK(clknet_leaf_41_clk),
    .D(_0304_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[11] ));
 sky130_fd_sc_hd__dfxtp_2 _8193_ (.CLK(clknet_leaf_41_clk),
    .D(_0305_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[12] ));
 sky130_fd_sc_hd__dfxtp_2 _8194_ (.CLK(clknet_leaf_41_clk),
    .D(_0306_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[13] ));
 sky130_fd_sc_hd__dfxtp_2 _8195_ (.CLK(clknet_leaf_40_clk),
    .D(_0307_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[14] ));
 sky130_fd_sc_hd__dfxtp_1 _8196_ (.CLK(clknet_leaf_41_clk),
    .D(_0308_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[15] ));
 sky130_fd_sc_hd__dfxtp_1 _8197_ (.CLK(clknet_leaf_41_clk),
    .D(_0309_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[16] ));
 sky130_fd_sc_hd__dfxtp_1 _8198_ (.CLK(clknet_leaf_40_clk),
    .D(_0310_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[17] ));
 sky130_fd_sc_hd__dfxtp_1 _8199_ (.CLK(clknet_leaf_40_clk),
    .D(_0311_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[18] ));
 sky130_fd_sc_hd__dfxtp_1 _8200_ (.CLK(clknet_leaf_40_clk),
    .D(_0312_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[19] ));
 sky130_fd_sc_hd__dfxtp_1 _8201_ (.CLK(clknet_leaf_40_clk),
    .D(_0313_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[20] ));
 sky130_fd_sc_hd__dfxtp_1 _8202_ (.CLK(clknet_leaf_40_clk),
    .D(_0314_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[21] ));
 sky130_fd_sc_hd__dfxtp_1 _8203_ (.CLK(clknet_leaf_40_clk),
    .D(_0315_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[22] ));
 sky130_fd_sc_hd__dfxtp_1 _8204_ (.CLK(clknet_leaf_40_clk),
    .D(_0316_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[23] ));
 sky130_fd_sc_hd__dfxtp_1 _8205_ (.CLK(clknet_leaf_40_clk),
    .D(_0317_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[24] ));
 sky130_fd_sc_hd__dfxtp_1 _8206_ (.CLK(clknet_leaf_40_clk),
    .D(_0318_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[25] ));
 sky130_fd_sc_hd__dfxtp_1 _8207_ (.CLK(clknet_leaf_40_clk),
    .D(_0319_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[26] ));
 sky130_fd_sc_hd__dfxtp_1 _8208_ (.CLK(clknet_leaf_40_clk),
    .D(_0320_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[27] ));
 sky130_fd_sc_hd__dfxtp_2 _8209_ (.CLK(clknet_leaf_39_clk),
    .D(_0321_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[30] ));
 sky130_fd_sc_hd__dfxtp_2 _8210_ (.CLK(clknet_leaf_40_clk),
    .D(_0322_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[31] ));
 sky130_fd_sc_hd__dfxtp_1 _8211_ (.CLK(clknet_leaf_9_clk),
    .D(_0323_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.instr_data[0][0] ));
 sky130_fd_sc_hd__dfxtp_1 _8212_ (.CLK(clknet_leaf_13_clk),
    .D(_0324_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.instr_data[0][1] ));
 sky130_fd_sc_hd__dfxtp_2 _8213_ (.CLK(clknet_leaf_40_clk),
    .D(_0325_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_shift.adjusted_shift_amt[0] ));
 sky130_fd_sc_hd__dfxtp_2 _8214_ (.CLK(clknet_leaf_39_clk),
    .D(_0326_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_shift.adjusted_shift_amt[1] ));
 sky130_fd_sc_hd__dfxtp_1 _8215_ (.CLK(clknet_leaf_39_clk),
    .D(_0327_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_shift.b[2] ));
 sky130_fd_sc_hd__dfxtp_1 _8216_ (.CLK(clknet_leaf_39_clk),
    .D(_0328_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_shift.b[3] ));
 sky130_fd_sc_hd__dfxtp_1 _8217_ (.CLK(clknet_leaf_39_clk),
    .D(_0016_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.multiplier.accum[0] ));
 sky130_fd_sc_hd__dfxtp_1 _8218_ (.CLK(clknet_leaf_39_clk),
    .D(_0019_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.multiplier.accum[1] ));
 sky130_fd_sc_hd__dfxtp_1 _8219_ (.CLK(clknet_leaf_42_clk),
    .D(_0020_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.multiplier.accum[2] ));
 sky130_fd_sc_hd__dfxtp_1 _8220_ (.CLK(clknet_leaf_42_clk),
    .D(_0021_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.multiplier.accum[3] ));
 sky130_fd_sc_hd__dfxtp_1 _8221_ (.CLK(clknet_leaf_45_clk),
    .D(_0022_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.multiplier.accum[4] ));
 sky130_fd_sc_hd__dfxtp_1 _8222_ (.CLK(clknet_leaf_44_clk),
    .D(_0023_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.multiplier.accum[5] ));
 sky130_fd_sc_hd__dfxtp_1 _8223_ (.CLK(clknet_leaf_44_clk),
    .D(_0024_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.multiplier.accum[6] ));
 sky130_fd_sc_hd__dfxtp_1 _8224_ (.CLK(clknet_leaf_44_clk),
    .D(_0025_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.multiplier.accum[7] ));
 sky130_fd_sc_hd__dfxtp_1 _8225_ (.CLK(clknet_leaf_44_clk),
    .D(_0026_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.multiplier.accum[8] ));
 sky130_fd_sc_hd__dfxtp_1 _8226_ (.CLK(clknet_leaf_44_clk),
    .D(_0027_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.multiplier.accum[9] ));
 sky130_fd_sc_hd__dfxtp_1 _8227_ (.CLK(clknet_leaf_43_clk),
    .D(_0017_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.multiplier.accum[10] ));
 sky130_fd_sc_hd__dfxtp_1 _8228_ (.CLK(clknet_leaf_43_clk),
    .D(_0018_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.multiplier.accum[11] ));
 sky130_fd_sc_hd__dfxtp_1 _8229_ (.CLK(clknet_leaf_35_clk),
    .D(_0329_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.mepc[0] ));
 sky130_fd_sc_hd__dfxtp_1 _8230_ (.CLK(clknet_leaf_35_clk),
    .D(_0330_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.mepc[1] ));
 sky130_fd_sc_hd__dfxtp_2 _8231_ (.CLK(clknet_leaf_34_clk),
    .D(_0331_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.mepc[2] ));
 sky130_fd_sc_hd__dfxtp_1 _8232_ (.CLK(clknet_leaf_35_clk),
    .D(_0332_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.mepc[3] ));
 sky130_fd_sc_hd__dfxtp_1 _8233_ (.CLK(clknet_leaf_35_clk),
    .D(_0333_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.mepc[4] ));
 sky130_fd_sc_hd__dfxtp_1 _8234_ (.CLK(clknet_leaf_40_clk),
    .D(_0334_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.mepc[5] ));
 sky130_fd_sc_hd__dfxtp_1 _8235_ (.CLK(clknet_leaf_34_clk),
    .D(_0335_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.mepc[6] ));
 sky130_fd_sc_hd__dfxtp_1 _8236_ (.CLK(clknet_leaf_35_clk),
    .D(_0336_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.mepc[7] ));
 sky130_fd_sc_hd__dfxtp_1 _8237_ (.CLK(clknet_leaf_40_clk),
    .D(_0337_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.mepc[8] ));
 sky130_fd_sc_hd__dfxtp_1 _8238_ (.CLK(clknet_leaf_40_clk),
    .D(_0338_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.mepc[9] ));
 sky130_fd_sc_hd__dfxtp_1 _8239_ (.CLK(clknet_leaf_34_clk),
    .D(_0339_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.mepc[10] ));
 sky130_fd_sc_hd__dfxtp_1 _8240_ (.CLK(clknet_leaf_35_clk),
    .D(_0340_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.mepc[11] ));
 sky130_fd_sc_hd__dfxtp_1 _8241_ (.CLK(clknet_leaf_35_clk),
    .D(_0341_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.mepc[12] ));
 sky130_fd_sc_hd__dfxtp_1 _8242_ (.CLK(clknet_leaf_35_clk),
    .D(_0342_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.mepc[13] ));
 sky130_fd_sc_hd__dfxtp_1 _8243_ (.CLK(clknet_leaf_34_clk),
    .D(_0343_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.mepc[14] ));
 sky130_fd_sc_hd__dfxtp_1 _8244_ (.CLK(clknet_leaf_35_clk),
    .D(_0344_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.mepc[15] ));
 sky130_fd_sc_hd__dfxtp_1 _8245_ (.CLK(clknet_leaf_35_clk),
    .D(_0345_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.mepc[16] ));
 sky130_fd_sc_hd__dfxtp_1 _8246_ (.CLK(clknet_leaf_35_clk),
    .D(_0346_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.mepc[17] ));
 sky130_fd_sc_hd__dfxtp_1 _8247_ (.CLK(clknet_leaf_34_clk),
    .D(_0347_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.mepc[18] ));
 sky130_fd_sc_hd__dfxtp_1 _8248_ (.CLK(clknet_leaf_35_clk),
    .D(_0348_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.mepc[19] ));
 sky130_fd_sc_hd__dfxtp_2 _8249_ (.CLK(clknet_leaf_20_clk),
    .D(_0349_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.mem.instr_active ));
 sky130_fd_sc_hd__dfxtp_1 _8250_ (.CLK(clknet_leaf_22_clk),
    .D(_0350_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.load_top_bit ));
 sky130_fd_sc_hd__dfxtp_2 _8251_ (.CLK(clknet_leaf_19_clk),
    .D(_0351_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(debug_register_data));
 sky130_fd_sc_hd__dfxtp_1 _8252_ (.CLK(clknet_leaf_17_clk),
    .D(_0352_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.mem.data_stall ));
 sky130_fd_sc_hd__dfxtp_1 _8253_ (.CLK(clknet_leaf_17_clk),
    .D(_0082_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.mem.qspi_write_done ));
 sky130_fd_sc_hd__dfxtp_1 _8254_ (.CLK(clknet_leaf_43_clk),
    .D(_0353_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.multiplier.accum[12] ));
 sky130_fd_sc_hd__dfxtp_1 _8255_ (.CLK(clknet_leaf_43_clk),
    .D(_0354_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.multiplier.accum[13] ));
 sky130_fd_sc_hd__dfxtp_1 _8256_ (.CLK(clknet_leaf_43_clk),
    .D(_0355_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.multiplier.accum[14] ));
 sky130_fd_sc_hd__dfxtp_1 _8257_ (.CLK(clknet_leaf_42_clk),
    .D(_0356_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.multiplier.accum[15] ));
 sky130_fd_sc_hd__dfxtp_1 _8258_ (.CLK(clknet_leaf_17_clk),
    .D(_0357_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.mem.qspi_data_byte_idx[0] ));
 sky130_fd_sc_hd__dfxtp_4 _8259_ (.CLK(clknet_leaf_17_clk),
    .D(_0358_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.mem.qspi_data_byte_idx[1] ));
 sky130_fd_sc_hd__dfxtp_1 _8260_ (.CLK(clknet_leaf_13_clk),
    .D(_0359_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.instr_data_in[0] ));
 sky130_fd_sc_hd__dfxtp_1 _8261_ (.CLK(clknet_leaf_13_clk),
    .D(_0360_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.instr_data_in[1] ));
 sky130_fd_sc_hd__dfxtp_1 _8262_ (.CLK(clknet_leaf_14_clk),
    .D(_0361_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.instr_data_in[2] ));
 sky130_fd_sc_hd__dfxtp_2 _8263_ (.CLK(clknet_leaf_14_clk),
    .D(_0362_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.instr_data_in[3] ));
 sky130_fd_sc_hd__dfxtp_1 _8264_ (.CLK(clknet_leaf_14_clk),
    .D(_0363_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.instr_data_in[4] ));
 sky130_fd_sc_hd__dfxtp_2 _8265_ (.CLK(clknet_leaf_14_clk),
    .D(_0364_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.instr_data_in[5] ));
 sky130_fd_sc_hd__dfxtp_1 _8266_ (.CLK(clknet_leaf_14_clk),
    .D(_0365_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.instr_data_in[6] ));
 sky130_fd_sc_hd__dfxtp_2 _8267_ (.CLK(clknet_leaf_14_clk),
    .D(_0366_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.instr_data_in[7] ));
 sky130_fd_sc_hd__dfxtp_1 _8268_ (.CLK(clknet_leaf_14_clk),
    .D(_0367_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.mem.qspi_data_buf[8] ));
 sky130_fd_sc_hd__dfxtp_1 _8269_ (.CLK(clknet_leaf_14_clk),
    .D(_0368_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.mem.qspi_data_buf[9] ));
 sky130_fd_sc_hd__dfxtp_1 _8270_ (.CLK(clknet_leaf_14_clk),
    .D(_0369_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.mem.qspi_data_buf[10] ));
 sky130_fd_sc_hd__dfxtp_1 _8271_ (.CLK(clknet_leaf_21_clk),
    .D(_0370_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.mem.qspi_data_buf[11] ));
 sky130_fd_sc_hd__dfxtp_1 _8272_ (.CLK(clknet_leaf_14_clk),
    .D(_0371_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.mem.qspi_data_buf[12] ));
 sky130_fd_sc_hd__dfxtp_1 _8273_ (.CLK(clknet_leaf_14_clk),
    .D(_0372_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.mem.qspi_data_buf[13] ));
 sky130_fd_sc_hd__dfxtp_1 _8274_ (.CLK(clknet_leaf_14_clk),
    .D(_0373_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.mem.qspi_data_buf[14] ));
 sky130_fd_sc_hd__dfxtp_1 _8275_ (.CLK(clknet_leaf_17_clk),
    .D(_0374_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.mem.qspi_data_buf[15] ));
 sky130_fd_sc_hd__dfxtp_1 _8276_ (.CLK(clknet_leaf_13_clk),
    .D(_0375_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.mem.data_from_read[16] ));
 sky130_fd_sc_hd__dfxtp_1 _8277_ (.CLK(clknet_leaf_13_clk),
    .D(_0376_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.mem.data_from_read[17] ));
 sky130_fd_sc_hd__dfxtp_1 _8278_ (.CLK(clknet_leaf_17_clk),
    .D(_0377_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.mem.data_from_read[18] ));
 sky130_fd_sc_hd__dfxtp_1 _8279_ (.CLK(clknet_leaf_21_clk),
    .D(_0378_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.mem.data_from_read[19] ));
 sky130_fd_sc_hd__dfxtp_1 _8280_ (.CLK(clknet_leaf_13_clk),
    .D(_0379_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.mem.data_from_read[20] ));
 sky130_fd_sc_hd__dfxtp_1 _8281_ (.CLK(clknet_leaf_13_clk),
    .D(_0380_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.mem.data_from_read[21] ));
 sky130_fd_sc_hd__dfxtp_1 _8282_ (.CLK(clknet_leaf_13_clk),
    .D(_0381_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.mem.data_from_read[22] ));
 sky130_fd_sc_hd__dfxtp_1 _8283_ (.CLK(clknet_leaf_17_clk),
    .D(_0382_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.mem.data_from_read[23] ));
 sky130_fd_sc_hd__dfxtp_1 _8284_ (.CLK(clknet_leaf_14_clk),
    .D(_0383_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.mem.qspi_data_buf[24] ));
 sky130_fd_sc_hd__dfxtp_1 _8285_ (.CLK(clknet_leaf_14_clk),
    .D(_0384_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.mem.qspi_data_buf[25] ));
 sky130_fd_sc_hd__dfxtp_1 _8286_ (.CLK(clknet_leaf_14_clk),
    .D(_0385_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.mem.qspi_data_buf[26] ));
 sky130_fd_sc_hd__dfxtp_1 _8287_ (.CLK(clknet_leaf_17_clk),
    .D(_0386_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.mem.qspi_data_buf[27] ));
 sky130_fd_sc_hd__dfxtp_1 _8288_ (.CLK(clknet_leaf_14_clk),
    .D(_0387_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.mem.qspi_data_buf[28] ));
 sky130_fd_sc_hd__dfxtp_1 _8289_ (.CLK(clknet_leaf_14_clk),
    .D(_0388_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.mem.qspi_data_buf[29] ));
 sky130_fd_sc_hd__dfxtp_1 _8290_ (.CLK(clknet_leaf_14_clk),
    .D(_0389_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.mem.qspi_data_buf[30] ));
 sky130_fd_sc_hd__dfxtp_1 _8291_ (.CLK(clknet_leaf_16_clk),
    .D(_0390_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.mem.qspi_data_buf[31] ));
 sky130_fd_sc_hd__dfxtp_1 _8292_ (.CLK(clknet_leaf_20_clk),
    .D(_0391_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.instr_fetch_started ));
 sky130_fd_sc_hd__dfxtp_2 _8293_ (.CLK(clknet_leaf_15_clk),
    .D(_0392_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.mem.q_ctrl.read_cycles_count[0] ));
 sky130_fd_sc_hd__dfxtp_1 _8294_ (.CLK(clknet_leaf_15_clk),
    .D(_0393_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.mem.q_ctrl.read_cycles_count[1] ));
 sky130_fd_sc_hd__dfxtp_1 _8295_ (.CLK(clknet_leaf_15_clk),
    .D(_0394_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.mem.q_ctrl.read_cycles_count[2] ));
 sky130_fd_sc_hd__dfxtp_2 _8296_ (.CLK(clknet_leaf_16_clk),
    .D(_0395_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.mem.q_ctrl.data_req ));
 sky130_fd_sc_hd__dfxtp_1 _8297_ (.CLK(clknet_leaf_14_clk),
    .D(_0396_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.mem.q_ctrl.nibbles_remaining[0] ));
 sky130_fd_sc_hd__dfxtp_1 _8298_ (.CLK(clknet_leaf_14_clk),
    .D(_0397_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.mem.q_ctrl.nibbles_remaining[1] ));
 sky130_fd_sc_hd__dfxtp_1 _8299_ (.CLK(clknet_leaf_14_clk),
    .D(_0398_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.mem.q_ctrl.nibbles_remaining[2] ));
 sky130_fd_sc_hd__dfxtp_1 _8300_ (.CLK(clknet_leaf_16_clk),
    .D(_0399_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.mem.q_ctrl.is_writing ));
 sky130_fd_sc_hd__dfxtp_1 _8301_ (.CLK(clknet_leaf_15_clk),
    .D(_0400_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.mem.q_ctrl.fsm_state[0] ));
 sky130_fd_sc_hd__dfxtp_2 _8302_ (.CLK(clknet_leaf_15_clk),
    .D(_0401_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.mem.q_ctrl.fsm_state[1] ));
 sky130_fd_sc_hd__dfxtp_1 _8303_ (.CLK(clknet_leaf_15_clk),
    .D(_0402_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.mem.q_ctrl.fsm_state[2] ));
 sky130_fd_sc_hd__dfxtp_2 _8304_ (.CLK(clknet_leaf_16_clk),
    .D(_0403_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.mem.q_ctrl.data_ready ));
 sky130_fd_sc_hd__dfxtp_1 _8305_ (.CLK(clknet_leaf_16_clk),
    .D(_0404_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.mem.q_ctrl.spi_ram_b_select ));
 sky130_fd_sc_hd__dfxtp_1 _8306_ (.CLK(clknet_leaf_17_clk),
    .D(_0405_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.mem.q_ctrl.spi_ram_a_select ));
 sky130_fd_sc_hd__dfxtp_1 _8307_ (.CLK(clknet_leaf_16_clk),
    .D(_0406_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.mem.q_ctrl.spi_flash_select ));
 sky130_fd_sc_hd__dfxtp_2 _8308_ (.CLK(clknet_leaf_15_clk),
    .D(_0407_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.mem.q_ctrl.spi_clk_out ));
 sky130_fd_sc_hd__dfxtp_1 _8309_ (.CLK(clknet_leaf_15_clk),
    .D(_0408_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.mem.q_ctrl.spi_data_oe[0] ));
 sky130_fd_sc_hd__dfxtp_2 _8310_ (.CLK(clknet_leaf_39_clk),
    .D(_0409_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[28] ));
 sky130_fd_sc_hd__dfxtp_2 _8311_ (.CLK(clknet_leaf_39_clk),
    .D(_0410_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[29] ));
 sky130_fd_sc_hd__dfxtp_1 _8312_ (.CLK(clknet_leaf_16_clk),
    .D(_0411_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.mem.q_ctrl.spi_in_buffer[0] ));
 sky130_fd_sc_hd__dfxtp_1 _8313_ (.CLK(clknet_leaf_15_clk),
    .D(_0412_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.mem.q_ctrl.spi_in_buffer[1] ));
 sky130_fd_sc_hd__dfxtp_1 _8314_ (.CLK(clknet_leaf_16_clk),
    .D(_0413_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.mem.q_ctrl.spi_in_buffer[2] ));
 sky130_fd_sc_hd__dfxtp_1 _8315_ (.CLK(clknet_leaf_16_clk),
    .D(_0414_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.mem.q_ctrl.spi_in_buffer[3] ));
 sky130_fd_sc_hd__dfxtp_1 _8316_ (.CLK(clknet_leaf_18_clk),
    .D(_0415_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.mem.q_ctrl.spi_in_buffer[4] ));
 sky130_fd_sc_hd__dfxtp_1 _8317_ (.CLK(clknet_leaf_16_clk),
    .D(_0416_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.mem.q_ctrl.spi_in_buffer[5] ));
 sky130_fd_sc_hd__dfxtp_1 _8318_ (.CLK(clknet_leaf_16_clk),
    .D(_0417_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.mem.q_ctrl.spi_in_buffer[6] ));
 sky130_fd_sc_hd__dfxtp_1 _8319_ (.CLK(clknet_leaf_16_clk),
    .D(_0418_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.mem.q_ctrl.spi_in_buffer[7] ));
 sky130_fd_sc_hd__dfxtp_1 _8320_ (.CLK(clknet_leaf_16_clk),
    .D(_0419_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.instr_data_in[8] ));
 sky130_fd_sc_hd__dfxtp_1 _8321_ (.CLK(clknet_leaf_14_clk),
    .D(_0420_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.instr_data_in[9] ));
 sky130_fd_sc_hd__dfxtp_1 _8322_ (.CLK(clknet_leaf_13_clk),
    .D(_0421_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.instr_data_in[10] ));
 sky130_fd_sc_hd__dfxtp_1 _8323_ (.CLK(clknet_leaf_16_clk),
    .D(_0422_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.instr_data_in[11] ));
 sky130_fd_sc_hd__dfxtp_1 _8324_ (.CLK(clknet_leaf_13_clk),
    .D(_0423_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.instr_data_in[12] ));
 sky130_fd_sc_hd__dfxtp_1 _8325_ (.CLK(clknet_leaf_14_clk),
    .D(_0424_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.instr_data_in[13] ));
 sky130_fd_sc_hd__dfxtp_1 _8326_ (.CLK(clknet_leaf_13_clk),
    .D(_0425_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.instr_data_in[14] ));
 sky130_fd_sc_hd__dfxtp_1 _8327_ (.CLK(clknet_leaf_16_clk),
    .D(_0426_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.instr_data_in[15] ));
 sky130_fd_sc_hd__dfxtp_1 _8328_ (.CLK(clknet_leaf_17_clk),
    .D(_0427_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.mem.q_ctrl.last_ram_b_sel ));
 sky130_fd_sc_hd__dfxtp_1 _8329_ (.CLK(clknet_leaf_17_clk),
    .D(_0428_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.mem.q_ctrl.last_ram_a_sel ));
 sky130_fd_sc_hd__dfxtp_1 _8330_ (.CLK(clknet_leaf_17_clk),
    .D(_0429_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.instr_fetch_stopped ));
 sky130_fd_sc_hd__dfxtp_1 _8331_ (.CLK(clknet_leaf_13_clk),
    .D(_0430_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.instr_data[2][0] ));
 sky130_fd_sc_hd__dfxtp_1 _8332_ (.CLK(clknet_leaf_13_clk),
    .D(_0431_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.instr_data[2][1] ));
 sky130_fd_sc_hd__dfxtp_1 _8333_ (.CLK(clknet_leaf_18_clk),
    .D(_0432_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.mem.q_ctrl.delay_cycles_cfg[0] ));
 sky130_fd_sc_hd__dfxtp_1 _8334_ (.CLK(clknet_leaf_15_clk),
    .D(_0433_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.mem.q_ctrl.delay_cycles_cfg[1] ));
 sky130_fd_sc_hd__dfxtp_1 _8335_ (.CLK(clknet_leaf_16_clk),
    .D(_0434_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.mem.q_ctrl.delay_cycles_cfg[2] ));
 sky130_fd_sc_hd__dfxtp_1 _8336_ (.CLK(clknet_leaf_21_clk),
    .D(_0435_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.instr_write_offset[1] ));
 sky130_fd_sc_hd__dfxtp_2 _8337_ (.CLK(clknet_leaf_22_clk),
    .D(_0436_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.instr_write_offset[2] ));
 sky130_fd_sc_hd__dfxtp_1 _8338_ (.CLK(clknet_leaf_29_clk),
    .D(_0437_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.mem.q_ctrl.addr[0] ));
 sky130_fd_sc_hd__dfxtp_1 _8339_ (.CLK(clknet_leaf_33_clk),
    .D(_0438_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.mem.q_ctrl.addr[1] ));
 sky130_fd_sc_hd__dfxtp_1 _8340_ (.CLK(clknet_leaf_33_clk),
    .D(_0439_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.mem.q_ctrl.addr[2] ));
 sky130_fd_sc_hd__dfxtp_1 _8341_ (.CLK(clknet_leaf_29_clk),
    .D(_0440_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.mem.q_ctrl.addr[3] ));
 sky130_fd_sc_hd__dfxtp_1 _8342_ (.CLK(clknet_leaf_22_clk),
    .D(_0441_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.pc[1] ));
 sky130_fd_sc_hd__dfxtp_2 _8343_ (.CLK(clknet_leaf_22_clk),
    .D(_0442_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.pc[2] ));
 sky130_fd_sc_hd__dfxtp_1 _8344_ (.CLK(clknet_leaf_26_clk),
    .D(_0443_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_spi.end_txn_reg ));
 sky130_fd_sc_hd__dfxtp_1 _8345_ (.CLK(clknet_leaf_24_clk),
    .D(_0444_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.instr_data_start[3] ));
 sky130_fd_sc_hd__dfxtp_2 _8346_ (.CLK(clknet_leaf_24_clk),
    .D(_0445_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.instr_data_start[4] ));
 sky130_fd_sc_hd__dfxtp_2 _8347_ (.CLK(clknet_leaf_24_clk),
    .D(_0446_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.instr_data_start[5] ));
 sky130_fd_sc_hd__dfxtp_1 _8348_ (.CLK(clknet_leaf_24_clk),
    .D(_0447_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.instr_data_start[6] ));
 sky130_fd_sc_hd__dfxtp_2 _8349_ (.CLK(clknet_leaf_36_clk),
    .D(_0448_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.instr_data_start[7] ));
 sky130_fd_sc_hd__dfxtp_2 _8350_ (.CLK(clknet_leaf_33_clk),
    .D(_0449_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.instr_data_start[8] ));
 sky130_fd_sc_hd__dfxtp_1 _8351_ (.CLK(clknet_leaf_25_clk),
    .D(_0450_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.instr_data_start[9] ));
 sky130_fd_sc_hd__dfxtp_2 _8352_ (.CLK(clknet_leaf_25_clk),
    .D(_0451_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.instr_data_start[10] ));
 sky130_fd_sc_hd__dfxtp_2 _8353_ (.CLK(clknet_leaf_33_clk),
    .D(_0452_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.instr_data_start[11] ));
 sky130_fd_sc_hd__dfxtp_1 _8354_ (.CLK(clknet_leaf_36_clk),
    .D(_0453_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.instr_data_start[12] ));
 sky130_fd_sc_hd__dfxtp_2 _8355_ (.CLK(clknet_leaf_36_clk),
    .D(_0454_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.instr_data_start[13] ));
 sky130_fd_sc_hd__dfxtp_2 _8356_ (.CLK(clknet_leaf_36_clk),
    .D(_0455_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.instr_data_start[14] ));
 sky130_fd_sc_hd__dfxtp_1 _8357_ (.CLK(clknet_leaf_36_clk),
    .D(_0456_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.instr_data_start[15] ));
 sky130_fd_sc_hd__dfxtp_2 _8358_ (.CLK(clknet_leaf_36_clk),
    .D(_0457_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.instr_data_start[16] ));
 sky130_fd_sc_hd__dfxtp_2 _8359_ (.CLK(clknet_leaf_36_clk),
    .D(_0458_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.instr_data_start[17] ));
 sky130_fd_sc_hd__dfxtp_1 _8360_ (.CLK(clknet_leaf_36_clk),
    .D(_0459_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.instr_data_start[18] ));
 sky130_fd_sc_hd__dfxtp_2 _8361_ (.CLK(clknet_leaf_36_clk),
    .D(_0460_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.instr_data_start[19] ));
 sky130_fd_sc_hd__dfxtp_2 _8362_ (.CLK(clknet_leaf_36_clk),
    .D(_0461_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.instr_data_start[20] ));
 sky130_fd_sc_hd__dfxtp_2 _8363_ (.CLK(clknet_leaf_36_clk),
    .D(_0462_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.instr_data_start[21] ));
 sky130_fd_sc_hd__dfxtp_2 _8364_ (.CLK(clknet_leaf_36_clk),
    .D(_0463_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.instr_data_start[22] ));
 sky130_fd_sc_hd__dfxtp_2 _8365_ (.CLK(clknet_leaf_36_clk),
    .D(_0464_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.instr_data_start[23] ));
 sky130_fd_sc_hd__dfxtp_1 _8366_ (.CLK(clknet_leaf_22_clk),
    .D(_0465_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.instr_fetch_running ));
 sky130_fd_sc_hd__dfxtp_2 _8367_ (.CLK(clknet_leaf_24_clk),
    .D(_0466_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.was_early_branch ));
 sky130_fd_sc_hd__dfxtp_2 _8368_ (.CLK(clknet_leaf_21_clk),
    .D(_0467_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.data_write_n[0] ));
 sky130_fd_sc_hd__dfxtp_2 _8369_ (.CLK(clknet_leaf_21_clk),
    .D(_0468_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.data_write_n[1] ));
 sky130_fd_sc_hd__dfxtp_2 _8370_ (.CLK(clknet_leaf_21_clk),
    .D(_0469_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.data_read_n[0] ));
 sky130_fd_sc_hd__dfxtp_1 _8371_ (.CLK(clknet_leaf_20_clk),
    .D(_0470_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.data_read_n[1] ));
 sky130_fd_sc_hd__dfxtp_1 _8372_ (.CLK(clknet_leaf_21_clk),
    .D(_0028_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.data_continue ));
 sky130_fd_sc_hd__dfxtp_2 _8373_ (.CLK(clknet_leaf_22_clk),
    .D(_0471_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.no_write_in_progress ));
 sky130_fd_sc_hd__dfxtp_1 _8374_ (.CLK(clknet_leaf_21_clk),
    .D(_0472_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.load_started ));
 sky130_fd_sc_hd__dfxtp_2 _8375_ (.CLK(clknet_leaf_25_clk),
    .D(_0473_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_debug_uart_tx.uart_tx_data[0] ));
 sky130_fd_sc_hd__dfxtp_1 _8376_ (.CLK(clknet_leaf_25_clk),
    .D(_0474_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_debug_uart_tx.uart_tx_data[1] ));
 sky130_fd_sc_hd__dfxtp_1 _8377_ (.CLK(clknet_leaf_25_clk),
    .D(_0475_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_debug_uart_tx.uart_tx_data[2] ));
 sky130_fd_sc_hd__dfxtp_2 _8378_ (.CLK(clknet_leaf_26_clk),
    .D(_0476_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_debug_uart_tx.uart_tx_data[3] ));
 sky130_fd_sc_hd__dfxtp_2 _8379_ (.CLK(clknet_leaf_19_clk),
    .D(_0477_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_debug_uart_tx.uart_tx_data[4] ));
 sky130_fd_sc_hd__dfxtp_2 _8380_ (.CLK(clknet_leaf_19_clk),
    .D(_0478_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_debug_uart_tx.uart_tx_data[5] ));
 sky130_fd_sc_hd__dfxtp_1 _8381_ (.CLK(clknet_leaf_19_clk),
    .D(_0479_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_debug_uart_tx.uart_tx_data[6] ));
 sky130_fd_sc_hd__dfxtp_2 _8382_ (.CLK(clknet_leaf_19_clk),
    .D(_0480_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_debug_uart_tx.uart_tx_data[7] ));
 sky130_fd_sc_hd__dfxtp_1 _8383_ (.CLK(clknet_leaf_26_clk),
    .D(_0481_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_spi.end_txn ));
 sky130_fd_sc_hd__dfxtp_1 _8384_ (.CLK(clknet_leaf_26_clk),
    .D(_0482_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_spi.dc_in ));
 sky130_fd_sc_hd__dfxtp_1 _8385_ (.CLK(clknet_leaf_26_clk),
    .D(_0483_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.data_out[10] ));
 sky130_fd_sc_hd__dfxtp_1 _8386_ (.CLK(clknet_leaf_26_clk),
    .D(_0484_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.data_out[11] ));
 sky130_fd_sc_hd__dfxtp_1 _8387_ (.CLK(clknet_leaf_19_clk),
    .D(_0485_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.data_out[12] ));
 sky130_fd_sc_hd__dfxtp_1 _8388_ (.CLK(clknet_leaf_19_clk),
    .D(_0486_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.data_out[13] ));
 sky130_fd_sc_hd__dfxtp_1 _8389_ (.CLK(clknet_leaf_19_clk),
    .D(_0487_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.data_out[14] ));
 sky130_fd_sc_hd__dfxtp_1 _8390_ (.CLK(clknet_leaf_20_clk),
    .D(_0488_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.data_out[15] ));
 sky130_fd_sc_hd__dfxtp_1 _8391_ (.CLK(clknet_leaf_26_clk),
    .D(_0489_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.data_out[16] ));
 sky130_fd_sc_hd__dfxtp_1 _8392_ (.CLK(clknet_leaf_26_clk),
    .D(_0490_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.data_out[17] ));
 sky130_fd_sc_hd__dfxtp_1 _8393_ (.CLK(clknet_leaf_26_clk),
    .D(_0491_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.data_out[18] ));
 sky130_fd_sc_hd__dfxtp_1 _8394_ (.CLK(clknet_leaf_26_clk),
    .D(_0492_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.data_out[19] ));
 sky130_fd_sc_hd__dfxtp_1 _8395_ (.CLK(clknet_leaf_19_clk),
    .D(_0493_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.data_out[20] ));
 sky130_fd_sc_hd__dfxtp_1 _8396_ (.CLK(clknet_leaf_20_clk),
    .D(_0494_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.data_out[21] ));
 sky130_fd_sc_hd__dfxtp_1 _8397_ (.CLK(clknet_leaf_20_clk),
    .D(_0495_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.data_out[22] ));
 sky130_fd_sc_hd__dfxtp_1 _8398_ (.CLK(clknet_leaf_20_clk),
    .D(_0496_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.data_out[23] ));
 sky130_fd_sc_hd__dfxtp_1 _8399_ (.CLK(clknet_leaf_20_clk),
    .D(_0497_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.data_out[24] ));
 sky130_fd_sc_hd__dfxtp_1 _8400_ (.CLK(clknet_leaf_26_clk),
    .D(_0498_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.data_out[25] ));
 sky130_fd_sc_hd__dfxtp_1 _8401_ (.CLK(clknet_leaf_19_clk),
    .D(_0499_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.data_out[26] ));
 sky130_fd_sc_hd__dfxtp_1 _8402_ (.CLK(clknet_leaf_26_clk),
    .D(_0500_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.data_out[27] ));
 sky130_fd_sc_hd__dfxtp_1 _8403_ (.CLK(clknet_leaf_20_clk),
    .D(_0501_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.data_out[28] ));
 sky130_fd_sc_hd__dfxtp_1 _8404_ (.CLK(clknet_leaf_20_clk),
    .D(_0502_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.data_out[29] ));
 sky130_fd_sc_hd__dfxtp_1 _8405_ (.CLK(clknet_leaf_20_clk),
    .D(_0503_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.data_out[30] ));
 sky130_fd_sc_hd__dfxtp_1 _8406_ (.CLK(clknet_leaf_20_clk),
    .D(_0504_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.data_out[31] ));
 sky130_fd_sc_hd__dfxtp_2 _8407_ (.CLK(clknet_leaf_22_clk),
    .D(_0505_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.counter[2] ));
 sky130_fd_sc_hd__dfxtp_1 _8408_ (.CLK(clknet_leaf_24_clk),
    .D(_0506_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.counter[3] ));
 sky130_fd_sc_hd__dfxtp_4 _8409_ (.CLK(clknet_leaf_22_clk),
    .D(_0507_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.counter[4] ));
 sky130_fd_sc_hd__dfxtp_1 _8410_ (.CLK(clknet_leaf_7_clk),
    .D(_0508_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.data_ready_core ));
 sky130_fd_sc_hd__dfxtp_1 _8411_ (.CLK(clknet_leaf_22_clk),
    .D(_0509_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.data_ready_latch ));
 sky130_fd_sc_hd__dfxtp_1 _8412_ (.CLK(clknet_leaf_7_clk),
    .D(_0510_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.is_load ));
 sky130_fd_sc_hd__dfxtp_1 _8413_ (.CLK(clknet_leaf_6_clk),
    .D(_0511_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.is_alu_imm ));
 sky130_fd_sc_hd__dfxtp_1 _8414_ (.CLK(clknet_leaf_6_clk),
    .D(_0512_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.is_auipc ));
 sky130_fd_sc_hd__dfxtp_2 _8415_ (.CLK(clknet_leaf_7_clk),
    .D(_0513_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.is_store ));
 sky130_fd_sc_hd__dfxtp_1 _8416_ (.CLK(clknet_leaf_6_clk),
    .D(_0514_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.is_alu_reg ));
 sky130_fd_sc_hd__dfxtp_1 _8417_ (.CLK(clknet_leaf_7_clk),
    .D(_0515_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.is_lui ));
 sky130_fd_sc_hd__dfxtp_2 _8418_ (.CLK(clknet_leaf_6_clk),
    .D(_0516_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.is_branch ));
 sky130_fd_sc_hd__dfxtp_1 _8419_ (.CLK(clknet_leaf_7_clk),
    .D(_0517_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.is_jalr ));
 sky130_fd_sc_hd__dfxtp_2 _8420_ (.CLK(clknet_leaf_7_clk),
    .D(_0518_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.is_jal ));
 sky130_fd_sc_hd__dfxtp_1 _8421_ (.CLK(clknet_leaf_7_clk),
    .D(_0519_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.is_system ));
 sky130_fd_sc_hd__dfxtp_1 _8422_ (.CLK(clknet_leaf_23_clk),
    .D(_0520_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.imm_lo[0] ));
 sky130_fd_sc_hd__dfxtp_2 _8423_ (.CLK(clknet_leaf_7_clk),
    .D(_0521_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.imm_lo[1] ));
 sky130_fd_sc_hd__dfxtp_2 _8424_ (.CLK(clknet_leaf_9_clk),
    .D(_0522_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.imm_lo[2] ));
 sky130_fd_sc_hd__dfxtp_2 _8425_ (.CLK(clknet_leaf_23_clk),
    .D(_0523_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.imm_lo[3] ));
 sky130_fd_sc_hd__dfxtp_2 _8426_ (.CLK(clknet_leaf_9_clk),
    .D(_0524_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.imm_lo[4] ));
 sky130_fd_sc_hd__dfxtp_2 _8427_ (.CLK(clknet_leaf_9_clk),
    .D(_0525_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.imm_lo[5] ));
 sky130_fd_sc_hd__dfxtp_2 _8428_ (.CLK(clknet_leaf_9_clk),
    .D(_0526_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.imm_lo[6] ));
 sky130_fd_sc_hd__dfxtp_2 _8429_ (.CLK(clknet_leaf_22_clk),
    .D(_0527_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.imm_lo[7] ));
 sky130_fd_sc_hd__dfxtp_2 _8430_ (.CLK(clknet_leaf_23_clk),
    .D(_0528_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.imm_lo[8] ));
 sky130_fd_sc_hd__dfxtp_4 _8431_ (.CLK(clknet_leaf_8_clk),
    .D(_0529_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.imm_lo[9] ));
 sky130_fd_sc_hd__dfxtp_2 _8432_ (.CLK(clknet_leaf_8_clk),
    .D(_0530_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.imm_lo[10] ));
 sky130_fd_sc_hd__dfxtp_2 _8433_ (.CLK(clknet_leaf_22_clk),
    .D(_0531_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.imm_lo[11] ));
 sky130_fd_sc_hd__dfxtp_2 _8434_ (.CLK(clknet_leaf_8_clk),
    .D(_0532_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.imm[12] ));
 sky130_fd_sc_hd__dfxtp_2 _8435_ (.CLK(clknet_leaf_8_clk),
    .D(_0533_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.imm[13] ));
 sky130_fd_sc_hd__dfxtp_2 _8436_ (.CLK(clknet_leaf_21_clk),
    .D(_0534_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.imm[14] ));
 sky130_fd_sc_hd__dfxtp_2 _8437_ (.CLK(clknet_leaf_8_clk),
    .D(_0535_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.imm[15] ));
 sky130_fd_sc_hd__dfxtp_2 _8438_ (.CLK(clknet_leaf_8_clk),
    .D(_0536_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.imm[16] ));
 sky130_fd_sc_hd__dfxtp_2 _8439_ (.CLK(clknet_leaf_22_clk),
    .D(_0537_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.imm[17] ));
 sky130_fd_sc_hd__dfxtp_2 _8440_ (.CLK(clknet_leaf_22_clk),
    .D(_0538_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.imm[18] ));
 sky130_fd_sc_hd__dfxtp_2 _8441_ (.CLK(clknet_leaf_21_clk),
    .D(_0539_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.imm[19] ));
 sky130_fd_sc_hd__dfxtp_2 _8442_ (.CLK(clknet_leaf_7_clk),
    .D(_0540_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.imm[20] ));
 sky130_fd_sc_hd__dfxtp_2 _8443_ (.CLK(clknet_leaf_7_clk),
    .D(_0541_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.imm[21] ));
 sky130_fd_sc_hd__dfxtp_1 _8444_ (.CLK(clknet_leaf_22_clk),
    .D(_0542_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.imm[22] ));
 sky130_fd_sc_hd__dfxtp_2 _8445_ (.CLK(clknet_leaf_7_clk),
    .D(_0543_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.imm[23] ));
 sky130_fd_sc_hd__dfxtp_1 _8446_ (.CLK(clknet_leaf_8_clk),
    .D(_0544_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.imm[24] ));
 sky130_fd_sc_hd__dfxtp_1 _8447_ (.CLK(clknet_leaf_9_clk),
    .D(_0545_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.imm[25] ));
 sky130_fd_sc_hd__dfxtp_1 _8448_ (.CLK(clknet_leaf_7_clk),
    .D(_0546_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.imm[26] ));
 sky130_fd_sc_hd__dfxtp_1 _8449_ (.CLK(clknet_leaf_8_clk),
    .D(_0547_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.imm[27] ));
 sky130_fd_sc_hd__dfxtp_1 _8450_ (.CLK(clknet_leaf_9_clk),
    .D(_0548_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.imm[28] ));
 sky130_fd_sc_hd__dfxtp_1 _8451_ (.CLK(clknet_leaf_22_clk),
    .D(_0549_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.imm[29] ));
 sky130_fd_sc_hd__dfxtp_1 _8452_ (.CLK(clknet_leaf_22_clk),
    .D(_0550_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.imm[30] ));
 sky130_fd_sc_hd__dfxtp_1 _8453_ (.CLK(clknet_leaf_22_clk),
    .D(_0551_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.imm[31] ));
 sky130_fd_sc_hd__dfxtp_2 _8454_ (.CLK(clknet_leaf_6_clk),
    .D(_0552_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.alu_op[0] ));
 sky130_fd_sc_hd__dfxtp_1 _8455_ (.CLK(clknet_leaf_38_clk),
    .D(_0553_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.alu_op[1] ));
 sky130_fd_sc_hd__dfxtp_1 _8456_ (.CLK(clknet_leaf_39_clk),
    .D(_0554_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.alu_op[2] ));
 sky130_fd_sc_hd__dfxtp_4 _8457_ (.CLK(clknet_leaf_6_clk),
    .D(_0555_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.alu_op[3] ));
 sky130_fd_sc_hd__dfxtp_4 _8458_ (.CLK(clknet_leaf_6_clk),
    .D(_0556_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.mem_op[0] ));
 sky130_fd_sc_hd__dfxtp_1 _8459_ (.CLK(clknet_leaf_8_clk),
    .D(_0557_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.mem_op[1] ));
 sky130_fd_sc_hd__dfxtp_1 _8460_ (.CLK(clknet_leaf_7_clk),
    .D(_0558_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.mem_op[2] ));
 sky130_fd_sc_hd__dfxtp_2 _8461_ (.CLK(clknet_leaf_51_clk),
    .D(_0559_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.rs1[0] ));
 sky130_fd_sc_hd__dfxtp_2 _8462_ (.CLK(clknet_leaf_51_clk),
    .D(_0560_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.rs1[1] ));
 sky130_fd_sc_hd__dfxtp_2 _8463_ (.CLK(clknet_leaf_51_clk),
    .D(_0561_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.rs1[2] ));
 sky130_fd_sc_hd__dfxtp_2 _8464_ (.CLK(clknet_leaf_51_clk),
    .D(_0562_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.rs1[3] ));
 sky130_fd_sc_hd__dfxtp_2 _8465_ (.CLK(clknet_leaf_52_clk),
    .D(_0563_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.rs2[0] ));
 sky130_fd_sc_hd__dfxtp_2 _8466_ (.CLK(clknet_leaf_5_clk),
    .D(_0564_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.rs2[1] ));
 sky130_fd_sc_hd__dfxtp_2 _8467_ (.CLK(clknet_leaf_52_clk),
    .D(_0565_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.rs2[2] ));
 sky130_fd_sc_hd__dfxtp_2 _8468_ (.CLK(clknet_leaf_52_clk),
    .D(_0566_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_registers.rs2[3] ));
 sky130_fd_sc_hd__dfxtp_1 _8469_ (.CLK(clknet_leaf_7_clk),
    .D(_0567_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.instr_len[1] ));
 sky130_fd_sc_hd__dfxtp_1 _8470_ (.CLK(clknet_leaf_7_clk),
    .D(_0568_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.instr_len[2] ));
 sky130_fd_sc_hd__dfxtp_1 _8471_ (.CLK(clknet_leaf_6_clk),
    .D(_0569_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.additional_mem_ops[0] ));
 sky130_fd_sc_hd__dfxtp_1 _8472_ (.CLK(clknet_leaf_6_clk),
    .D(_0570_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.additional_mem_ops[1] ));
 sky130_fd_sc_hd__dfxtp_1 _8473_ (.CLK(clknet_leaf_6_clk),
    .D(_0571_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.additional_mem_ops[2] ));
 sky130_fd_sc_hd__dfxtp_1 _8474_ (.CLK(clknet_leaf_6_clk),
    .D(_0572_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.mem_op_increment_reg ));
 sky130_fd_sc_hd__dfxtp_2 _8475_ (.CLK(clknet_leaf_7_clk),
    .D(_0573_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.is_interrupt ));
 sky130_fd_sc_hd__dfxtp_4 _8476_ (.CLK(clknet_leaf_23_clk),
    .D(_0574_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.debug_instr_valid ));
 sky130_fd_sc_hd__dfxtp_2 _8477_ (.CLK(clknet_leaf_22_clk),
    .D(_0575_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.instr_write_offset[3] ));
 sky130_fd_sc_hd__dfxtp_1 _8478_ (.CLK(clknet_leaf_29_clk),
    .D(_0576_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.mem.q_ctrl.addr[4] ));
 sky130_fd_sc_hd__dfxtp_1 _8479_ (.CLK(clknet_leaf_32_clk),
    .D(_0577_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.mem.q_ctrl.addr[5] ));
 sky130_fd_sc_hd__dfxtp_1 _8480_ (.CLK(clknet_leaf_33_clk),
    .D(_0578_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.mem.q_ctrl.addr[6] ));
 sky130_fd_sc_hd__dfxtp_1 _8481_ (.CLK(clknet_leaf_32_clk),
    .D(_0579_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.mem.q_ctrl.addr[7] ));
 sky130_fd_sc_hd__dfxtp_1 _8482_ (.CLK(clknet_leaf_33_clk),
    .D(_0580_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.mem.q_ctrl.addr[8] ));
 sky130_fd_sc_hd__dfxtp_1 _8483_ (.CLK(clknet_leaf_32_clk),
    .D(_0581_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.mem.q_ctrl.addr[9] ));
 sky130_fd_sc_hd__dfxtp_1 _8484_ (.CLK(clknet_leaf_32_clk),
    .D(_0582_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.mem.q_ctrl.addr[10] ));
 sky130_fd_sc_hd__dfxtp_1 _8485_ (.CLK(clknet_leaf_32_clk),
    .D(_0583_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.mem.q_ctrl.addr[11] ));
 sky130_fd_sc_hd__dfxtp_1 _8486_ (.CLK(clknet_leaf_33_clk),
    .D(_0584_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.mem.q_ctrl.addr[12] ));
 sky130_fd_sc_hd__dfxtp_1 _8487_ (.CLK(clknet_leaf_32_clk),
    .D(_0585_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.mem.q_ctrl.addr[13] ));
 sky130_fd_sc_hd__dfxtp_1 _8488_ (.CLK(clknet_leaf_32_clk),
    .D(_0586_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.mem.q_ctrl.addr[14] ));
 sky130_fd_sc_hd__dfxtp_1 _8489_ (.CLK(clknet_leaf_32_clk),
    .D(_0587_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.mem.q_ctrl.addr[15] ));
 sky130_fd_sc_hd__dfxtp_1 _8490_ (.CLK(clknet_leaf_32_clk),
    .D(_0588_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.mem.q_ctrl.addr[16] ));
 sky130_fd_sc_hd__dfxtp_1 _8491_ (.CLK(clknet_leaf_32_clk),
    .D(_0589_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.mem.q_ctrl.addr[17] ));
 sky130_fd_sc_hd__dfxtp_1 _8492_ (.CLK(clknet_leaf_32_clk),
    .D(_0590_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.mem.q_ctrl.addr[18] ));
 sky130_fd_sc_hd__dfxtp_1 _8493_ (.CLK(clknet_leaf_32_clk),
    .D(_0591_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.mem.q_ctrl.addr[19] ));
 sky130_fd_sc_hd__dfxtp_2 _8494_ (.CLK(clknet_leaf_32_clk),
    .D(_0592_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.mem.q_ctrl.addr[20] ));
 sky130_fd_sc_hd__dfxtp_2 _8495_ (.CLK(clknet_leaf_32_clk),
    .D(_0593_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.mem.q_ctrl.addr[21] ));
 sky130_fd_sc_hd__dfxtp_2 _8496_ (.CLK(clknet_leaf_32_clk),
    .D(_0594_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.mem.q_ctrl.addr[22] ));
 sky130_fd_sc_hd__dfxtp_2 _8497_ (.CLK(clknet_leaf_29_clk),
    .D(_0595_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.mem.q_ctrl.addr[23] ));
 sky130_fd_sc_hd__dfxtp_1 _8498_ (.CLK(clknet_leaf_39_clk),
    .D(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.data[0] ));
 sky130_fd_sc_hd__dfxtp_1 _8499_ (.CLK(clknet_leaf_45_clk),
    .D(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.data[1] ));
 sky130_fd_sc_hd__dfxtp_1 _8500_ (.CLK(clknet_leaf_49_clk),
    .D(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.data[2] ));
 sky130_fd_sc_hd__dfxtp_1 _8501_ (.CLK(clknet_leaf_44_clk),
    .D(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.data[3] ));
 sky130_fd_sc_hd__dfxtp_1 _8502_ (.CLK(clknet_leaf_49_clk),
    .D(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.register[8] ));
 sky130_fd_sc_hd__dfxtp_1 _8503_ (.CLK(clknet_leaf_45_clk),
    .D(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.register[9] ));
 sky130_fd_sc_hd__dfxtp_1 _8504_ (.CLK(clknet_leaf_49_clk),
    .D(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.register[10] ));
 sky130_fd_sc_hd__dfxtp_1 _8505_ (.CLK(clknet_leaf_45_clk),
    .D(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.register[11] ));
 sky130_fd_sc_hd__dfxtp_1 _8506_ (.CLK(clknet_leaf_49_clk),
    .D(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.register[12] ));
 sky130_fd_sc_hd__dfxtp_1 _8507_ (.CLK(clknet_leaf_45_clk),
    .D(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.register[13] ));
 sky130_fd_sc_hd__dfxtp_1 _8508_ (.CLK(clknet_leaf_49_clk),
    .D(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.register[14] ));
 sky130_fd_sc_hd__dfxtp_1 _8509_ (.CLK(clknet_leaf_45_clk),
    .D(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.register[15] ));
 sky130_fd_sc_hd__dfxtp_1 _8510_ (.CLK(clknet_leaf_49_clk),
    .D(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.register[16] ));
 sky130_fd_sc_hd__dfxtp_1 _8511_ (.CLK(clknet_leaf_45_clk),
    .D(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.register[17] ));
 sky130_fd_sc_hd__dfxtp_1 _8512_ (.CLK(clknet_leaf_49_clk),
    .D(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.register[18] ));
 sky130_fd_sc_hd__dfxtp_1 _8513_ (.CLK(clknet_leaf_45_clk),
    .D(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.register[19] ));
 sky130_fd_sc_hd__dfxtp_1 _8514_ (.CLK(clknet_leaf_49_clk),
    .D(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.register[20] ));
 sky130_fd_sc_hd__dfxtp_1 _8515_ (.CLK(clknet_leaf_45_clk),
    .D(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.register[21] ));
 sky130_fd_sc_hd__dfxtp_1 _8516_ (.CLK(clknet_leaf_48_clk),
    .D(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.register[22] ));
 sky130_fd_sc_hd__dfxtp_1 _8517_ (.CLK(clknet_leaf_46_clk),
    .D(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.register[23] ));
 sky130_fd_sc_hd__dfxtp_1 _8518_ (.CLK(clknet_leaf_50_clk),
    .D(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.register[24] ));
 sky130_fd_sc_hd__dfxtp_1 _8519_ (.CLK(clknet_leaf_48_clk),
    .D(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.register[25] ));
 sky130_fd_sc_hd__dfxtp_1 _8520_ (.CLK(clknet_leaf_50_clk),
    .D(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.register[26] ));
 sky130_fd_sc_hd__dfxtp_1 _8521_ (.CLK(clknet_leaf_46_clk),
    .D(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.register[27] ));
 sky130_fd_sc_hd__dfxtp_1 _8522_ (.CLK(clknet_leaf_49_clk),
    .D(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.register[28] ));
 sky130_fd_sc_hd__dfxtp_1 _8523_ (.CLK(clknet_leaf_48_clk),
    .D(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.register[29] ));
 sky130_fd_sc_hd__dfxtp_1 _8524_ (.CLK(clknet_leaf_50_clk),
    .D(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.register[30] ));
 sky130_fd_sc_hd__dfxtp_1 _8525_ (.CLK(clknet_leaf_47_clk),
    .D(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.register[31] ));
 sky130_fd_sc_hd__dfxtp_1 _8526_ (.CLK(clknet_leaf_6_clk),
    .D(_0596_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.register[0] ));
 sky130_fd_sc_hd__dfxtp_1 _8527_ (.CLK(clknet_leaf_3_clk),
    .D(_0597_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.register[1] ));
 sky130_fd_sc_hd__dfxtp_1 _8528_ (.CLK(clknet_leaf_4_clk),
    .D(_0598_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.register[2] ));
 sky130_fd_sc_hd__dfxtp_1 _8529_ (.CLK(clknet_leaf_51_clk),
    .D(_0599_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.register[3] ));
 sky130_fd_sc_hd__dfxtp_1 _8530_ (.CLK(clknet_leaf_50_clk),
    .D(_0600_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.cy ));
 sky130_fd_sc_hd__dfxtp_1 _8531_ (.CLK(clknet_leaf_50_clk),
    .D(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.cycle_count[0] ));
 sky130_fd_sc_hd__dfxtp_1 _8532_ (.CLK(clknet_leaf_6_clk),
    .D(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.cycle_count[1] ));
 sky130_fd_sc_hd__dfxtp_1 _8533_ (.CLK(clknet_leaf_51_clk),
    .D(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.cycle_count[2] ));
 sky130_fd_sc_hd__dfxtp_1 _8534_ (.CLK(clknet_leaf_50_clk),
    .D(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.cycle_count[3] ));
 sky130_fd_sc_hd__dfxtp_1 _8535_ (.CLK(clknet_leaf_50_clk),
    .D(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.cycle_count_wide[4] ));
 sky130_fd_sc_hd__dfxtp_1 _8536_ (.CLK(clknet_leaf_6_clk),
    .D(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.cycle_count_wide[5] ));
 sky130_fd_sc_hd__dfxtp_1 _8537_ (.CLK(clknet_leaf_5_clk),
    .D(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.cycle_count_wide[6] ));
 sky130_fd_sc_hd__dfxtp_1 _8538_ (.CLK(clknet_leaf_50_clk),
    .D(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.register[11] ));
 sky130_fd_sc_hd__dfxtp_1 _8539_ (.CLK(clknet_leaf_51_clk),
    .D(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.register[12] ));
 sky130_fd_sc_hd__dfxtp_1 _8540_ (.CLK(clknet_leaf_4_clk),
    .D(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.register[13] ));
 sky130_fd_sc_hd__dfxtp_1 _8541_ (.CLK(clknet_leaf_5_clk),
    .D(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.register[14] ));
 sky130_fd_sc_hd__dfxtp_1 _8542_ (.CLK(clknet_leaf_50_clk),
    .D(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.register[15] ));
 sky130_fd_sc_hd__dfxtp_1 _8543_ (.CLK(clknet_leaf_51_clk),
    .D(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.register[16] ));
 sky130_fd_sc_hd__dfxtp_1 _8544_ (.CLK(clknet_leaf_4_clk),
    .D(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.register[17] ));
 sky130_fd_sc_hd__dfxtp_1 _8545_ (.CLK(clknet_leaf_5_clk),
    .D(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.register[18] ));
 sky130_fd_sc_hd__dfxtp_1 _8546_ (.CLK(clknet_leaf_50_clk),
    .D(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.register[19] ));
 sky130_fd_sc_hd__dfxtp_1 _8547_ (.CLK(clknet_leaf_51_clk),
    .D(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.register[20] ));
 sky130_fd_sc_hd__dfxtp_1 _8548_ (.CLK(clknet_leaf_3_clk),
    .D(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.register[21] ));
 sky130_fd_sc_hd__dfxtp_1 _8549_ (.CLK(clknet_leaf_4_clk),
    .D(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.register[22] ));
 sky130_fd_sc_hd__dfxtp_1 _8550_ (.CLK(clknet_leaf_50_clk),
    .D(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.register[23] ));
 sky130_fd_sc_hd__dfxtp_1 _8551_ (.CLK(clknet_leaf_51_clk),
    .D(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.register[24] ));
 sky130_fd_sc_hd__dfxtp_1 _8552_ (.CLK(clknet_leaf_3_clk),
    .D(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.register[25] ));
 sky130_fd_sc_hd__dfxtp_1 _8553_ (.CLK(clknet_leaf_4_clk),
    .D(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.register[26] ));
 sky130_fd_sc_hd__dfxtp_1 _8554_ (.CLK(clknet_leaf_51_clk),
    .D(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.register[27] ));
 sky130_fd_sc_hd__dfxtp_1 _8555_ (.CLK(clknet_leaf_6_clk),
    .D(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.register[28] ));
 sky130_fd_sc_hd__dfxtp_1 _8556_ (.CLK(clknet_leaf_3_clk),
    .D(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.register[29] ));
 sky130_fd_sc_hd__dfxtp_1 _8557_ (.CLK(clknet_leaf_4_clk),
    .D(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.register[30] ));
 sky130_fd_sc_hd__dfxtp_1 _8558_ (.CLK(clknet_leaf_51_clk),
    .D(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.register[31] ));
 sky130_fd_sc_hd__dfxtp_1 _8559_ (.CLK(clknet_leaf_40_clk),
    .D(_0601_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_shift.b[4] ));
 sky130_fd_sc_hd__dfxtp_1 _8560_ (.CLK(clknet_leaf_51_clk),
    .D(_0602_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.cy ));
 sky130_fd_sc_hd__dfxtp_1 _8561_ (.CLK(clknet_leaf_50_clk),
    .D(_0603_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.register[0] ));
 sky130_fd_sc_hd__dfxtp_1 _8562_ (.CLK(clknet_leaf_48_clk),
    .D(_0604_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.register[1] ));
 sky130_fd_sc_hd__dfxtp_1 _8563_ (.CLK(clknet_leaf_50_clk),
    .D(_0605_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.register[2] ));
 sky130_fd_sc_hd__dfxtp_1 _8564_ (.CLK(clknet_leaf_47_clk),
    .D(_0606_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.register[3] ));
 sky130_fd_sc_hd__clkbuf_4 _8565_ (.A(net1),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uio_oe[0]));
 sky130_fd_sc_hd__clkbuf_4 _8566_ (.A(uio_oe[5]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uio_oe[1]));
 sky130_fd_sc_hd__clkbuf_4 _8567_ (.A(uio_oe[5]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uio_oe[2]));
 sky130_fd_sc_hd__clkbuf_4 _8568_ (.A(net1),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uio_oe[3]));
 sky130_fd_sc_hd__clkbuf_4 _8569_ (.A(uio_oe[5]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uio_oe[4]));
 sky130_fd_sc_hd__clkbuf_4 _8570_ (.A(net1),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uio_oe[6]));
 sky130_fd_sc_hd__clkbuf_4 _8571_ (.A(net1),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uio_oe[7]));
 sky130_fd_sc_hd__clkbuf_4 _8572_ (.A(\i_tinyqv.mem.q_ctrl.spi_flash_select ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uio_out[0]));
 sky130_fd_sc_hd__clkbuf_4 _8573_ (.A(\i_tinyqv.mem.q_ctrl.spi_clk_out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uio_out[3]));
 sky130_fd_sc_hd__clkbuf_4 _8574_ (.A(\i_tinyqv.mem.q_ctrl.spi_ram_a_select ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uio_out[6]));
 sky130_fd_sc_hd__clkbuf_4 _8575_ (.A(\i_tinyqv.mem.q_ctrl.spi_ram_b_select ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uio_out[7]));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_0_clk (.A(clknet_3_0__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_10_clk (.A(clknet_3_2__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_10_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_11_clk (.A(clknet_3_2__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_11_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_12_clk (.A(clknet_3_2__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_12_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_13_clk (.A(clknet_3_2__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_13_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_14_clk (.A(clknet_3_2__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_14_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_15_clk (.A(clknet_3_2__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_15_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_16_clk (.A(clknet_3_2__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_16_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_17_clk (.A(clknet_3_3__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_17_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_18_clk (.A(clknet_3_3__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_18_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_19_clk (.A(clknet_3_3__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_19_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_1_clk (.A(clknet_3_0__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_1_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_20_clk (.A(clknet_3_3__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_20_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_21_clk (.A(clknet_3_3__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_21_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_22_clk (.A(clknet_3_3__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_22_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_23_clk (.A(clknet_3_6__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_23_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_24_clk (.A(clknet_3_6__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_24_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_25_clk (.A(clknet_3_6__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_25_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_26_clk (.A(clknet_3_6__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_26_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_27_clk (.A(clknet_3_6__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_27_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_28_clk (.A(clknet_3_6__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_28_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_29_clk (.A(clknet_3_7__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_29_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_2_clk (.A(clknet_3_0__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_2_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_30_clk (.A(clknet_3_7__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_30_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_31_clk (.A(clknet_3_7__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_31_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_32_clk (.A(clknet_3_7__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_32_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_33_clk (.A(clknet_3_7__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_33_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_34_clk (.A(clknet_3_7__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_34_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_35_clk (.A(clknet_3_7__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_35_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_36_clk (.A(clknet_3_6__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_36_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_37_clk (.A(clknet_3_4__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_37_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_38_clk (.A(clknet_3_4__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_38_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_39_clk (.A(clknet_3_5__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_39_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_3_clk (.A(clknet_3_0__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_3_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_40_clk (.A(clknet_3_5__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_40_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_41_clk (.A(clknet_3_5__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_41_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_42_clk (.A(clknet_3_5__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_42_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_43_clk (.A(clknet_3_5__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_43_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_44_clk (.A(clknet_3_5__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_44_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_45_clk (.A(clknet_3_4__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_45_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_46_clk (.A(clknet_3_4__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_46_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_47_clk (.A(clknet_3_4__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_47_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_48_clk (.A(clknet_3_4__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_48_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_49_clk (.A(clknet_3_4__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_49_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_4_clk (.A(clknet_3_0__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_4_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_50_clk (.A(clknet_3_4__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_50_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_51_clk (.A(clknet_3_1__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_51_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_52_clk (.A(clknet_3_1__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_52_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_53_clk (.A(clknet_3_1__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_53_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_54_clk (.A(clknet_3_1__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_54_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_55_clk (.A(clknet_3_1__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_55_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_56_clk (.A(clknet_3_1__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_56_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_57_clk (.A(clknet_3_0__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_57_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_58_clk (.A(clknet_3_0__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_58_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_59_clk (.A(clknet_3_0__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_59_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_5_clk (.A(clknet_3_0__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_5_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_6_clk (.A(clknet_3_1__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_6_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_7_clk (.A(clknet_3_3__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_7_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_8_clk (.A(clknet_3_3__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_8_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_9_clk (.A(clknet_3_2__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_9_clk));
 sky130_fd_sc_hd__clkbuf_2 clone11 (.A(_1398_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net40));
 sky130_fd_sc_hd__buf_6 clone3 (.A(_1638_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net32));
 sky130_fd_sc_hd__o21a_1 clone7 (.A1(_1410_),
    .A2(_1339_),
    .B1(_1411_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net36));
 sky130_fd_sc_hd__buf_2 clone8 (.A(\i_tinyqv.cpu.i_core.i_registers.rs1[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net324));
 sky130_fd_sc_hd__dlygate4sd3_1 hold100 (.A(\i_tinyqv.cpu.data_out[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net129));
 sky130_fd_sc_hd__dlygate4sd3_1 hold101 (.A(\i_tinyqv.cpu.data_out[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net130));
 sky130_fd_sc_hd__dlygate4sd3_1 hold102 (.A(\i_tinyqv.cpu.data_out[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net131));
 sky130_fd_sc_hd__dlygate4sd3_1 hold103 (.A(\i_tinyqv.cpu.data_out[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net132));
 sky130_fd_sc_hd__dlygate4sd3_1 hold104 (.A(\i_tinyqv.mem.q_ctrl.spi_in_buffer[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net133));
 sky130_fd_sc_hd__dlygate4sd3_1 hold105 (.A(_2903_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net134));
 sky130_fd_sc_hd__dlygate4sd3_1 hold106 (.A(\i_tinyqv.cpu.imm[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net135));
 sky130_fd_sc_hd__dlygate4sd3_1 hold107 (.A(\i_tinyqv.cpu.data_out[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net136));
 sky130_fd_sc_hd__dlygate4sd3_1 hold108 (.A(\i_tinyqv.cpu.data_addr[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net137));
 sky130_fd_sc_hd__dlygate4sd3_1 hold109 (.A(\i_tinyqv.cpu.i_core.load_done ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net138));
 sky130_fd_sc_hd__dlygate4sd3_1 hold110 (.A(_0084_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net139));
 sky130_fd_sc_hd__dlygate4sd3_1 hold111 (.A(\i_tinyqv.cpu.data_out[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net140));
 sky130_fd_sc_hd__dlygate4sd3_1 hold112 (.A(\i_tinyqv.cpu.alu_op[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net141));
 sky130_fd_sc_hd__dlygate4sd3_1 hold113 (.A(\i_uart_rx.cycle_counter[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net142));
 sky130_fd_sc_hd__dlygate4sd3_1 hold114 (.A(\i_tinyqv.cpu.data_out[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net143));
 sky130_fd_sc_hd__dlygate4sd3_1 hold115 (.A(\i_tinyqv.cpu.load_started ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net144));
 sky130_fd_sc_hd__dlygate4sd3_1 hold116 (.A(\i_tinyqv.mem.q_ctrl.spi_data_oe[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net145));
 sky130_fd_sc_hd__dlygate4sd3_1 hold117 (.A(\i_tinyqv.cpu.imm[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net146));
 sky130_fd_sc_hd__dlygate4sd3_1 hold118 (.A(\i_tinyqv.mem.q_ctrl.addr[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net147));
 sky130_fd_sc_hd__dlygate4sd3_1 hold119 (.A(\i_uart_rx.cycle_counter[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net148));
 sky130_fd_sc_hd__dlygate4sd3_1 hold120 (.A(\i_tinyqv.cpu.data_out[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net149));
 sky130_fd_sc_hd__dlygate4sd3_1 hold121 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[7][2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net150));
 sky130_fd_sc_hd__dlygate4sd3_1 hold122 (.A(\i_tinyqv.mem.q_ctrl.addr[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net151));
 sky130_fd_sc_hd__dlygate4sd3_1 hold123 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[6][3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net152));
 sky130_fd_sc_hd__dlygate4sd3_1 hold124 (.A(\i_tinyqv.mem.q_ctrl.addr[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net153));
 sky130_fd_sc_hd__dlygate4sd3_1 hold125 (.A(\i_tinyqv.cpu.additional_mem_ops[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net154));
 sky130_fd_sc_hd__clkbuf_2 hold126 (.A(\i_tinyqv.mem.q_ctrl.spi_clk_out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net155));
 sky130_fd_sc_hd__dlygate4sd3_1 hold127 (.A(\i_tinyqv.cpu.data_out[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net156));
 sky130_fd_sc_hd__dlygate4sd3_1 hold128 (.A(\i_uart_tx.cycle_counter[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net157));
 sky130_fd_sc_hd__dlygate4sd3_1 hold129 (.A(\i_tinyqv.cpu.i_core.mcause[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net158));
 sky130_fd_sc_hd__dlygate4sd3_1 hold130 (.A(\i_tinyqv.cpu.i_core.mcause[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net159));
 sky130_fd_sc_hd__dlygate4sd3_1 hold131 (.A(\i_uart_rx.recieved_data[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net160));
 sky130_fd_sc_hd__dlygate4sd3_1 hold132 (.A(\i_tinyqv.cpu.data_addr[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net161));
 sky130_fd_sc_hd__dlygate4sd3_1 hold133 (.A(\i_spi.clock_divider[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net162));
 sky130_fd_sc_hd__dlygate4sd3_1 hold134 (.A(_0203_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net163));
 sky130_fd_sc_hd__dlygate4sd3_1 hold135 (.A(\i_uart_tx.fsm_state[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net164));
 sky130_fd_sc_hd__dlygate4sd3_1 hold136 (.A(_2232_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net165));
 sky130_fd_sc_hd__dlygate4sd3_1 hold137 (.A(_0130_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net166));
 sky130_fd_sc_hd__dlygate4sd3_1 hold138 (.A(\i_tinyqv.mem.q_ctrl.spi_in_buffer[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net167));
 sky130_fd_sc_hd__dlygate4sd3_1 hold139 (.A(_2902_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net168));
 sky130_fd_sc_hd__dlygate4sd3_1 hold140 (.A(\i_spi.dc_in ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net169));
 sky130_fd_sc_hd__dlygate4sd3_1 hold141 (.A(\i_uart_tx.cycle_counter[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net170));
 sky130_fd_sc_hd__dlygate4sd3_1 hold142 (.A(_2219_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net171));
 sky130_fd_sc_hd__dlygate4sd3_1 hold143 (.A(\i_uart_rx.recieved_data[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net172));
 sky130_fd_sc_hd__dlygate4sd3_1 hold144 (.A(\i_tinyqv.cpu.data_addr[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net173));
 sky130_fd_sc_hd__dlygate4sd3_1 hold145 (.A(\i_uart_tx.cycle_counter[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net174));
 sky130_fd_sc_hd__dlygate4sd3_1 hold146 (.A(\i_tinyqv.cpu.data_out[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net175));
 sky130_fd_sc_hd__dlygate4sd3_1 hold147 (.A(\i_tinyqv.cpu.i_core.i_instrret.data[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net176));
 sky130_fd_sc_hd__dlygate4sd3_1 hold148 (.A(\i_tinyqv.cpu.data_addr[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net177));
 sky130_fd_sc_hd__dlygate4sd3_1 hold149 (.A(\i_uart_rx.cycle_counter[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net178));
 sky130_fd_sc_hd__dlygate4sd3_1 hold150 (.A(\i_tinyqv.cpu.i_core.mie[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net179));
 sky130_fd_sc_hd__dlygate4sd3_1 hold151 (.A(\i_tinyqv.cpu.data_ready_latch ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net180));
 sky130_fd_sc_hd__dlygate4sd3_1 hold152 (.A(\i_tinyqv.cpu.data_addr[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net181));
 sky130_fd_sc_hd__dlygate4sd3_1 hold153 (.A(\i_tinyqv.cpu.i_core.mie[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net182));
 sky130_fd_sc_hd__dlygate4sd3_1 hold154 (.A(\i_tinyqv.cpu.instr_fetch_started ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net183));
 sky130_fd_sc_hd__dlygate4sd3_1 hold155 (.A(\i_spi.end_txn_reg ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net184));
 sky130_fd_sc_hd__dlygate4sd3_1 hold156 (.A(_0199_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net185));
 sky130_fd_sc_hd__dlygate4sd3_1 hold157 (.A(\i_spi.end_txn ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net186));
 sky130_fd_sc_hd__dlygate4sd3_1 hold158 (.A(\i_tinyqv.mem.q_ctrl.addr[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net187));
 sky130_fd_sc_hd__dlygate4sd3_1 hold159 (.A(\i_debug_uart_tx.cycle_counter[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net188));
 sky130_fd_sc_hd__dlygate4sd3_1 hold160 (.A(\i_tinyqv.mem.q_ctrl.addr[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net189));
 sky130_fd_sc_hd__dlygate4sd3_1 hold161 (.A(\i_tinyqv.cpu.imm[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net190));
 sky130_fd_sc_hd__dlygate4sd3_1 hold162 (.A(\i_uart_rx.bit_sample ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net191));
 sky130_fd_sc_hd__dlygate4sd3_1 hold163 (.A(\i_tinyqv.cpu.i_core.mip[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net192));
 sky130_fd_sc_hd__dlygate4sd3_1 hold164 (.A(\i_uart_rx.rxd_reg[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net193));
 sky130_fd_sc_hd__dlygate4sd3_1 hold165 (.A(\i_spi.bits_remaining[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net194));
 sky130_fd_sc_hd__dlygate4sd3_1 hold166 (.A(_0196_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net195));
 sky130_fd_sc_hd__dlygate4sd3_1 hold167 (.A(\i_tinyqv.cpu.instr_len[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net196));
 sky130_fd_sc_hd__buf_1 hold168 (.A(\i_debug_uart_tx.uart_tx_data[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net197));
 sky130_fd_sc_hd__dlygate4sd3_1 hold169 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[1][0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net198));
 sky130_fd_sc_hd__dlygate4sd3_1 hold170 (.A(\i_uart_rx.cycle_counter[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net199));
 sky130_fd_sc_hd__dlygate4sd3_1 hold171 (.A(\i_tinyqv.cpu.i_core.mie[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net200));
 sky130_fd_sc_hd__dlygate4sd3_1 hold172 (.A(\i_uart_rx.recieved_data[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net201));
 sky130_fd_sc_hd__dlygate4sd3_1 hold173 (.A(_0142_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net202));
 sky130_fd_sc_hd__dlygate4sd3_1 hold174 (.A(\i_tinyqv.cpu.i_core.i_registers.registers[1][25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net203));
 sky130_fd_sc_hd__dlygate4sd3_1 hold175 (.A(\i_spi.clock_divider[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net204));
 sky130_fd_sc_hd__dlygate4sd3_1 hold176 (.A(\i_debug_uart_tx.data_to_send[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net205));
 sky130_fd_sc_hd__buf_1 hold177 (.A(\i_uart_tx.cycle_counter[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net206));
 sky130_fd_sc_hd__dlygate4sd3_1 hold178 (.A(\i_uart_rx.recieved_data[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net207));
 sky130_fd_sc_hd__dlygate4sd3_1 hold179 (.A(\i_tinyqv.mem.q_ctrl.spi_ram_a_select ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net208));
 sky130_fd_sc_hd__dlygate4sd3_1 hold180 (.A(\i_tinyqv.cpu.is_system ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net209));
 sky130_fd_sc_hd__dlygate4sd3_1 hold181 (.A(\i_tinyqv.mem.q_ctrl.spi_ram_b_select ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net210));
 sky130_fd_sc_hd__dlygate4sd3_1 hold182 (.A(\i_tinyqv.cpu.i_core.mepc[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net211));
 sky130_fd_sc_hd__dlygate4sd3_1 hold183 (.A(\i_tinyqv.cpu.is_lui ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net212));
 sky130_fd_sc_hd__dlygate4sd3_1 hold184 (.A(\i_tinyqv.cpu.imm[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net213));
 sky130_fd_sc_hd__dlygate4sd3_1 hold185 (.A(\i_uart_tx.cycle_counter[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net214));
 sky130_fd_sc_hd__dlygate4sd3_1 hold186 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[12][0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net215));
 sky130_fd_sc_hd__dlygate4sd3_1 hold187 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[7][1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net216));
 sky130_fd_sc_hd__dlygate4sd3_1 hold188 (.A(\i_tinyqv.cpu.i_core.i_instrret.data[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net217));
 sky130_fd_sc_hd__dlygate4sd3_1 hold189 (.A(\i_tinyqv.cpu.i_core.time_hi[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net218));
 sky130_fd_sc_hd__dlygate4sd3_1 hold190 (.A(\i_uart_tx.cycle_counter[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net219));
 sky130_fd_sc_hd__dlygate4sd3_1 hold191 (.A(\i_spi.read_latency ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net220));
 sky130_fd_sc_hd__dlygate4sd3_1 hold192 (.A(\i_tinyqv.cpu.i_core.imm_lo[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net221));
 sky130_fd_sc_hd__dlygate4sd3_1 hold193 (.A(\i_tinyqv.cpu.i_core.mepc[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net222));
 sky130_fd_sc_hd__dlygate4sd3_1 hold194 (.A(\i_tinyqv.cpu.i_core.mepc[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net223));
 sky130_fd_sc_hd__dlygate4sd3_1 hold195 (.A(\i_uart_rx.cycle_counter[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net224));
 sky130_fd_sc_hd__dlygate4sd3_1 hold196 (.A(\i_uart_rx.recieved_data[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net225));
 sky130_fd_sc_hd__dlygate4sd3_1 hold197 (.A(\i_tinyqv.cpu.i_core.mepc[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net226));
 sky130_fd_sc_hd__dlygate4sd3_1 hold198 (.A(\i_tinyqv.cpu.imm[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net227));
 sky130_fd_sc_hd__dlygate4sd3_1 hold199 (.A(\i_tinyqv.cpu.i_core.mepc[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net228));
 sky130_fd_sc_hd__dlygate4sd3_1 hold200 (.A(\i_tinyqv.mem.qspi_data_buf[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net229));
 sky130_fd_sc_hd__dlygate4sd3_1 hold201 (.A(\i_tinyqv.cpu.i_core.mie[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net230));
 sky130_fd_sc_hd__dlygate4sd3_1 hold202 (.A(\i_tinyqv.cpu.imm[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net231));
 sky130_fd_sc_hd__dlygate4sd3_1 hold203 (.A(\i_tinyqv.cpu.i_core.mepc[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net232));
 sky130_fd_sc_hd__dlygate4sd3_1 hold204 (.A(\i_debug_uart_tx.data_to_send[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net233));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold205 (.A(\i_debug_uart_tx.uart_tx_data[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net234));
 sky130_fd_sc_hd__dlygate4sd3_1 hold206 (.A(\i_tinyqv.cpu.i_core.cycle_count[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net235));
 sky130_fd_sc_hd__dlygate4sd3_1 hold207 (.A(\i_tinyqv.cpu.data_ready_core ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net236));
 sky130_fd_sc_hd__dlygate4sd3_1 hold208 (.A(\i_debug_uart_tx.uart_tx_data[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net237));
 sky130_fd_sc_hd__dlygate4sd3_1 hold209 (.A(\i_debug_uart_tx.uart_tx_data[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net238));
 sky130_fd_sc_hd__dlygate4sd3_1 hold210 (.A(\i_spi.bits_remaining[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net239));
 sky130_fd_sc_hd__dlygate4sd3_1 hold211 (.A(\i_uart_rx.recieved_data[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net240));
 sky130_fd_sc_hd__dlygate4sd3_1 hold212 (.A(\i_uart_rx.recieved_data[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net241));
 sky130_fd_sc_hd__dlygate4sd3_1 hold213 (.A(\i_tinyqv.cpu.additional_mem_ops[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net242));
 sky130_fd_sc_hd__dlygate4sd3_1 hold214 (.A(\i_tinyqv.cpu.alu_op[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net243));
 sky130_fd_sc_hd__dlygate4sd3_1 hold215 (.A(\i_tinyqv.cpu.i_core.mepc[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net244));
 sky130_fd_sc_hd__dlygate4sd3_1 hold216 (.A(\i_tinyqv.mem.data_from_read[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net245));
 sky130_fd_sc_hd__dlygate4sd3_1 hold217 (.A(\i_tinyqv.cpu.i_core.time_hi[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net246));
 sky130_fd_sc_hd__dlygate4sd3_1 hold218 (.A(\i_uart_rx.cycle_counter[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net247));
 sky130_fd_sc_hd__dlygate4sd3_1 hold219 (.A(\i_tinyqv.cpu.i_core.i_cycles.cy ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net248));
 sky130_fd_sc_hd__dlygate4sd3_1 hold220 (.A(\i_tinyqv.cpu.is_alu_imm ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net249));
 sky130_fd_sc_hd__dlygate4sd3_1 hold221 (.A(\i_tinyqv.cpu.i_core.last_interrupt_req[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net250));
 sky130_fd_sc_hd__dlygate4sd3_1 hold222 (.A(_2085_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net251));
 sky130_fd_sc_hd__dlygate4sd3_1 hold223 (.A(\i_tinyqv.cpu.i_core.i_registers.rd[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net252));
 sky130_fd_sc_hd__dlygate4sd3_1 hold224 (.A(\i_tinyqv.mem.qspi_data_buf[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net253));
 sky130_fd_sc_hd__dlygate4sd3_1 hold225 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[9][1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net254));
 sky130_fd_sc_hd__dlygate4sd3_1 hold226 (.A(\i_debug_uart_tx.data_to_send[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net255));
 sky130_fd_sc_hd__dlygate4sd3_1 hold227 (.A(\i_tinyqv.mem.qspi_data_buf[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net256));
 sky130_fd_sc_hd__dlygate4sd3_1 hold228 (.A(\i_tinyqv.cpu.imm[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net257));
 sky130_fd_sc_hd__dlygate4sd3_1 hold229 (.A(\i_tinyqv.cpu.i_core.mem_op[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net258));
 sky130_fd_sc_hd__dlygate4sd3_1 hold230 (.A(\i_tinyqv.cpu.imm[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net259));
 sky130_fd_sc_hd__dlygate4sd3_1 hold231 (.A(\i_tinyqv.cpu.instr_data[3][3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net260));
 sky130_fd_sc_hd__dlygate4sd3_1 hold232 (.A(\i_tinyqv.mem.qspi_data_buf[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net261));
 sky130_fd_sc_hd__dlygate4sd3_1 hold233 (.A(\i_tinyqv.cpu.i_core.mstatus_mpie ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net262));
 sky130_fd_sc_hd__dlygate4sd3_1 hold234 (.A(\i_tinyqv.cpu.instr_data[3][2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net263));
 sky130_fd_sc_hd__dlygate4sd3_1 hold235 (.A(\i_tinyqv.cpu.i_core.mepc[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net264));
 sky130_fd_sc_hd__dlygate4sd3_1 hold236 (.A(\i_tinyqv.mem.q_ctrl.nibbles_remaining[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net265));
 sky130_fd_sc_hd__dlygate4sd3_1 hold237 (.A(\i_tinyqv.cpu.instr_data[0][14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net266));
 sky130_fd_sc_hd__dlygate4sd3_1 hold238 (.A(\i_tinyqv.mem.qspi_data_buf[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net267));
 sky130_fd_sc_hd__dlygate4sd3_1 hold239 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[1][1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net268));
 sky130_fd_sc_hd__dlygate4sd3_1 hold240 (.A(\i_tinyqv.mem.data_from_read[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net269));
 sky130_fd_sc_hd__dlygate4sd3_1 hold241 (.A(\i_uart_tx.fsm_state[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net270));
 sky130_fd_sc_hd__dlygate4sd3_1 hold242 (.A(\i_tinyqv.mem.q_ctrl.spi_in_buffer[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net271));
 sky130_fd_sc_hd__dlygate4sd3_1 hold243 (.A(\i_tinyqv.cpu.instr_data[3][13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net272));
 sky130_fd_sc_hd__dlygate4sd3_1 hold244 (.A(\i_debug_uart_tx.uart_tx_data[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net273));
 sky130_fd_sc_hd__dlygate4sd3_1 hold245 (.A(\i_tinyqv.mem.q_ctrl.spi_in_buffer[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net274));
 sky130_fd_sc_hd__dlygate4sd3_1 hold246 (.A(\i_tinyqv.mem.qspi_data_buf[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net275));
 sky130_fd_sc_hd__dlygate4sd3_1 hold247 (.A(\i_tinyqv.mem.qspi_data_buf[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net276));
 sky130_fd_sc_hd__dlygate4sd3_1 hold248 (.A(\i_tinyqv.mem.data_from_read[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net277));
 sky130_fd_sc_hd__dlygate4sd3_1 hold249 (.A(\i_debug_uart_tx.data_to_send[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net278));
 sky130_fd_sc_hd__dlygate4sd3_1 hold250 (.A(\i_tinyqv.mem.qspi_data_buf[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net279));
 sky130_fd_sc_hd__dlygate4sd3_1 hold251 (.A(\i_tinyqv.mem.data_from_read[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net280));
 sky130_fd_sc_hd__dlygate4sd3_1 hold252 (.A(\i_tinyqv.cpu.instr_data[3][15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net281));
 sky130_fd_sc_hd__dlygate4sd3_1 hold253 (.A(\i_spi.spi_dc ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net282));
 sky130_fd_sc_hd__dlygate4sd3_1 hold254 (.A(\i_tinyqv.cpu.instr_data[0][15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net283));
 sky130_fd_sc_hd__dlygate4sd3_1 hold255 (.A(\i_tinyqv.cpu.imm[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net284));
 sky130_fd_sc_hd__dlygate4sd3_1 hold256 (.A(\i_tinyqv.mem.data_from_read[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net285));
 sky130_fd_sc_hd__dlygate4sd3_1 hold257 (.A(\i_tinyqv.mem.qspi_data_buf[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net286));
 sky130_fd_sc_hd__dlygate4sd3_1 hold258 (.A(\i_tinyqv.mem.qspi_data_buf[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net287));
 sky130_fd_sc_hd__dlygate4sd3_1 hold259 (.A(\i_tinyqv.cpu.data_addr[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net288));
 sky130_fd_sc_hd__dlygate4sd3_1 hold260 (.A(\i_tinyqv.mem.q_ctrl.spi_flash_select ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net289));
 sky130_fd_sc_hd__dlygate4sd3_1 hold261 (.A(\i_tinyqv.mem.qspi_data_buf[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net290));
 sky130_fd_sc_hd__dlygate4sd3_1 hold262 (.A(\i_tinyqv.cpu.instr_data[0][3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net291));
 sky130_fd_sc_hd__dlygate4sd3_1 hold263 (.A(\i_tinyqv.mem.data_from_read[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net292));
 sky130_fd_sc_hd__dlygate4sd3_1 hold264 (.A(\i_tinyqv.mem.qspi_data_buf[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net293));
 sky130_fd_sc_hd__dlygate4sd3_1 hold265 (.A(\i_tinyqv.cpu.data_write_n[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net294));
 sky130_fd_sc_hd__dlygate4sd3_1 hold266 (.A(\i_tinyqv.cpu.i_core.imm_lo[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net295));
 sky130_fd_sc_hd__dlygate4sd3_1 hold267 (.A(\i_tinyqv.cpu.i_core.imm_lo[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net296));
 sky130_fd_sc_hd__dlygate4sd3_1 hold268 (.A(\i_tinyqv.cpu.data_addr[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net297));
 sky130_fd_sc_hd__dlygate4sd3_1 hold269 (.A(\i_tinyqv.cpu.data_addr[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net298));
 sky130_fd_sc_hd__dlygate4sd3_1 hold270 (.A(\i_tinyqv.cpu.data_addr[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net299));
 sky130_fd_sc_hd__dlygate4sd3_1 hold271 (.A(\i_tinyqv.cpu.data_addr[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net300));
 sky130_fd_sc_hd__dlygate4sd3_1 hold272 (.A(\i_tinyqv.mem.q_ctrl.addr[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net301));
 sky130_fd_sc_hd__dlygate4sd3_1 hold273 (.A(\i_tinyqv.mem.q_ctrl.addr[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net302));
 sky130_fd_sc_hd__dlygate4sd3_1 hold274 (.A(\i_tinyqv.mem.q_ctrl.addr[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net303));
 sky130_fd_sc_hd__dlygate4sd3_1 hold275 (.A(\i_tinyqv.mem.q_ctrl.addr[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net304));
 sky130_fd_sc_hd__dlygate4sd3_1 hold276 (.A(\i_tinyqv.mem.q_ctrl.addr[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net305));
 sky130_fd_sc_hd__dlygate4sd3_1 hold277 (.A(\i_uart_rx.cycle_counter[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net306));
 sky130_fd_sc_hd__dlygate4sd3_1 hold278 (.A(\i_uart_rx.cycle_counter[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net307));
 sky130_fd_sc_hd__dlygate4sd3_1 hold279 (.A(\i_spi.end_txn_reg ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net308));
 sky130_fd_sc_hd__dlygate4sd3_1 hold280 (.A(\i_debug_uart_tx.uart_tx_data[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net309));
 sky130_fd_sc_hd__dlygate4sd3_1 hold281 (.A(\i_tinyqv.mem.q_ctrl.addr[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net310));
 sky130_fd_sc_hd__dlygate4sd3_1 hold282 (.A(\i_tinyqv.mem.q_ctrl.spi_ram_b_select ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net311));
 sky130_fd_sc_hd__dlygate4sd3_1 hold283 (.A(\i_tinyqv.mem.q_ctrl.addr[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net312));
 sky130_fd_sc_hd__dlygate4sd3_1 hold284 (.A(\i_debug_uart_tx.uart_tx_data[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net313));
 sky130_fd_sc_hd__dlygate4sd3_1 hold285 (.A(\i_tinyqv.cpu.data_addr[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net314));
 sky130_fd_sc_hd__dlygate4sd3_1 hold286 (.A(\i_tinyqv.mem.q_ctrl.addr[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net315));
 sky130_fd_sc_hd__dlygate4sd3_1 hold287 (.A(\i_debug_uart_tx.uart_tx_data[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net316));
 sky130_fd_sc_hd__dlygate4sd3_1 hold288 (.A(\i_tinyqv.mem.q_ctrl.addr[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net317));
 sky130_fd_sc_hd__dlygate4sd3_1 hold289 (.A(\i_tinyqv.mem.q_ctrl.addr[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net318));
 sky130_fd_sc_hd__dlygate4sd3_1 hold290 (.A(\i_debug_uart_tx.uart_tx_data[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net319));
 sky130_fd_sc_hd__dlygate4sd3_1 hold60 (.A(\i_tinyqv.mem.q_ctrl.addr[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net89));
 sky130_fd_sc_hd__buf_1 hold61 (.A(\i_tinyqv.cpu.i_core.i_instrret.data[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net90));
 sky130_fd_sc_hd__dlygate4sd3_1 hold62 (.A(\i_uart_rx.cycle_counter[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net91));
 sky130_fd_sc_hd__dlygate4sd3_1 hold63 (.A(\i_tinyqv.cpu.i_core.i_instrret.data[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net92));
 sky130_fd_sc_hd__dlygate4sd3_1 hold64 (.A(\i_tinyqv.mem.q_ctrl.addr[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net93));
 sky130_fd_sc_hd__dlygate4sd3_1 hold65 (.A(\i_tinyqv.cpu.data_continue ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net94));
 sky130_fd_sc_hd__dlygate4sd3_1 hold66 (.A(\i_tinyqv.mem.q_ctrl.addr[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net95));
 sky130_fd_sc_hd__dlygate4sd3_1 hold67 (.A(\i_tinyqv.cpu.data_addr[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net96));
 sky130_fd_sc_hd__clkbuf_2 hold68 (.A(\i_debug_uart_tx.uart_tx_data[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net97));
 sky130_fd_sc_hd__clkbuf_2 hold69 (.A(\i_debug_uart_tx.uart_tx_data[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net98));
 sky130_fd_sc_hd__dlygate4sd3_1 hold70 (.A(\i_tinyqv.cpu.i_core.is_double_fault_r ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net99));
 sky130_fd_sc_hd__dlygate4sd3_1 hold71 (.A(\i_tinyqv.cpu.instr_data[3][0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net100));
 sky130_fd_sc_hd__dlygate4sd3_1 hold72 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[12][3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net101));
 sky130_fd_sc_hd__dlygate4sd3_1 hold73 (.A(\i_uart_tx.cycle_counter[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net102));
 sky130_fd_sc_hd__dlygate4sd3_1 hold74 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[12][2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net103));
 sky130_fd_sc_hd__dlygate4sd3_1 hold75 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[15][2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net104));
 sky130_fd_sc_hd__dlygate4sd3_1 hold76 (.A(\i_tinyqv.cpu.i_core.i_registers.registers[1][24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net105));
 sky130_fd_sc_hd__dlygate4sd3_1 hold77 (.A(\i_tinyqv.cpu.instr_data[3][1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net106));
 sky130_fd_sc_hd__dlygate4sd3_1 hold78 (.A(\i_tinyqv.cpu.data_out[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net107));
 sky130_fd_sc_hd__dlygate4sd3_1 hold79 (.A(\i_tinyqv.cpu.i_core.time_hi[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net108));
 sky130_fd_sc_hd__dlygate4sd3_1 hold80 (.A(\i_tinyqv.cpu.data_out[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net109));
 sky130_fd_sc_hd__dlygate4sd3_1 hold81 (.A(\i_tinyqv.cpu.data_out[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net110));
 sky130_fd_sc_hd__dlygate4sd3_1 hold82 (.A(\i_tinyqv.cpu.data_addr[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net111));
 sky130_fd_sc_hd__dlygate4sd3_1 hold83 (.A(\i_tinyqv.cpu.data_out[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net112));
 sky130_fd_sc_hd__dlygate4sd3_1 hold84 (.A(\i_tinyqv.cpu.data_out[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net113));
 sky130_fd_sc_hd__dlygate4sd3_1 hold85 (.A(\i_tinyqv.cpu.data_out[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net114));
 sky130_fd_sc_hd__dlygate4sd3_1 hold86 (.A(\i_tinyqv.cpu.data_out[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net115));
 sky130_fd_sc_hd__dlygate4sd3_1 hold87 (.A(\i_uart_tx.data_to_send[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net116));
 sky130_fd_sc_hd__clkbuf_2 hold88 (.A(\i_debug_uart_tx.uart_tx_data[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net117));
 sky130_fd_sc_hd__dlygate4sd3_1 hold89 (.A(\i_tinyqv.cpu.data_out[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net118));
 sky130_fd_sc_hd__dlygate4sd3_1 hold90 (.A(\i_tinyqv.cpu.data_out[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net119));
 sky130_fd_sc_hd__dlygate4sd3_1 hold91 (.A(\i_tinyqv.cpu.data_out[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net120));
 sky130_fd_sc_hd__dlygate4sd3_1 hold92 (.A(\i_tinyqv.cpu.i_core.cycle_count[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net121));
 sky130_fd_sc_hd__dlygate4sd3_1 hold93 (.A(\i_tinyqv.mem.q_ctrl.addr[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net122));
 sky130_fd_sc_hd__dlygate4sd3_1 hold94 (.A(\i_tinyqv.cpu.i_core.mcause[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net123));
 sky130_fd_sc_hd__dlygate4sd3_1 hold95 (.A(\i_tinyqv.cpu.data_out[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net124));
 sky130_fd_sc_hd__dlygate4sd3_1 hold96 (.A(\i_tinyqv.cpu.data_out[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net125));
 sky130_fd_sc_hd__dlygate4sd3_1 hold97 (.A(\i_tinyqv.mem.q_ctrl.addr[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net126));
 sky130_fd_sc_hd__dlygate4sd3_1 hold98 (.A(\i_tinyqv.cpu.i_core.is_interrupt ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net127));
 sky130_fd_sc_hd__dlygate4sd3_1 hold99 (.A(_0029_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net128));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_cycles.i_regbuf[10]  (.A(\i_tinyqv.cpu.i_core.i_cycles.register[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[10] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_cycles.i_regbuf[11]  (.A(\i_tinyqv.cpu.i_core.i_cycles.register[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[11] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_cycles.i_regbuf[12]  (.A(\i_tinyqv.cpu.i_core.i_cycles.register[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[12] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_cycles.i_regbuf[13]  (.A(\i_tinyqv.cpu.i_core.i_cycles.register[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[13] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_cycles.i_regbuf[14]  (.A(\i_tinyqv.cpu.i_core.i_cycles.register[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[14] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_cycles.i_regbuf[15]  (.A(\i_tinyqv.cpu.i_core.i_cycles.register[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[15] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_cycles.i_regbuf[16]  (.A(\i_tinyqv.cpu.i_core.i_cycles.register[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[16] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_cycles.i_regbuf[17]  (.A(\i_tinyqv.cpu.i_core.i_cycles.register[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[17] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_cycles.i_regbuf[18]  (.A(\i_tinyqv.cpu.i_core.i_cycles.register[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[18] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_cycles.i_regbuf[19]  (.A(\i_tinyqv.cpu.i_core.i_cycles.register[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[19] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_cycles.i_regbuf[20]  (.A(\i_tinyqv.cpu.i_core.i_cycles.register[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[20] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_cycles.i_regbuf[21]  (.A(\i_tinyqv.cpu.i_core.i_cycles.register[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[21] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_cycles.i_regbuf[22]  (.A(\i_tinyqv.cpu.i_core.i_cycles.register[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[22] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_cycles.i_regbuf[23]  (.A(\i_tinyqv.cpu.i_core.i_cycles.register[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[23] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_cycles.i_regbuf[24]  (.A(\i_tinyqv.cpu.i_core.i_cycles.register[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[24] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_cycles.i_regbuf[25]  (.A(\i_tinyqv.cpu.i_core.i_cycles.register[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[25] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_cycles.i_regbuf[26]  (.A(\i_tinyqv.cpu.i_core.i_cycles.register[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[26] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_cycles.i_regbuf[27]  (.A(\i_tinyqv.cpu.i_core.i_cycles.register[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[27] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_cycles.i_regbuf[28]  (.A(\i_tinyqv.cpu.i_core.i_cycles.register[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[28] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_cycles.i_regbuf[29]  (.A(\i_tinyqv.cpu.i_core.i_cycles.register[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[29] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_cycles.i_regbuf[30]  (.A(\i_tinyqv.cpu.i_core.i_cycles.register[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[30] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_cycles.i_regbuf[31]  (.A(\i_tinyqv.cpu.i_core.i_cycles.register[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[31] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_cycles.i_regbuf[4]  (.A(\i_tinyqv.cpu.i_core.cycle_count_wide[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[4] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_cycles.i_regbuf[5]  (.A(\i_tinyqv.cpu.i_core.cycle_count_wide[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[5] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_cycles.i_regbuf[6]  (.A(\i_tinyqv.cpu.i_core.cycle_count_wide[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[6] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_cycles.i_regbuf[7]  (.A(\i_tinyqv.cpu.i_core.i_cycles.register[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[7] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_cycles.i_regbuf[8]  (.A(\i_tinyqv.cpu.i_core.i_cycles.register[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[8] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_cycles.i_regbuf[9]  (.A(\i_tinyqv.cpu.i_core.i_cycles.register[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[9] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_instrret.i_regbuf[10]  (.A(\i_tinyqv.cpu.i_core.i_instrret.register[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[10] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_instrret.i_regbuf[11]  (.A(\i_tinyqv.cpu.i_core.i_instrret.register[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[11] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_instrret.i_regbuf[12]  (.A(\i_tinyqv.cpu.i_core.i_instrret.register[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[12] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_instrret.i_regbuf[13]  (.A(\i_tinyqv.cpu.i_core.i_instrret.register[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[13] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_instrret.i_regbuf[14]  (.A(\i_tinyqv.cpu.i_core.i_instrret.register[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[14] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_instrret.i_regbuf[15]  (.A(\i_tinyqv.cpu.i_core.i_instrret.register[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[15] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_instrret.i_regbuf[16]  (.A(\i_tinyqv.cpu.i_core.i_instrret.register[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[16] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_instrret.i_regbuf[17]  (.A(\i_tinyqv.cpu.i_core.i_instrret.register[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[17] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_instrret.i_regbuf[18]  (.A(\i_tinyqv.cpu.i_core.i_instrret.register[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[18] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_instrret.i_regbuf[19]  (.A(\i_tinyqv.cpu.i_core.i_instrret.register[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[19] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_instrret.i_regbuf[20]  (.A(\i_tinyqv.cpu.i_core.i_instrret.register[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[20] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_instrret.i_regbuf[21]  (.A(\i_tinyqv.cpu.i_core.i_instrret.register[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[21] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_instrret.i_regbuf[22]  (.A(\i_tinyqv.cpu.i_core.i_instrret.register[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[22] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_instrret.i_regbuf[23]  (.A(\i_tinyqv.cpu.i_core.i_instrret.register[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[23] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_instrret.i_regbuf[24]  (.A(\i_tinyqv.cpu.i_core.i_instrret.register[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[24] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_instrret.i_regbuf[25]  (.A(\i_tinyqv.cpu.i_core.i_instrret.register[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[25] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_instrret.i_regbuf[26]  (.A(\i_tinyqv.cpu.i_core.i_instrret.register[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[26] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_instrret.i_regbuf[27]  (.A(\i_tinyqv.cpu.i_core.i_instrret.register[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[27] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_instrret.i_regbuf[28]  (.A(\i_tinyqv.cpu.i_core.i_instrret.register[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[28] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_instrret.i_regbuf[29]  (.A(\i_tinyqv.cpu.i_core.i_instrret.register[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[29] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_instrret.i_regbuf[30]  (.A(\i_tinyqv.cpu.i_core.i_instrret.register[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[30] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_instrret.i_regbuf[31]  (.A(\i_tinyqv.cpu.i_core.i_instrret.register[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[31] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_instrret.i_regbuf[4]  (.A(\i_tinyqv.cpu.i_core.i_instrret.register[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[4] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_instrret.i_regbuf[5]  (.A(\i_tinyqv.cpu.i_core.i_instrret.register[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[5] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_instrret.i_regbuf[6]  (.A(\i_tinyqv.cpu.i_core.i_instrret.register[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[6] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_instrret.i_regbuf[7]  (.A(\i_tinyqv.cpu.i_core.i_instrret.register[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[7] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_instrret.i_regbuf[8]  (.A(\i_tinyqv.cpu.i_core.i_instrret.register[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[8] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_instrret.i_regbuf[9]  (.A(\i_tinyqv.cpu.i_core.i_instrret.register[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[9] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.i_regbuf[10]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[10][14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.reg_buf[10] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.i_regbuf[11]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[10][15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.reg_buf[11] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.i_regbuf[12]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[10][16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.reg_buf[12] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.i_regbuf[13]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[10][17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.reg_buf[13] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.i_regbuf[14]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[10][18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.reg_buf[14] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.i_regbuf[15]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[10][19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.reg_buf[15] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.i_regbuf[16]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[10][20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.reg_buf[16] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.i_regbuf[17]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[10][21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.reg_buf[17] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.i_regbuf[18]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[10][22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.reg_buf[18] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.i_regbuf[19]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[10][23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.reg_buf[19] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.i_regbuf[20]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[10][24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.reg_buf[20] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.i_regbuf[21]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[10][25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.reg_buf[21] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.i_regbuf[22]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[10][26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.reg_buf[22] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.i_regbuf[23]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[10][27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.reg_buf[23] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.i_regbuf[24]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[10][28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.reg_buf[24] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.i_regbuf[25]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[10][29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.reg_buf[25] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.i_regbuf[26]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[10][30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.reg_buf[26] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.i_regbuf[27]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[10][31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.reg_buf[27] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.i_regbuf[28]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[10][0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.reg_buf[28] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.i_regbuf[29]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[10][1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.reg_buf[29] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.i_regbuf[30]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[10][2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.reg_buf[30] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.i_regbuf[31]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[10][3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.reg_buf[31] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.i_regbuf[4]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[10][8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.reg_buf[4] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.i_regbuf[5]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[10][9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.reg_buf[5] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.i_regbuf[6]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[10][10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.reg_buf[6] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.i_regbuf[7]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[10][11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.reg_buf[7] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.i_regbuf[8]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[10][12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.reg_buf[8] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.i_regbuf[9]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[10][13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.genblk1.reg_buf[9] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.i_regbuf[10]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[11][14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.reg_buf[10] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.i_regbuf[11]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[11][15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.reg_buf[11] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.i_regbuf[12]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[11][16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.reg_buf[12] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.i_regbuf[13]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[11][17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.reg_buf[13] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.i_regbuf[14]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[11][18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.reg_buf[14] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.i_regbuf[15]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[11][19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.reg_buf[15] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.i_regbuf[16]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[11][20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.reg_buf[16] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.i_regbuf[17]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[11][21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.reg_buf[17] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.i_regbuf[18]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[11][22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.reg_buf[18] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.i_regbuf[19]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[11][23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.reg_buf[19] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.i_regbuf[20]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[11][24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.reg_buf[20] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.i_regbuf[21]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[11][25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.reg_buf[21] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.i_regbuf[22]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[11][26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.reg_buf[22] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.i_regbuf[23]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[11][27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.reg_buf[23] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.i_regbuf[24]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[11][28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.reg_buf[24] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.i_regbuf[25]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[11][29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.reg_buf[25] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.i_regbuf[26]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[11][30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.reg_buf[26] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.i_regbuf[27]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[11][31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.reg_buf[27] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.i_regbuf[28]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[11][0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.reg_buf[28] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.i_regbuf[29]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[11][1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.reg_buf[29] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.i_regbuf[30]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[11][2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.reg_buf[30] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.i_regbuf[31]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[11][3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.reg_buf[31] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.i_regbuf[4]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[11][8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.reg_buf[4] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.i_regbuf[5]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[11][9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.reg_buf[5] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.i_regbuf[6]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[11][10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.reg_buf[6] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.i_regbuf[7]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[11][11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.reg_buf[7] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.i_regbuf[8]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[11][12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.reg_buf[8] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.i_regbuf[9]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[11][13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.genblk1.reg_buf[9] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.i_regbuf[10]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[12][14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.reg_buf[10] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.i_regbuf[11]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[12][15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.reg_buf[11] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.i_regbuf[12]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[12][16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.reg_buf[12] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.i_regbuf[13]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[12][17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.reg_buf[13] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.i_regbuf[14]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[12][18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.reg_buf[14] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.i_regbuf[15]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[12][19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.reg_buf[15] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.i_regbuf[16]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[12][20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.reg_buf[16] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.i_regbuf[17]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[12][21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.reg_buf[17] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.i_regbuf[18]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[12][22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.reg_buf[18] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.i_regbuf[19]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[12][23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.reg_buf[19] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.i_regbuf[20]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[12][24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.reg_buf[20] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.i_regbuf[21]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[12][25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.reg_buf[21] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.i_regbuf[22]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[12][26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.reg_buf[22] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.i_regbuf[23]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[12][27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.reg_buf[23] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.i_regbuf[24]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[12][28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.reg_buf[24] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.i_regbuf[25]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[12][29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.reg_buf[25] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.i_regbuf[26]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[12][30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.reg_buf[26] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.i_regbuf[27]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[12][31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.reg_buf[27] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.i_regbuf[28]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[12][0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.reg_buf[28] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.i_regbuf[29]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[12][1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.reg_buf[29] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.i_regbuf[30]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[12][2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.reg_buf[30] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.i_regbuf[31]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[12][3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.reg_buf[31] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.i_regbuf[4]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[12][8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.reg_buf[4] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.i_regbuf[5]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[12][9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.reg_buf[5] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.i_regbuf[6]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[12][10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.reg_buf[6] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.i_regbuf[7]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[12][11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.reg_buf[7] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.i_regbuf[8]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[12][12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.reg_buf[8] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.i_regbuf[9]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[12][13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.genblk1.reg_buf[9] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.i_regbuf[10]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[13][14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.reg_buf[10] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.i_regbuf[11]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[13][15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.reg_buf[11] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.i_regbuf[12]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[13][16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.reg_buf[12] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.i_regbuf[13]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[13][17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.reg_buf[13] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.i_regbuf[14]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[13][18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.reg_buf[14] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.i_regbuf[15]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[13][19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.reg_buf[15] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.i_regbuf[16]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[13][20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.reg_buf[16] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.i_regbuf[17]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[13][21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.reg_buf[17] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.i_regbuf[18]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[13][22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.reg_buf[18] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.i_regbuf[19]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[13][23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.reg_buf[19] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.i_regbuf[20]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[13][24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.reg_buf[20] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.i_regbuf[21]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[13][25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.reg_buf[21] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.i_regbuf[22]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[13][26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.reg_buf[22] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.i_regbuf[23]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[13][27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.reg_buf[23] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.i_regbuf[24]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[13][28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.reg_buf[24] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.i_regbuf[25]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[13][29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.reg_buf[25] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.i_regbuf[26]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[13][30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.reg_buf[26] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.i_regbuf[27]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[13][31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.reg_buf[27] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.i_regbuf[28]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[13][0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.reg_buf[28] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.i_regbuf[29]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[13][1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.reg_buf[29] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.i_regbuf[30]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[13][2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.reg_buf[30] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.i_regbuf[31]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[13][3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.reg_buf[31] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.i_regbuf[4]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[13][8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.reg_buf[4] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.i_regbuf[5]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[13][9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.reg_buf[5] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.i_regbuf[6]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[13][10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.reg_buf[6] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.i_regbuf[7]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[13][11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.reg_buf[7] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.i_regbuf[8]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[13][12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.reg_buf[8] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.i_regbuf[9]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[13][13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.genblk1.reg_buf[9] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.i_regbuf[10]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[14][14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.reg_buf[10] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.i_regbuf[11]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[14][15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.reg_buf[11] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.i_regbuf[12]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[14][16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.reg_buf[12] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.i_regbuf[13]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[14][17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.reg_buf[13] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.i_regbuf[14]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[14][18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.reg_buf[14] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.i_regbuf[15]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[14][19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.reg_buf[15] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.i_regbuf[16]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[14][20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.reg_buf[16] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.i_regbuf[17]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[14][21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.reg_buf[17] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.i_regbuf[18]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[14][22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.reg_buf[18] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.i_regbuf[19]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[14][23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.reg_buf[19] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.i_regbuf[20]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[14][24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.reg_buf[20] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.i_regbuf[21]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[14][25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.reg_buf[21] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.i_regbuf[22]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[14][26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.reg_buf[22] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.i_regbuf[23]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[14][27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.reg_buf[23] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.i_regbuf[24]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[14][28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.reg_buf[24] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.i_regbuf[25]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[14][29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.reg_buf[25] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.i_regbuf[26]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[14][30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.reg_buf[26] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.i_regbuf[27]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[14][31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.reg_buf[27] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.i_regbuf[28]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[14][0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.reg_buf[28] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.i_regbuf[29]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[14][1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.reg_buf[29] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.i_regbuf[30]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[14][2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.reg_buf[30] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.i_regbuf[31]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[14][3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.reg_buf[31] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.i_regbuf[4]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[14][8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.reg_buf[4] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.i_regbuf[5]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[14][9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.reg_buf[5] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.i_regbuf[6]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[14][10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.reg_buf[6] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.i_regbuf[7]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[14][11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.reg_buf[7] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.i_regbuf[8]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[14][12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.reg_buf[8] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.i_regbuf[9]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[14][13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.genblk1.reg_buf[9] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.i_regbuf[10]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[15][14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.reg_buf[10] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.i_regbuf[11]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[15][15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.reg_buf[11] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.i_regbuf[12]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[15][16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.reg_buf[12] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.i_regbuf[13]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[15][17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.reg_buf[13] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.i_regbuf[14]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[15][18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.reg_buf[14] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.i_regbuf[15]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[15][19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.reg_buf[15] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.i_regbuf[16]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[15][20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.reg_buf[16] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.i_regbuf[17]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[15][21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.reg_buf[17] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.i_regbuf[18]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[15][22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.reg_buf[18] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.i_regbuf[19]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[15][23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.reg_buf[19] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.i_regbuf[20]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[15][24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.reg_buf[20] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.i_regbuf[21]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[15][25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.reg_buf[21] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.i_regbuf[22]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[15][26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.reg_buf[22] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.i_regbuf[23]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[15][27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.reg_buf[23] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.i_regbuf[24]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[15][28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.reg_buf[24] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.i_regbuf[25]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[15][29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.reg_buf[25] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.i_regbuf[26]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[15][30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.reg_buf[26] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.i_regbuf[27]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[15][31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.reg_buf[27] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.i_regbuf[28]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[15][0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.reg_buf[28] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.i_regbuf[29]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[15][1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.reg_buf[29] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.i_regbuf[30]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[15][2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.reg_buf[30] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.i_regbuf[31]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[15][3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.reg_buf[31] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.i_regbuf[4]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[15][8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.reg_buf[4] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.i_regbuf[5]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[15][9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.reg_buf[5] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.i_regbuf[6]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[15][10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.reg_buf[6] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.i_regbuf[7]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[15][11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.reg_buf[7] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.i_regbuf[8]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[15][12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.reg_buf[8] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.i_regbuf[9]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[15][13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.genblk1.reg_buf[9] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.i_regbuf[10]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[1][14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.reg_buf[10] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.i_regbuf[11]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[1][15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.reg_buf[11] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.i_regbuf[12]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[1][16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.reg_buf[12] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.i_regbuf[13]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[1][17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.reg_buf[13] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.i_regbuf[14]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[1][18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.reg_buf[14] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.i_regbuf[15]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[1][19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.reg_buf[15] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.i_regbuf[16]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[1][20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.reg_buf[16] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.i_regbuf[17]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[1][21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.reg_buf[17] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.i_regbuf[18]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[1][22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.reg_buf[18] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.i_regbuf[19]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[1][23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.reg_buf[19] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.i_regbuf[20]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[1][24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.reg_buf[20] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.i_regbuf[21]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[1][25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.reg_buf[21] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.i_regbuf[22]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[1][26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.reg_buf[22] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.i_regbuf[23]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[1][27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.reg_buf[23] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.i_regbuf[24]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[1][28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.reg_buf[24] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.i_regbuf[25]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[1][29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.reg_buf[25] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.i_regbuf[26]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[1][30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.reg_buf[26] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.i_regbuf[27]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[1][31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.reg_buf[27] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.i_regbuf[28]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[1][0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.reg_buf[28] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.i_regbuf[29]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[1][1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.reg_buf[29] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.i_regbuf[30]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[1][2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.reg_buf[30] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.i_regbuf[31]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[1][3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.reg_buf[31] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.i_regbuf[4]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[1][8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.reg_buf[4] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.i_regbuf[5]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[1][9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.reg_buf[5] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.i_regbuf[6]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[1][10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.reg_buf[6] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.i_regbuf[7]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[1][11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.reg_buf[7] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.i_regbuf[8]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[1][12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.reg_buf[8] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.i_regbuf[9]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[1][13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.genblk1.reg_buf[9] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.i_regbuf[10]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[2][14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.reg_buf[10] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.i_regbuf[11]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[2][15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.reg_buf[11] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.i_regbuf[12]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[2][16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.reg_buf[12] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.i_regbuf[13]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[2][17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.reg_buf[13] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.i_regbuf[14]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[2][18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.reg_buf[14] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.i_regbuf[15]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[2][19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.reg_buf[15] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.i_regbuf[16]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[2][20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.reg_buf[16] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.i_regbuf[17]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[2][21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.reg_buf[17] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.i_regbuf[18]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[2][22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.reg_buf[18] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.i_regbuf[19]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[2][23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.reg_buf[19] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.i_regbuf[20]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[2][24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.reg_buf[20] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.i_regbuf[21]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[2][25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.reg_buf[21] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.i_regbuf[22]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[2][26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.reg_buf[22] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.i_regbuf[23]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[2][27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.reg_buf[23] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.i_regbuf[24]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[2][28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.reg_buf[24] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.i_regbuf[25]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[2][29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.reg_buf[25] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.i_regbuf[26]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[2][30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.reg_buf[26] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.i_regbuf[27]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[2][31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.reg_buf[27] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.i_regbuf[28]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[2][0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.reg_buf[28] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.i_regbuf[29]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[2][1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.reg_buf[29] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.i_regbuf[30]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[2][2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.reg_buf[30] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.i_regbuf[31]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[2][3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.reg_buf[31] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.i_regbuf[4]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[2][8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.reg_buf[4] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.i_regbuf[5]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[2][9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.reg_buf[5] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.i_regbuf[6]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[2][10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.reg_buf[6] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.i_regbuf[7]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[2][11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.reg_buf[7] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.i_regbuf[8]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[2][12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.reg_buf[8] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.i_regbuf[9]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[2][13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.genblk1.reg_buf[9] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.i_regbuf[10]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[5][14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.reg_buf[10] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.i_regbuf[11]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[5][15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.reg_buf[11] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.i_regbuf[12]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[5][16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.reg_buf[12] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.i_regbuf[13]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[5][17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.reg_buf[13] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.i_regbuf[14]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[5][18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.reg_buf[14] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.i_regbuf[15]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[5][19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.reg_buf[15] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.i_regbuf[16]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[5][20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.reg_buf[16] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.i_regbuf[17]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[5][21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.reg_buf[17] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.i_regbuf[18]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[5][22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.reg_buf[18] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.i_regbuf[19]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[5][23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.reg_buf[19] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.i_regbuf[20]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[5][24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.reg_buf[20] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.i_regbuf[21]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[5][25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.reg_buf[21] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.i_regbuf[22]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[5][26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.reg_buf[22] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.i_regbuf[23]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[5][27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.reg_buf[23] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.i_regbuf[24]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[5][28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.reg_buf[24] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.i_regbuf[25]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[5][29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.reg_buf[25] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.i_regbuf[26]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[5][30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.reg_buf[26] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.i_regbuf[27]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[5][31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.reg_buf[27] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.i_regbuf[28]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[5][0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.reg_buf[28] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.i_regbuf[29]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[5][1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.reg_buf[29] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.i_regbuf[30]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[5][2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.reg_buf[30] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.i_regbuf[31]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[5][3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.reg_buf[31] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.i_regbuf[4]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[5][8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.reg_buf[4] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.i_regbuf[5]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[5][9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.reg_buf[5] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.i_regbuf[6]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[5][10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.reg_buf[6] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.i_regbuf[7]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[5][11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.reg_buf[7] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.i_regbuf[8]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[5][12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.reg_buf[8] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.i_regbuf[9]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[5][13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.genblk1.reg_buf[9] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.i_regbuf[10]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[6][14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.reg_buf[10] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.i_regbuf[11]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[6][15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.reg_buf[11] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.i_regbuf[12]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[6][16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.reg_buf[12] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.i_regbuf[13]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[6][17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.reg_buf[13] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.i_regbuf[14]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[6][18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.reg_buf[14] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.i_regbuf[15]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[6][19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.reg_buf[15] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.i_regbuf[16]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[6][20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.reg_buf[16] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.i_regbuf[17]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[6][21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.reg_buf[17] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.i_regbuf[18]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[6][22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.reg_buf[18] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.i_regbuf[19]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[6][23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.reg_buf[19] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.i_regbuf[20]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[6][24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.reg_buf[20] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.i_regbuf[21]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[6][25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.reg_buf[21] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.i_regbuf[22]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[6][26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.reg_buf[22] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.i_regbuf[23]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[6][27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.reg_buf[23] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.i_regbuf[24]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[6][28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.reg_buf[24] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.i_regbuf[25]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[6][29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.reg_buf[25] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.i_regbuf[26]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[6][30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.reg_buf[26] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.i_regbuf[27]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[6][31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.reg_buf[27] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.i_regbuf[28]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[6][0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.reg_buf[28] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.i_regbuf[29]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[6][1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.reg_buf[29] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.i_regbuf[30]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[6][2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.reg_buf[30] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.i_regbuf[31]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[6][3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.reg_buf[31] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.i_regbuf[4]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[6][8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.reg_buf[4] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.i_regbuf[5]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[6][9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.reg_buf[5] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.i_regbuf[6]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[6][10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.reg_buf[6] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.i_regbuf[7]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[6][11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.reg_buf[7] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.i_regbuf[8]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[6][12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.reg_buf[8] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.i_regbuf[9]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[6][13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.genblk1.reg_buf[9] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.i_regbuf[10]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[7][14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.reg_buf[10] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.i_regbuf[11]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[7][15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.reg_buf[11] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.i_regbuf[12]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[7][16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.reg_buf[12] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.i_regbuf[13]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[7][17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.reg_buf[13] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.i_regbuf[14]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[7][18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.reg_buf[14] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.i_regbuf[15]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[7][19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.reg_buf[15] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.i_regbuf[16]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[7][20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.reg_buf[16] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.i_regbuf[17]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[7][21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.reg_buf[17] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.i_regbuf[18]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[7][22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.reg_buf[18] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.i_regbuf[19]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[7][23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.reg_buf[19] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.i_regbuf[20]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[7][24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.reg_buf[20] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.i_regbuf[21]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[7][25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.reg_buf[21] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.i_regbuf[22]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[7][26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.reg_buf[22] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.i_regbuf[23]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[7][27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.reg_buf[23] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.i_regbuf[24]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[7][28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.reg_buf[24] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.i_regbuf[25]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[7][29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.reg_buf[25] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.i_regbuf[26]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[7][30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.reg_buf[26] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.i_regbuf[27]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[7][31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.reg_buf[27] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.i_regbuf[28]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[7][0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.reg_buf[28] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.i_regbuf[29]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[7][1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.reg_buf[29] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.i_regbuf[30]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[7][2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.reg_buf[30] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.i_regbuf[31]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[7][3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.reg_buf[31] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.i_regbuf[4]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[7][8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.reg_buf[4] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.i_regbuf[5]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[7][9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.reg_buf[5] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.i_regbuf[6]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[7][10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.reg_buf[6] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.i_regbuf[7]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[7][11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.reg_buf[7] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.i_regbuf[8]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[7][12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.reg_buf[8] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.i_regbuf[9]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[7][13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.genblk1.reg_buf[9] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.i_regbuf[10]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[8][14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.reg_buf[10] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.i_regbuf[11]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[8][15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.reg_buf[11] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.i_regbuf[12]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[8][16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.reg_buf[12] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.i_regbuf[13]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[8][17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.reg_buf[13] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.i_regbuf[14]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[8][18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.reg_buf[14] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.i_regbuf[15]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[8][19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.reg_buf[15] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.i_regbuf[16]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[8][20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.reg_buf[16] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.i_regbuf[17]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[8][21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.reg_buf[17] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.i_regbuf[18]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[8][22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.reg_buf[18] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.i_regbuf[19]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[8][23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.reg_buf[19] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.i_regbuf[20]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[8][24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.reg_buf[20] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.i_regbuf[21]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[8][25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.reg_buf[21] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.i_regbuf[22]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[8][26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.reg_buf[22] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.i_regbuf[23]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[8][27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.reg_buf[23] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.i_regbuf[24]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[8][28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.reg_buf[24] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.i_regbuf[25]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[8][29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.reg_buf[25] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.i_regbuf[26]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[8][30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.reg_buf[26] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.i_regbuf[27]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[8][31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.reg_buf[27] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.i_regbuf[28]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[8][0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.reg_buf[28] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.i_regbuf[29]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[8][1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.reg_buf[29] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.i_regbuf[30]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[8][2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.reg_buf[30] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.i_regbuf[31]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[8][3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.reg_buf[31] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.i_regbuf[4]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[8][8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.reg_buf[4] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.i_regbuf[5]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[8][9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.reg_buf[5] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.i_regbuf[6]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[8][10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.reg_buf[6] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.i_regbuf[7]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[8][11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.reg_buf[7] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.i_regbuf[8]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[8][12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.reg_buf[8] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.i_regbuf[9]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[8][13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.genblk1.reg_buf[9] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.i_regbuf[10]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[9][14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.reg_buf[10] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.i_regbuf[11]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[9][15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.reg_buf[11] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.i_regbuf[12]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[9][16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.reg_buf[12] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.i_regbuf[13]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[9][17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.reg_buf[13] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.i_regbuf[14]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[9][18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.reg_buf[14] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.i_regbuf[15]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[9][19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.reg_buf[15] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.i_regbuf[16]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[9][20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.reg_buf[16] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.i_regbuf[17]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[9][21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.reg_buf[17] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.i_regbuf[18]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[9][22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.reg_buf[18] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.i_regbuf[19]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[9][23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.reg_buf[19] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.i_regbuf[20]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[9][24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.reg_buf[20] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.i_regbuf[21]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[9][25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.reg_buf[21] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.i_regbuf[22]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[9][26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.reg_buf[22] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.i_regbuf[23]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[9][27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.reg_buf[23] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.i_regbuf[24]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[9][28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.reg_buf[24] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.i_regbuf[25]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[9][29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.reg_buf[25] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.i_regbuf[26]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[9][30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.reg_buf[26] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.i_regbuf[27]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[9][31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.reg_buf[27] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.i_regbuf[28]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[9][0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.reg_buf[28] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.i_regbuf[29]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[9][1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.reg_buf[29] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.i_regbuf[30]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[9][2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.reg_buf[30] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.i_regbuf[31]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[9][3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.reg_buf[31] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.i_regbuf[4]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[9][8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.reg_buf[4] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.i_regbuf[5]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[9][9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.reg_buf[5] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.i_regbuf[6]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[9][10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.reg_buf[6] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.i_regbuf[7]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[9][11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.reg_buf[7] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.i_regbuf[8]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[9][12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.reg_buf[8] ));
 sky130_fd_sc_hd__dlygate4sd3_1 \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.i_regbuf[9]  (.A(\i_tinyqv.cpu.i_core.i_registers.registers[9][13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.genblk1.reg_buf[9] ));
 sky130_fd_sc_hd__buf_2 input1 (.A(rst_n),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net1));
 sky130_fd_sc_hd__buf_1 input10 (.A(uio_in[1]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net10));
 sky130_fd_sc_hd__buf_1 input11 (.A(uio_in[2]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net11));
 sky130_fd_sc_hd__buf_1 input12 (.A(uio_in[4]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net12));
 sky130_fd_sc_hd__buf_1 input13 (.A(uio_in[5]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net13));
 sky130_fd_sc_hd__buf_1 input2 (.A(ui_in[0]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(ui_in[1]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(ui_in[2]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net4));
 sky130_fd_sc_hd__buf_2 input5 (.A(ui_in[3]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_2 input6 (.A(ui_in[4]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net6));
 sky130_fd_sc_hd__dlymetal6s2s_1 input7 (.A(ui_in[5]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net7));
 sky130_fd_sc_hd__buf_1 input8 (.A(ui_in[6]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net8));
 sky130_fd_sc_hd__buf_1 input9 (.A(ui_in[7]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_1 max_cap1 (.A(_0683_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net320));
 sky130_fd_sc_hd__buf_2 max_cap14 (.A(_1003_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net14));
 sky130_fd_sc_hd__buf_1 max_cap15 (.A(_0943_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_2 max_cap18 (.A(_2089_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net18));
 sky130_fd_sc_hd__buf_1 max_cap19 (.A(_0948_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net19));
 sky130_fd_sc_hd__buf_1 max_cap2 (.A(_0634_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net321));
 sky130_fd_sc_hd__clkbuf_1 max_cap21 (.A(net22),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_1 max_cap23 (.A(_0714_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_2 max_cap24 (.A(_0683_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net24));
 sky130_fd_sc_hd__buf_1 max_cap26 (.A(_0638_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net26));
 sky130_fd_sc_hd__buf_1 max_cap27 (.A(_0634_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_1 rebuffer1 (.A(\i_tinyqv.cpu.i_core.i_registers.rs1[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_1 rebuffer10 (.A(net38),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net39));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer11 (.A(_1339_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net325));
 sky130_fd_sc_hd__buf_1 rebuffer12 (.A(_0652_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_1 rebuffer13 (.A(net41),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_1 rebuffer14 (.A(_0652_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_1 rebuffer15 (.A(net20),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net44));
 sky130_fd_sc_hd__buf_1 rebuffer16 (.A(net44),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_1 rebuffer17 (.A(_0643_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net46));
 sky130_fd_sc_hd__buf_1 rebuffer18 (.A(_0643_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_1 rebuffer19 (.A(net47),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net48));
 sky130_fd_sc_hd__buf_2 rebuffer2 (.A(_1546_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net31));
 sky130_fd_sc_hd__buf_1 rebuffer20 (.A(_0687_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net49));
 sky130_fd_sc_hd__buf_1 rebuffer21 (.A(net49),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_1 rebuffer22 (.A(\i_tinyqv.cpu.i_core.i_registers.rs1[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_1 rebuffer23 (.A(\i_tinyqv.cpu.i_core.i_registers.rs1[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_1 rebuffer24 (.A(\i_tinyqv.cpu.i_core.i_registers.rs1[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_1 rebuffer25 (.A(_0642_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_1 rebuffer26 (.A(_0649_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net55));
 sky130_fd_sc_hd__clkbuf_1 rebuffer27 (.A(\i_tinyqv.cpu.i_core.i_registers.rs1[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net56));
 sky130_fd_sc_hd__clkbuf_1 rebuffer28 (.A(_0645_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net57));
 sky130_fd_sc_hd__clkbuf_1 rebuffer29 (.A(_0645_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net58));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer3 (.A(_1412_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net322));
 sky130_fd_sc_hd__clkbuf_1 rebuffer30 (.A(net22),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net59));
 sky130_fd_sc_hd__clkbuf_1 rebuffer32 (.A(_0668_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net61));
 sky130_fd_sc_hd__buf_1 rebuffer33 (.A(_0628_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net62));
 sky130_fd_sc_hd__clkbuf_1 rebuffer34 (.A(net62),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net63));
 sky130_fd_sc_hd__buf_1 rebuffer35 (.A(_0740_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net64));
 sky130_fd_sc_hd__clkbuf_1 rebuffer36 (.A(_0740_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net65));
 sky130_fd_sc_hd__clkbuf_2 rebuffer37 (.A(_0762_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net66));
 sky130_fd_sc_hd__clkbuf_1 rebuffer38 (.A(net66),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net67));
 sky130_fd_sc_hd__clkbuf_1 rebuffer39 (.A(_0762_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net68));
 sky130_fd_sc_hd__clkbuf_1 rebuffer4 (.A(_1397_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_1 rebuffer41 (.A(\i_tinyqv.cpu.i_core.i_registers.rs1[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net70));
 sky130_fd_sc_hd__buf_1 rebuffer42 (.A(net323),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net71));
 sky130_fd_sc_hd__clkbuf_1 rebuffer43 (.A(net71),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net72));
 sky130_fd_sc_hd__clkbuf_1 rebuffer44 (.A(net71),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net73));
 sky130_fd_sc_hd__buf_1 rebuffer45 (.A(_0631_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net74));
 sky130_fd_sc_hd__clkbuf_1 rebuffer46 (.A(net74),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net75));
 sky130_fd_sc_hd__buf_1 rebuffer47 (.A(_0793_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net76));
 sky130_fd_sc_hd__buf_1 rebuffer48 (.A(_0720_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net77));
 sky130_fd_sc_hd__clkbuf_1 rebuffer49 (.A(net77),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net78));
 sky130_fd_sc_hd__clkbuf_1 rebuffer5 (.A(net36),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_1 rebuffer50 (.A(net77),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net79));
 sky130_fd_sc_hd__clkbuf_1 rebuffer51 (.A(_0655_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net80));
 sky130_fd_sc_hd__buf_1 rebuffer52 (.A(_0798_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net81));
 sky130_fd_sc_hd__clkbuf_1 rebuffer53 (.A(_1583_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net82));
 sky130_fd_sc_hd__clkbuf_1 rebuffer54 (.A(_0633_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net83));
 sky130_fd_sc_hd__clkbuf_1 rebuffer55 (.A(_0633_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net84));
 sky130_fd_sc_hd__clkbuf_2 rebuffer56 (.A(\i_tinyqv.cpu.pc[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net85));
 sky130_fd_sc_hd__buf_1 rebuffer57 (.A(_0799_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net86));
 sky130_fd_sc_hd__clkbuf_1 rebuffer58 (.A(\i_tinyqv.cpu.i_core.i_registers.rs1[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net87));
 sky130_fd_sc_hd__clkbuf_1 rebuffer59 (.A(_0649_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net88));
 sky130_fd_sc_hd__clkbuf_1 rebuffer6 (.A(net36),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net35));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer7 (.A(_0651_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net323));
 sky130_fd_sc_hd__buf_6 rebuffer8 (.A(\i_tinyqv.cpu.i_core.i_registers.rs2[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net37));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer9 (.A(\i_tinyqv.cpu.i_core.i_registers.rs2[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net38));
 sky130_fd_sc_hd__buf_1 split31 (.A(\i_tinyqv.cpu.pc[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net60));
 sky130_fd_sc_hd__buf_2 split40 (.A(\i_tinyqv.cpu.alu_op[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net69));
 sky130_fd_sc_hd__buf_4 wire16 (.A(_0808_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net16));
 sky130_fd_sc_hd__buf_1 wire17 (.A(_2241_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net17));
 sky130_fd_sc_hd__buf_1 wire20 (.A(_0736_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net20));
 sky130_fd_sc_hd__buf_2 wire22 (.A(_0719_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net22));
 sky130_fd_sc_hd__buf_1 wire25 (.A(_0671_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net25));
 sky130_fd_sc_hd__buf_2 wire28 (.A(_0972_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net28));
endmodule
