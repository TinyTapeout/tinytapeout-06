VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_emilian_rf_playground
  CLASS BLOCK ;
  FOREIGN tt_um_emilian_rf_playground ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 154.870 224.760 155.170 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 158.550 224.760 158.850 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 151.190 224.760 151.490 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.000000 ;
    ANTENNADIFFAREA 1.740000 ;
    PORT
      LAYER met4 ;
        RECT 156.560 0.000 157.160 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.160000 ;
    PORT
      LAYER met4 ;
        RECT 134.480 0.000 135.080 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.000000 ;
    PORT
      LAYER met4 ;
        RECT 112.400 0.000 113.000 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 90.320 0.000 90.920 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 68.240 0.000 68.840 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 46.160 0.000 46.760 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 24.080 0.000 24.680 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 2.000 0.000 2.600 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 147.510 224.760 147.810 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 140.150 224.760 140.450 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 136.470 224.760 136.770 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 129.110 224.760 129.410 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 125.430 224.760 125.730 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.070 224.760 118.370 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 114.390 224.760 114.690 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.030 224.760 107.330 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 103.350 224.760 103.650 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 95.990 224.760 96.290 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 92.310 224.760 92.610 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 137.678391 ;
    PORT
      LAYER met4 ;
        RECT 29.750 224.760 30.050 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 26.070 224.760 26.370 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 22.390 224.760 22.690 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 18.710 224.760 19.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 15.030 224.760 15.330 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 11.350 224.760 11.650 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 7.670 224.760 7.970 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 3.990 224.760 4.290 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 137.678391 ;
    PORT
      LAYER met4 ;
        RECT 59.190 224.760 59.490 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 137.678391 ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 137.678391 ;
    PORT
      LAYER met4 ;
        RECT 51.830 224.760 52.130 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 137.678391 ;
    PORT
      LAYER met4 ;
        RECT 48.150 224.760 48.450 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 40.790 224.760 41.090 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 37.110 224.760 37.410 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 84.950 224.760 85.250 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 81.270 224.760 81.570 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 73.910 224.760 74.210 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 70.230 224.760 70.530 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 62.870 224.760 63.170 225.760 ;
    END
  END uo_out[7]
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 2.500 220.760 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 49.000 5.000 50.500 220.760 ;
    END
  END VGND
  OBS
      LAYER pwell ;
        RECT 132.130 68.460 143.030 69.460 ;
        RECT 128.130 68.220 143.030 68.460 ;
        RECT 128.080 65.260 143.030 68.220 ;
        RECT 128.130 65.160 143.030 65.260 ;
      LAYER nwell ;
        RECT 125.440 64.410 131.630 64.420 ;
        RECT 125.430 58.460 131.630 64.410 ;
      LAYER pwell ;
        RECT 132.230 61.760 143.030 65.160 ;
      LAYER nwell ;
        RECT 143.630 62.510 149.830 68.460 ;
        RECT 143.630 62.500 149.820 62.510 ;
      LAYER pwell ;
        RECT 132.230 61.660 147.130 61.760 ;
        RECT 132.230 58.700 147.180 61.660 ;
        RECT 132.230 58.460 147.130 58.700 ;
        RECT 132.230 57.460 143.130 58.460 ;
        RECT 132.130 56.460 143.030 57.460 ;
        RECT 128.130 56.220 143.030 56.460 ;
        RECT 128.080 53.260 143.030 56.220 ;
        RECT 128.130 53.160 143.030 53.260 ;
      LAYER nwell ;
        RECT 125.440 52.410 131.630 52.420 ;
        RECT 125.430 46.460 131.630 52.410 ;
      LAYER pwell ;
        RECT 132.230 49.760 143.030 53.160 ;
      LAYER nwell ;
        RECT 143.630 50.510 149.830 56.460 ;
        RECT 143.630 50.500 149.820 50.510 ;
      LAYER pwell ;
        RECT 132.230 49.660 147.130 49.760 ;
        RECT 132.230 46.700 147.180 49.660 ;
        RECT 132.230 46.460 147.130 46.700 ;
        RECT 132.230 45.460 143.130 46.460 ;
        RECT 132.130 44.460 143.030 45.460 ;
        RECT 128.130 44.220 143.030 44.460 ;
        RECT 128.080 41.260 143.030 44.220 ;
        RECT 128.130 41.160 143.030 41.260 ;
      LAYER nwell ;
        RECT 125.440 40.410 131.630 40.420 ;
        RECT 125.430 34.460 131.630 40.410 ;
      LAYER pwell ;
        RECT 132.230 37.760 143.030 41.160 ;
      LAYER nwell ;
        RECT 143.630 38.510 149.830 44.460 ;
        RECT 143.630 38.500 149.820 38.510 ;
      LAYER pwell ;
        RECT 132.230 37.660 147.130 37.760 ;
        RECT 132.230 34.700 147.180 37.660 ;
        RECT 132.230 34.460 147.130 34.700 ;
        RECT 132.230 33.460 143.130 34.460 ;
        RECT 132.130 32.460 143.030 33.460 ;
        RECT 128.130 32.220 143.030 32.460 ;
        RECT 128.080 29.260 143.030 32.220 ;
        RECT 128.130 29.160 143.030 29.260 ;
      LAYER nwell ;
        RECT 125.440 28.410 131.630 28.420 ;
        RECT 125.430 22.460 131.630 28.410 ;
      LAYER pwell ;
        RECT 132.230 25.760 143.030 29.160 ;
      LAYER nwell ;
        RECT 143.630 26.510 149.830 32.460 ;
        RECT 143.630 26.500 149.820 26.510 ;
      LAYER pwell ;
        RECT 132.230 25.660 147.130 25.760 ;
        RECT 132.230 22.700 147.180 25.660 ;
        RECT 132.230 22.460 147.130 22.700 ;
        RECT 132.230 21.460 143.130 22.460 ;
      LAYER nwell ;
        RECT 135.130 19.470 143.330 19.560 ;
        RECT 131.640 19.360 143.380 19.470 ;
        RECT 131.640 16.560 143.430 19.360 ;
        RECT 131.640 16.510 143.380 16.560 ;
      LAYER li1 ;
        RECT 121.730 20.060 123.830 74.060 ;
        RECT 124.630 70.460 150.630 72.460 ;
        RECT 124.630 69.460 126.130 70.460 ;
        RECT 149.130 69.460 150.630 70.460 ;
        RECT 124.630 68.390 126.380 69.460 ;
        RECT 132.130 68.960 143.130 69.460 ;
        RECT 148.880 69.260 150.630 69.460 ;
        RECT 132.130 68.660 139.030 68.960 ;
        RECT 139.730 68.710 141.230 68.960 ;
        RECT 132.130 68.460 133.030 68.660 ;
        RECT 124.630 64.560 127.750 68.390 ;
        RECT 128.130 67.860 133.030 68.460 ;
        RECT 133.560 68.200 135.600 68.370 ;
        RECT 128.130 65.660 128.430 67.860 ;
        RECT 129.110 67.300 131.150 67.470 ;
        RECT 128.770 66.240 128.940 67.240 ;
        RECT 131.320 66.240 131.490 67.240 ;
        RECT 131.730 66.560 133.030 67.860 ;
        RECT 133.220 67.140 133.390 68.140 ;
        RECT 134.030 67.080 135.530 67.160 ;
        RECT 135.770 67.140 135.940 68.140 ;
        RECT 133.560 66.910 135.600 67.080 ;
        RECT 134.030 66.560 135.530 66.910 ;
        RECT 136.230 66.860 139.030 68.660 ;
        RECT 139.660 68.540 141.700 68.710 ;
        RECT 139.320 68.260 139.490 68.480 ;
        RECT 141.870 68.260 142.040 68.480 ;
        RECT 139.320 67.480 142.040 68.260 ;
        RECT 139.330 67.260 142.030 67.480 ;
        RECT 139.660 67.250 141.700 67.260 ;
        RECT 142.230 66.860 143.130 68.960 ;
        RECT 136.230 66.560 143.130 66.860 ;
        RECT 129.110 66.010 131.150 66.180 ;
        RECT 131.730 66.160 143.130 66.560 ;
        RECT 131.730 65.870 139.030 66.160 ;
        RECT 131.730 65.660 133.030 65.870 ;
        RECT 128.130 65.160 133.030 65.660 ;
        RECT 133.580 65.470 135.580 65.610 ;
        RECT 133.560 65.300 135.600 65.470 ;
        RECT 124.630 63.960 131.530 64.560 ;
        RECT 124.630 61.860 125.930 63.960 ;
        RECT 126.515 63.610 130.555 63.670 ;
        RECT 126.230 63.440 130.880 63.610 ;
        RECT 126.130 63.060 130.940 63.440 ;
        RECT 126.130 62.440 126.300 63.060 ;
        RECT 130.770 62.440 130.940 63.060 ;
        RECT 126.515 62.210 130.555 62.380 ;
        RECT 126.730 61.860 130.380 62.210 ;
        RECT 131.230 61.860 131.530 63.960 ;
        RECT 124.630 60.960 131.530 61.860 ;
        RECT 124.630 58.860 125.930 60.960 ;
        RECT 126.730 60.670 130.380 60.960 ;
        RECT 126.515 60.500 130.555 60.670 ;
        RECT 126.130 59.440 126.300 60.440 ;
        RECT 130.770 59.440 130.940 60.440 ;
        RECT 126.515 59.210 130.555 59.380 ;
        RECT 131.230 58.860 131.530 60.960 ;
        RECT 124.630 57.660 131.530 58.860 ;
        RECT 132.130 63.660 133.030 65.160 ;
        RECT 133.220 64.240 133.390 65.240 ;
        RECT 134.030 64.180 135.530 64.260 ;
        RECT 135.770 64.240 135.940 65.240 ;
        RECT 133.560 64.010 135.600 64.180 ;
        RECT 134.030 63.660 135.530 64.010 ;
        RECT 136.230 63.960 139.030 65.870 ;
        RECT 139.730 65.810 141.230 66.160 ;
        RECT 139.660 65.640 141.700 65.810 ;
        RECT 139.320 65.360 139.490 65.580 ;
        RECT 141.870 65.360 142.040 65.580 ;
        RECT 139.320 64.580 142.040 65.360 ;
        RECT 139.330 64.360 142.030 64.580 ;
        RECT 139.660 64.350 141.700 64.360 ;
        RECT 142.230 63.960 143.130 66.160 ;
        RECT 136.230 63.660 143.130 63.960 ;
        RECT 132.130 63.260 143.130 63.660 ;
        RECT 132.130 62.960 139.030 63.260 ;
        RECT 132.130 60.760 133.030 62.960 ;
        RECT 133.560 62.560 135.600 62.570 ;
        RECT 133.230 62.340 135.930 62.560 ;
        RECT 133.220 61.560 135.940 62.340 ;
        RECT 133.220 61.340 133.390 61.560 ;
        RECT 135.770 61.340 135.940 61.560 ;
        RECT 133.560 61.110 135.600 61.280 ;
        RECT 134.030 60.760 135.530 61.110 ;
        RECT 136.230 61.050 139.030 62.960 ;
        RECT 139.730 62.910 141.230 63.260 ;
        RECT 139.660 62.740 141.700 62.910 ;
        RECT 139.320 61.680 139.490 62.680 ;
        RECT 139.730 62.660 141.230 62.740 ;
        RECT 141.870 61.680 142.040 62.680 ;
        RECT 142.230 61.760 143.130 63.260 ;
        RECT 143.730 68.060 150.630 69.260 ;
        RECT 143.730 65.960 144.030 68.060 ;
        RECT 144.705 67.540 148.745 67.710 ;
        RECT 144.320 66.480 144.490 67.480 ;
        RECT 148.960 66.480 149.130 67.480 ;
        RECT 144.705 66.250 148.745 66.420 ;
        RECT 144.880 65.960 148.530 66.250 ;
        RECT 149.330 65.960 150.630 68.060 ;
        RECT 143.730 65.060 150.630 65.960 ;
        RECT 143.730 62.960 144.030 65.060 ;
        RECT 144.880 64.710 148.530 65.060 ;
        RECT 144.705 64.540 148.745 64.710 ;
        RECT 144.320 63.860 144.490 64.480 ;
        RECT 148.960 63.860 149.130 64.480 ;
        RECT 144.320 63.480 149.130 63.860 ;
        RECT 144.380 63.310 149.030 63.480 ;
        RECT 144.705 63.250 148.745 63.310 ;
        RECT 149.330 62.960 150.630 65.060 ;
        RECT 143.730 62.360 150.630 62.960 ;
        RECT 139.660 61.450 141.700 61.620 ;
        RECT 139.680 61.310 141.680 61.450 ;
        RECT 142.230 61.260 147.130 61.760 ;
        RECT 142.230 61.050 143.530 61.260 ;
        RECT 136.230 60.760 143.530 61.050 ;
        RECT 132.130 60.360 143.530 60.760 ;
        RECT 144.110 60.740 146.150 60.910 ;
        RECT 132.130 60.060 139.030 60.360 ;
        RECT 132.130 57.960 133.030 60.060 ;
        RECT 133.560 59.660 135.600 59.670 ;
        RECT 133.230 59.440 135.930 59.660 ;
        RECT 133.220 58.660 135.940 59.440 ;
        RECT 133.220 58.440 133.390 58.660 ;
        RECT 135.770 58.440 135.940 58.660 ;
        RECT 133.560 58.210 135.600 58.380 ;
        RECT 136.230 58.260 139.030 60.060 ;
        RECT 139.730 60.010 141.230 60.360 ;
        RECT 139.660 59.840 141.700 60.010 ;
        RECT 139.320 58.780 139.490 59.780 ;
        RECT 139.730 59.760 141.230 59.840 ;
        RECT 141.870 58.780 142.040 59.780 ;
        RECT 142.230 59.060 143.530 60.360 ;
        RECT 143.770 59.680 143.940 60.680 ;
        RECT 146.320 59.680 146.490 60.680 ;
        RECT 144.110 59.450 146.150 59.620 ;
        RECT 146.830 59.060 147.130 61.260 ;
        RECT 139.660 58.550 141.700 58.720 ;
        RECT 142.230 58.460 147.130 59.060 ;
        RECT 147.510 58.530 150.630 62.360 ;
        RECT 142.230 58.260 143.130 58.460 ;
        RECT 134.030 57.960 135.530 58.210 ;
        RECT 136.230 57.960 143.130 58.260 ;
        RECT 124.630 56.390 126.380 57.660 ;
        RECT 132.130 56.960 143.130 57.960 ;
        RECT 148.880 57.260 150.630 58.530 ;
        RECT 132.130 56.660 139.030 56.960 ;
        RECT 139.730 56.710 141.230 56.960 ;
        RECT 132.130 56.460 133.030 56.660 ;
        RECT 124.630 52.560 127.750 56.390 ;
        RECT 128.130 55.860 133.030 56.460 ;
        RECT 133.560 56.200 135.600 56.370 ;
        RECT 128.130 53.660 128.430 55.860 ;
        RECT 129.110 55.300 131.150 55.470 ;
        RECT 128.770 54.240 128.940 55.240 ;
        RECT 131.320 54.240 131.490 55.240 ;
        RECT 131.730 54.560 133.030 55.860 ;
        RECT 133.220 55.140 133.390 56.140 ;
        RECT 134.030 55.080 135.530 55.160 ;
        RECT 135.770 55.140 135.940 56.140 ;
        RECT 133.560 54.910 135.600 55.080 ;
        RECT 134.030 54.560 135.530 54.910 ;
        RECT 136.230 54.860 139.030 56.660 ;
        RECT 139.660 56.540 141.700 56.710 ;
        RECT 139.320 56.260 139.490 56.480 ;
        RECT 141.870 56.260 142.040 56.480 ;
        RECT 139.320 55.480 142.040 56.260 ;
        RECT 139.330 55.260 142.030 55.480 ;
        RECT 139.660 55.250 141.700 55.260 ;
        RECT 142.230 54.860 143.130 56.960 ;
        RECT 136.230 54.560 143.130 54.860 ;
        RECT 129.110 54.010 131.150 54.180 ;
        RECT 131.730 54.160 143.130 54.560 ;
        RECT 131.730 53.870 139.030 54.160 ;
        RECT 131.730 53.660 133.030 53.870 ;
        RECT 128.130 53.160 133.030 53.660 ;
        RECT 133.580 53.470 135.580 53.610 ;
        RECT 133.560 53.300 135.600 53.470 ;
        RECT 124.630 51.960 131.530 52.560 ;
        RECT 124.630 49.860 125.930 51.960 ;
        RECT 126.515 51.610 130.555 51.670 ;
        RECT 126.230 51.440 130.880 51.610 ;
        RECT 126.130 51.060 130.940 51.440 ;
        RECT 126.130 50.440 126.300 51.060 ;
        RECT 130.770 50.440 130.940 51.060 ;
        RECT 126.515 50.210 130.555 50.380 ;
        RECT 126.730 49.860 130.380 50.210 ;
        RECT 131.230 49.860 131.530 51.960 ;
        RECT 124.630 48.960 131.530 49.860 ;
        RECT 124.630 46.860 125.930 48.960 ;
        RECT 126.730 48.670 130.380 48.960 ;
        RECT 126.515 48.500 130.555 48.670 ;
        RECT 126.130 47.440 126.300 48.440 ;
        RECT 130.770 47.440 130.940 48.440 ;
        RECT 126.515 47.210 130.555 47.380 ;
        RECT 131.230 46.860 131.530 48.960 ;
        RECT 124.630 45.660 131.530 46.860 ;
        RECT 132.130 51.660 133.030 53.160 ;
        RECT 133.220 52.240 133.390 53.240 ;
        RECT 134.030 52.180 135.530 52.260 ;
        RECT 135.770 52.240 135.940 53.240 ;
        RECT 133.560 52.010 135.600 52.180 ;
        RECT 134.030 51.660 135.530 52.010 ;
        RECT 136.230 51.960 139.030 53.870 ;
        RECT 139.730 53.810 141.230 54.160 ;
        RECT 139.660 53.640 141.700 53.810 ;
        RECT 139.320 53.360 139.490 53.580 ;
        RECT 141.870 53.360 142.040 53.580 ;
        RECT 139.320 52.580 142.040 53.360 ;
        RECT 139.330 52.360 142.030 52.580 ;
        RECT 139.660 52.350 141.700 52.360 ;
        RECT 142.230 51.960 143.130 54.160 ;
        RECT 136.230 51.660 143.130 51.960 ;
        RECT 132.130 51.260 143.130 51.660 ;
        RECT 132.130 50.960 139.030 51.260 ;
        RECT 132.130 48.760 133.030 50.960 ;
        RECT 133.560 50.560 135.600 50.570 ;
        RECT 133.230 50.340 135.930 50.560 ;
        RECT 133.220 49.560 135.940 50.340 ;
        RECT 133.220 49.340 133.390 49.560 ;
        RECT 135.770 49.340 135.940 49.560 ;
        RECT 133.560 49.110 135.600 49.280 ;
        RECT 134.030 48.760 135.530 49.110 ;
        RECT 136.230 49.050 139.030 50.960 ;
        RECT 139.730 50.910 141.230 51.260 ;
        RECT 139.660 50.740 141.700 50.910 ;
        RECT 139.320 49.680 139.490 50.680 ;
        RECT 139.730 50.660 141.230 50.740 ;
        RECT 141.870 49.680 142.040 50.680 ;
        RECT 142.230 49.760 143.130 51.260 ;
        RECT 143.730 56.060 150.630 57.260 ;
        RECT 143.730 53.960 144.030 56.060 ;
        RECT 144.705 55.540 148.745 55.710 ;
        RECT 144.320 54.480 144.490 55.480 ;
        RECT 148.960 54.480 149.130 55.480 ;
        RECT 144.705 54.250 148.745 54.420 ;
        RECT 144.880 53.960 148.530 54.250 ;
        RECT 149.330 53.960 150.630 56.060 ;
        RECT 143.730 53.060 150.630 53.960 ;
        RECT 143.730 50.960 144.030 53.060 ;
        RECT 144.880 52.710 148.530 53.060 ;
        RECT 144.705 52.540 148.745 52.710 ;
        RECT 144.320 51.860 144.490 52.480 ;
        RECT 148.960 51.860 149.130 52.480 ;
        RECT 144.320 51.480 149.130 51.860 ;
        RECT 144.380 51.310 149.030 51.480 ;
        RECT 144.705 51.250 148.745 51.310 ;
        RECT 149.330 50.960 150.630 53.060 ;
        RECT 143.730 50.360 150.630 50.960 ;
        RECT 139.660 49.450 141.700 49.620 ;
        RECT 139.680 49.310 141.680 49.450 ;
        RECT 142.230 49.260 147.130 49.760 ;
        RECT 142.230 49.050 143.530 49.260 ;
        RECT 136.230 48.760 143.530 49.050 ;
        RECT 132.130 48.360 143.530 48.760 ;
        RECT 144.110 48.740 146.150 48.910 ;
        RECT 132.130 48.060 139.030 48.360 ;
        RECT 132.130 45.960 133.030 48.060 ;
        RECT 133.560 47.660 135.600 47.670 ;
        RECT 133.230 47.440 135.930 47.660 ;
        RECT 133.220 46.660 135.940 47.440 ;
        RECT 133.220 46.440 133.390 46.660 ;
        RECT 135.770 46.440 135.940 46.660 ;
        RECT 133.560 46.210 135.600 46.380 ;
        RECT 136.230 46.260 139.030 48.060 ;
        RECT 139.730 48.010 141.230 48.360 ;
        RECT 139.660 47.840 141.700 48.010 ;
        RECT 139.320 46.780 139.490 47.780 ;
        RECT 139.730 47.760 141.230 47.840 ;
        RECT 141.870 46.780 142.040 47.780 ;
        RECT 142.230 47.060 143.530 48.360 ;
        RECT 143.770 47.680 143.940 48.680 ;
        RECT 146.320 47.680 146.490 48.680 ;
        RECT 144.110 47.450 146.150 47.620 ;
        RECT 146.830 47.060 147.130 49.260 ;
        RECT 139.660 46.550 141.700 46.720 ;
        RECT 142.230 46.460 147.130 47.060 ;
        RECT 147.510 46.530 150.630 50.360 ;
        RECT 142.230 46.260 143.130 46.460 ;
        RECT 134.030 45.960 135.530 46.210 ;
        RECT 136.230 45.960 143.130 46.260 ;
        RECT 124.630 44.390 126.380 45.660 ;
        RECT 132.130 44.960 143.130 45.960 ;
        RECT 148.880 45.260 150.630 46.530 ;
        RECT 132.130 44.660 139.030 44.960 ;
        RECT 139.730 44.710 141.230 44.960 ;
        RECT 132.130 44.460 133.030 44.660 ;
        RECT 124.630 40.560 127.750 44.390 ;
        RECT 128.130 43.860 133.030 44.460 ;
        RECT 133.560 44.200 135.600 44.370 ;
        RECT 128.130 41.660 128.430 43.860 ;
        RECT 129.110 43.300 131.150 43.470 ;
        RECT 128.770 42.240 128.940 43.240 ;
        RECT 131.320 42.240 131.490 43.240 ;
        RECT 131.730 42.560 133.030 43.860 ;
        RECT 133.220 43.140 133.390 44.140 ;
        RECT 134.030 43.080 135.530 43.160 ;
        RECT 135.770 43.140 135.940 44.140 ;
        RECT 133.560 42.910 135.600 43.080 ;
        RECT 134.030 42.560 135.530 42.910 ;
        RECT 136.230 42.860 139.030 44.660 ;
        RECT 139.660 44.540 141.700 44.710 ;
        RECT 139.320 44.260 139.490 44.480 ;
        RECT 141.870 44.260 142.040 44.480 ;
        RECT 139.320 43.480 142.040 44.260 ;
        RECT 139.330 43.260 142.030 43.480 ;
        RECT 139.660 43.250 141.700 43.260 ;
        RECT 142.230 42.860 143.130 44.960 ;
        RECT 136.230 42.560 143.130 42.860 ;
        RECT 129.110 42.010 131.150 42.180 ;
        RECT 131.730 42.160 143.130 42.560 ;
        RECT 131.730 41.870 139.030 42.160 ;
        RECT 131.730 41.660 133.030 41.870 ;
        RECT 128.130 41.160 133.030 41.660 ;
        RECT 133.580 41.470 135.580 41.610 ;
        RECT 133.560 41.300 135.600 41.470 ;
        RECT 124.630 39.960 131.530 40.560 ;
        RECT 124.630 37.860 125.930 39.960 ;
        RECT 126.515 39.610 130.555 39.670 ;
        RECT 126.230 39.440 130.880 39.610 ;
        RECT 126.130 39.060 130.940 39.440 ;
        RECT 126.130 38.440 126.300 39.060 ;
        RECT 130.770 38.440 130.940 39.060 ;
        RECT 126.515 38.210 130.555 38.380 ;
        RECT 126.730 37.860 130.380 38.210 ;
        RECT 131.230 37.860 131.530 39.960 ;
        RECT 124.630 36.960 131.530 37.860 ;
        RECT 124.630 34.860 125.930 36.960 ;
        RECT 126.730 36.670 130.380 36.960 ;
        RECT 126.515 36.500 130.555 36.670 ;
        RECT 126.130 35.440 126.300 36.440 ;
        RECT 130.770 35.440 130.940 36.440 ;
        RECT 126.515 35.210 130.555 35.380 ;
        RECT 131.230 34.860 131.530 36.960 ;
        RECT 124.630 33.660 131.530 34.860 ;
        RECT 132.130 39.660 133.030 41.160 ;
        RECT 133.220 40.240 133.390 41.240 ;
        RECT 134.030 40.180 135.530 40.260 ;
        RECT 135.770 40.240 135.940 41.240 ;
        RECT 133.560 40.010 135.600 40.180 ;
        RECT 134.030 39.660 135.530 40.010 ;
        RECT 136.230 39.960 139.030 41.870 ;
        RECT 139.730 41.810 141.230 42.160 ;
        RECT 139.660 41.640 141.700 41.810 ;
        RECT 139.320 41.360 139.490 41.580 ;
        RECT 141.870 41.360 142.040 41.580 ;
        RECT 139.320 40.580 142.040 41.360 ;
        RECT 139.330 40.360 142.030 40.580 ;
        RECT 139.660 40.350 141.700 40.360 ;
        RECT 142.230 39.960 143.130 42.160 ;
        RECT 136.230 39.660 143.130 39.960 ;
        RECT 132.130 39.260 143.130 39.660 ;
        RECT 132.130 38.960 139.030 39.260 ;
        RECT 132.130 36.760 133.030 38.960 ;
        RECT 133.560 38.560 135.600 38.570 ;
        RECT 133.230 38.340 135.930 38.560 ;
        RECT 133.220 37.560 135.940 38.340 ;
        RECT 133.220 37.340 133.390 37.560 ;
        RECT 135.770 37.340 135.940 37.560 ;
        RECT 133.560 37.110 135.600 37.280 ;
        RECT 134.030 36.760 135.530 37.110 ;
        RECT 136.230 37.050 139.030 38.960 ;
        RECT 139.730 38.910 141.230 39.260 ;
        RECT 139.660 38.740 141.700 38.910 ;
        RECT 139.320 37.680 139.490 38.680 ;
        RECT 139.730 38.660 141.230 38.740 ;
        RECT 141.870 37.680 142.040 38.680 ;
        RECT 142.230 37.760 143.130 39.260 ;
        RECT 143.730 44.060 150.630 45.260 ;
        RECT 143.730 41.960 144.030 44.060 ;
        RECT 144.705 43.540 148.745 43.710 ;
        RECT 144.320 42.480 144.490 43.480 ;
        RECT 148.960 42.480 149.130 43.480 ;
        RECT 144.705 42.250 148.745 42.420 ;
        RECT 144.880 41.960 148.530 42.250 ;
        RECT 149.330 41.960 150.630 44.060 ;
        RECT 143.730 41.060 150.630 41.960 ;
        RECT 143.730 38.960 144.030 41.060 ;
        RECT 144.880 40.710 148.530 41.060 ;
        RECT 144.705 40.540 148.745 40.710 ;
        RECT 144.320 39.860 144.490 40.480 ;
        RECT 148.960 39.860 149.130 40.480 ;
        RECT 144.320 39.480 149.130 39.860 ;
        RECT 144.380 39.310 149.030 39.480 ;
        RECT 144.705 39.250 148.745 39.310 ;
        RECT 149.330 38.960 150.630 41.060 ;
        RECT 143.730 38.360 150.630 38.960 ;
        RECT 139.660 37.450 141.700 37.620 ;
        RECT 139.680 37.310 141.680 37.450 ;
        RECT 142.230 37.260 147.130 37.760 ;
        RECT 142.230 37.050 143.530 37.260 ;
        RECT 136.230 36.760 143.530 37.050 ;
        RECT 132.130 36.360 143.530 36.760 ;
        RECT 144.110 36.740 146.150 36.910 ;
        RECT 132.130 36.060 139.030 36.360 ;
        RECT 132.130 33.960 133.030 36.060 ;
        RECT 133.560 35.660 135.600 35.670 ;
        RECT 133.230 35.440 135.930 35.660 ;
        RECT 133.220 34.660 135.940 35.440 ;
        RECT 133.220 34.440 133.390 34.660 ;
        RECT 135.770 34.440 135.940 34.660 ;
        RECT 133.560 34.210 135.600 34.380 ;
        RECT 136.230 34.260 139.030 36.060 ;
        RECT 139.730 36.010 141.230 36.360 ;
        RECT 139.660 35.840 141.700 36.010 ;
        RECT 139.320 34.780 139.490 35.780 ;
        RECT 139.730 35.760 141.230 35.840 ;
        RECT 141.870 34.780 142.040 35.780 ;
        RECT 142.230 35.060 143.530 36.360 ;
        RECT 143.770 35.680 143.940 36.680 ;
        RECT 146.320 35.680 146.490 36.680 ;
        RECT 144.110 35.450 146.150 35.620 ;
        RECT 146.830 35.060 147.130 37.260 ;
        RECT 139.660 34.550 141.700 34.720 ;
        RECT 142.230 34.460 147.130 35.060 ;
        RECT 147.510 34.530 150.630 38.360 ;
        RECT 142.230 34.260 143.130 34.460 ;
        RECT 134.030 33.960 135.530 34.210 ;
        RECT 136.230 33.960 143.130 34.260 ;
        RECT 124.630 32.390 126.380 33.660 ;
        RECT 132.130 32.960 143.130 33.960 ;
        RECT 148.880 33.260 150.630 34.530 ;
        RECT 132.130 32.660 139.030 32.960 ;
        RECT 139.730 32.710 141.230 32.960 ;
        RECT 132.130 32.460 133.030 32.660 ;
        RECT 124.630 28.560 127.750 32.390 ;
        RECT 128.130 31.860 133.030 32.460 ;
        RECT 133.560 32.200 135.600 32.370 ;
        RECT 128.130 29.660 128.430 31.860 ;
        RECT 129.110 31.300 131.150 31.470 ;
        RECT 128.770 30.240 128.940 31.240 ;
        RECT 131.320 30.240 131.490 31.240 ;
        RECT 131.730 30.560 133.030 31.860 ;
        RECT 133.220 31.140 133.390 32.140 ;
        RECT 134.030 31.080 135.530 31.160 ;
        RECT 135.770 31.140 135.940 32.140 ;
        RECT 133.560 30.910 135.600 31.080 ;
        RECT 134.030 30.560 135.530 30.910 ;
        RECT 136.230 30.860 139.030 32.660 ;
        RECT 139.660 32.540 141.700 32.710 ;
        RECT 139.320 32.260 139.490 32.480 ;
        RECT 141.870 32.260 142.040 32.480 ;
        RECT 139.320 31.480 142.040 32.260 ;
        RECT 139.330 31.260 142.030 31.480 ;
        RECT 139.660 31.250 141.700 31.260 ;
        RECT 142.230 30.860 143.130 32.960 ;
        RECT 136.230 30.560 143.130 30.860 ;
        RECT 129.110 30.010 131.150 30.180 ;
        RECT 131.730 30.160 143.130 30.560 ;
        RECT 131.730 29.870 139.030 30.160 ;
        RECT 131.730 29.660 133.030 29.870 ;
        RECT 128.130 29.160 133.030 29.660 ;
        RECT 133.580 29.470 135.580 29.610 ;
        RECT 133.560 29.300 135.600 29.470 ;
        RECT 124.630 27.960 131.530 28.560 ;
        RECT 124.630 25.860 125.930 27.960 ;
        RECT 126.515 27.610 130.555 27.670 ;
        RECT 126.230 27.440 130.880 27.610 ;
        RECT 126.130 27.060 130.940 27.440 ;
        RECT 126.130 26.440 126.300 27.060 ;
        RECT 130.770 26.440 130.940 27.060 ;
        RECT 126.515 26.210 130.555 26.380 ;
        RECT 126.730 25.860 130.380 26.210 ;
        RECT 131.230 25.860 131.530 27.960 ;
        RECT 124.630 24.960 131.530 25.860 ;
        RECT 124.630 22.860 125.930 24.960 ;
        RECT 126.730 24.670 130.380 24.960 ;
        RECT 126.515 24.500 130.555 24.670 ;
        RECT 126.130 23.440 126.300 24.440 ;
        RECT 130.770 23.440 130.940 24.440 ;
        RECT 126.515 23.210 130.555 23.380 ;
        RECT 131.230 22.860 131.530 24.960 ;
        RECT 124.630 21.960 131.530 22.860 ;
        RECT 132.130 27.660 133.030 29.160 ;
        RECT 133.220 28.240 133.390 29.240 ;
        RECT 134.030 28.180 135.530 28.260 ;
        RECT 135.770 28.240 135.940 29.240 ;
        RECT 133.560 28.010 135.600 28.180 ;
        RECT 134.030 27.660 135.530 28.010 ;
        RECT 136.230 27.960 139.030 29.870 ;
        RECT 139.730 29.810 141.230 30.160 ;
        RECT 139.660 29.640 141.700 29.810 ;
        RECT 139.320 29.360 139.490 29.580 ;
        RECT 141.870 29.360 142.040 29.580 ;
        RECT 139.320 28.580 142.040 29.360 ;
        RECT 139.330 28.360 142.030 28.580 ;
        RECT 139.660 28.350 141.700 28.360 ;
        RECT 142.230 27.960 143.130 30.160 ;
        RECT 136.230 27.660 143.130 27.960 ;
        RECT 132.130 27.260 143.130 27.660 ;
        RECT 132.130 26.960 139.030 27.260 ;
        RECT 132.130 24.760 133.030 26.960 ;
        RECT 133.560 26.560 135.600 26.570 ;
        RECT 133.230 26.340 135.930 26.560 ;
        RECT 133.220 25.560 135.940 26.340 ;
        RECT 133.220 25.340 133.390 25.560 ;
        RECT 135.770 25.340 135.940 25.560 ;
        RECT 133.560 25.110 135.600 25.280 ;
        RECT 134.030 24.760 135.530 25.110 ;
        RECT 136.230 25.050 139.030 26.960 ;
        RECT 139.730 26.910 141.230 27.260 ;
        RECT 139.660 26.740 141.700 26.910 ;
        RECT 139.320 25.680 139.490 26.680 ;
        RECT 139.730 26.660 141.230 26.740 ;
        RECT 141.870 25.680 142.040 26.680 ;
        RECT 142.230 25.760 143.130 27.260 ;
        RECT 143.730 32.060 150.630 33.260 ;
        RECT 143.730 29.960 144.030 32.060 ;
        RECT 144.705 31.540 148.745 31.710 ;
        RECT 144.320 30.480 144.490 31.480 ;
        RECT 148.960 30.480 149.130 31.480 ;
        RECT 144.705 30.250 148.745 30.420 ;
        RECT 144.880 29.960 148.530 30.250 ;
        RECT 149.330 29.960 150.630 32.060 ;
        RECT 143.730 29.060 150.630 29.960 ;
        RECT 143.730 26.960 144.030 29.060 ;
        RECT 144.880 28.710 148.530 29.060 ;
        RECT 144.705 28.540 148.745 28.710 ;
        RECT 144.320 27.860 144.490 28.480 ;
        RECT 148.960 27.860 149.130 28.480 ;
        RECT 144.320 27.480 149.130 27.860 ;
        RECT 144.380 27.310 149.030 27.480 ;
        RECT 144.705 27.250 148.745 27.310 ;
        RECT 149.330 26.960 150.630 29.060 ;
        RECT 143.730 26.360 150.630 26.960 ;
        RECT 139.660 25.450 141.700 25.620 ;
        RECT 139.680 25.310 141.680 25.450 ;
        RECT 142.230 25.260 147.130 25.760 ;
        RECT 142.230 25.050 143.530 25.260 ;
        RECT 136.230 24.760 143.530 25.050 ;
        RECT 132.130 24.360 143.530 24.760 ;
        RECT 144.110 24.740 146.150 24.910 ;
        RECT 132.130 24.060 139.030 24.360 ;
        RECT 132.130 21.960 133.030 24.060 ;
        RECT 133.560 23.660 135.600 23.670 ;
        RECT 133.230 23.440 135.930 23.660 ;
        RECT 133.220 22.660 135.940 23.440 ;
        RECT 133.220 22.440 133.390 22.660 ;
        RECT 135.770 22.440 135.940 22.660 ;
        RECT 133.560 22.210 135.600 22.380 ;
        RECT 136.230 22.260 139.030 24.060 ;
        RECT 139.730 24.010 141.230 24.360 ;
        RECT 139.660 23.840 141.700 24.010 ;
        RECT 139.320 22.780 139.490 23.780 ;
        RECT 139.730 23.760 141.230 23.840 ;
        RECT 141.870 22.780 142.040 23.780 ;
        RECT 142.230 23.060 143.530 24.360 ;
        RECT 143.770 23.680 143.940 24.680 ;
        RECT 146.320 23.680 146.490 24.680 ;
        RECT 144.110 23.450 146.150 23.620 ;
        RECT 146.830 23.060 147.130 25.260 ;
        RECT 139.660 22.550 141.700 22.720 ;
        RECT 142.230 22.460 147.130 23.060 ;
        RECT 147.510 22.530 150.630 26.360 ;
        RECT 142.230 22.260 143.130 22.460 ;
        RECT 134.030 21.960 135.530 22.210 ;
        RECT 136.230 21.960 143.130 22.260 ;
        RECT 124.630 20.460 131.630 21.960 ;
        RECT 132.130 20.960 143.130 21.960 ;
        RECT 148.880 21.460 150.630 22.530 ;
        RECT 148.885 20.960 150.630 21.460 ;
        RECT 151.130 20.960 154.130 72.160 ;
        RECT 124.630 20.360 131.530 20.460 ;
        RECT 124.530 20.060 131.530 20.360 ;
        RECT 121.730 19.760 131.530 20.060 ;
        RECT 132.130 19.960 146.930 20.960 ;
        RECT 116.780 19.560 131.530 19.760 ;
        RECT 116.780 19.360 143.330 19.560 ;
        RECT 116.780 19.120 143.430 19.360 ;
        RECT 116.780 16.960 132.030 19.120 ;
        RECT 135.130 19.060 143.430 19.120 ;
        RECT 132.730 18.720 136.630 18.760 ;
        RECT 132.715 18.550 136.755 18.720 ;
        RECT 132.330 17.490 132.500 18.490 ;
        RECT 132.730 18.060 136.630 18.550 ;
        RECT 136.970 17.490 137.140 18.490 ;
        RECT 133.230 17.430 136.330 17.460 ;
        RECT 132.715 17.260 136.755 17.430 ;
        RECT 133.230 16.960 136.330 17.260 ;
        RECT 137.370 16.960 137.650 19.060 ;
        RECT 138.265 18.550 142.305 18.720 ;
        RECT 137.880 17.490 138.050 18.490 ;
        RECT 142.520 17.490 142.690 18.490 ;
        RECT 138.430 17.430 142.130 17.460 ;
        RECT 138.265 17.260 142.305 17.430 ;
        RECT 138.430 16.960 142.130 17.260 ;
        RECT 142.930 16.960 143.430 19.060 ;
        RECT 144.030 17.760 146.930 19.960 ;
        RECT 148.885 19.460 154.130 20.960 ;
        RECT 149.130 16.960 154.130 19.460 ;
        RECT 116.780 15.160 154.130 16.960 ;
        RECT 116.780 14.460 138.030 15.160 ;
        RECT 141.930 14.460 154.130 15.160 ;
        RECT 116.780 12.380 124.050 14.460 ;
      LAYER met1 ;
        RECT 121.730 20.060 123.830 74.060 ;
        RECT 124.630 70.460 150.630 72.460 ;
        RECT 124.630 69.460 126.130 70.460 ;
        RECT 149.130 69.460 150.630 70.460 ;
        RECT 124.630 68.390 126.380 69.460 ;
        RECT 132.130 68.960 143.030 69.460 ;
        RECT 148.880 69.260 150.630 69.460 ;
        RECT 132.130 68.710 139.030 68.960 ;
        RECT 139.730 68.740 141.230 68.960 ;
        RECT 132.130 68.660 133.080 68.710 ;
        RECT 132.130 68.460 133.030 68.660 ;
        RECT 124.630 64.560 127.750 68.390 ;
        RECT 128.130 67.860 133.030 68.460 ;
        RECT 133.630 68.400 135.580 68.510 ;
        RECT 133.580 68.170 135.580 68.400 ;
        RECT 128.130 65.660 128.430 67.860 ;
        RECT 129.330 67.500 131.130 67.660 ;
        RECT 129.130 67.270 131.130 67.500 ;
        RECT 128.740 67.110 128.970 67.220 ;
        RECT 129.330 67.210 131.130 67.270 ;
        RECT 129.330 67.110 130.880 67.210 ;
        RECT 128.730 67.060 129.030 67.110 ;
        RECT 131.290 67.060 131.520 67.220 ;
        RECT 128.730 66.960 129.130 67.060 ;
        RECT 131.130 66.960 131.530 67.060 ;
        RECT 128.730 66.510 131.530 66.960 ;
        RECT 128.730 66.360 129.130 66.510 ;
        RECT 131.180 66.360 131.530 66.510 ;
        RECT 131.730 66.560 133.030 67.860 ;
        RECT 133.190 67.960 133.420 68.120 ;
        RECT 135.740 67.960 135.970 68.120 ;
        RECT 133.190 67.360 135.970 67.960 ;
        RECT 133.190 67.160 133.420 67.360 ;
        RECT 135.740 67.160 135.970 67.360 ;
        RECT 134.030 67.110 135.530 67.160 ;
        RECT 133.580 66.880 135.580 67.110 ;
        RECT 134.030 66.560 135.530 66.880 ;
        RECT 136.230 66.860 139.030 68.710 ;
        RECT 139.680 68.510 141.680 68.740 ;
        RECT 139.290 68.260 139.520 68.460 ;
        RECT 141.840 68.450 142.070 68.460 ;
        RECT 141.840 68.310 142.130 68.450 ;
        RECT 141.730 68.260 142.130 68.310 ;
        RECT 139.290 67.500 142.130 68.260 ;
        RECT 139.330 67.310 142.130 67.500 ;
        RECT 139.330 67.260 142.030 67.310 ;
        RECT 139.680 67.220 141.680 67.260 ;
        RECT 142.330 66.860 143.030 68.960 ;
        RECT 136.230 66.560 143.030 66.860 ;
        RECT 128.730 66.310 129.030 66.360 ;
        RECT 128.740 66.260 128.970 66.310 ;
        RECT 131.290 66.260 131.520 66.360 ;
        RECT 129.430 66.210 131.030 66.260 ;
        RECT 129.130 65.980 131.130 66.210 ;
        RECT 131.730 66.160 143.030 66.560 ;
        RECT 129.430 65.810 131.080 65.980 ;
        RECT 131.730 65.960 139.030 66.160 ;
        RECT 131.730 65.660 133.030 65.960 ;
        RECT 136.180 65.910 139.030 65.960 ;
        RECT 133.630 65.760 134.130 65.810 ;
        RECT 128.130 65.160 133.030 65.660 ;
        RECT 133.580 65.270 135.580 65.760 ;
        RECT 124.630 63.990 131.530 64.560 ;
        RECT 124.630 62.260 125.930 63.990 ;
        RECT 131.210 63.960 131.530 63.990 ;
        RECT 126.535 63.660 130.535 63.700 ;
        RECT 126.130 63.420 130.930 63.660 ;
        RECT 126.100 62.560 130.970 63.420 ;
        RECT 126.100 62.460 126.330 62.560 ;
        RECT 130.740 62.460 130.970 62.560 ;
        RECT 126.535 62.260 130.535 62.410 ;
        RECT 131.230 62.260 131.530 63.960 ;
        RECT 124.630 60.660 131.530 62.260 ;
        RECT 124.630 60.560 130.535 60.660 ;
        RECT 124.630 58.860 125.930 60.560 ;
        RECT 126.535 60.470 130.535 60.560 ;
        RECT 126.100 60.260 126.330 60.420 ;
        RECT 130.740 60.260 130.970 60.420 ;
        RECT 126.100 59.760 130.970 60.260 ;
        RECT 126.100 59.660 126.430 59.760 ;
        RECT 126.100 59.460 126.330 59.660 ;
        RECT 127.230 59.610 127.530 59.760 ;
        RECT 130.730 59.660 130.970 59.760 ;
        RECT 128.530 59.410 130.330 59.510 ;
        RECT 130.740 59.460 130.970 59.660 ;
        RECT 126.535 59.180 130.535 59.410 ;
        RECT 128.530 59.010 130.330 59.180 ;
        RECT 131.230 58.860 131.530 60.660 ;
        RECT 124.630 57.660 131.530 58.860 ;
        RECT 132.230 63.660 133.030 65.160 ;
        RECT 133.190 65.060 133.420 65.220 ;
        RECT 135.740 65.060 135.970 65.220 ;
        RECT 133.190 64.460 135.970 65.060 ;
        RECT 133.190 64.260 133.420 64.460 ;
        RECT 135.740 64.260 135.970 64.460 ;
        RECT 134.030 64.210 135.530 64.260 ;
        RECT 133.580 63.980 135.580 64.210 ;
        RECT 134.030 63.660 135.530 63.980 ;
        RECT 136.230 63.960 139.030 65.910 ;
        RECT 139.730 65.840 141.230 66.160 ;
        RECT 139.680 65.610 141.680 65.840 ;
        RECT 139.290 65.360 139.520 65.560 ;
        RECT 141.840 65.360 142.070 65.560 ;
        RECT 139.290 64.600 142.070 65.360 ;
        RECT 139.330 64.360 142.030 64.600 ;
        RECT 139.680 64.320 141.680 64.360 ;
        RECT 142.230 63.960 143.030 66.160 ;
        RECT 136.230 63.660 143.030 63.960 ;
        RECT 132.230 63.260 143.030 63.660 ;
        RECT 132.230 62.960 139.030 63.260 ;
        RECT 132.230 60.760 133.030 62.960 ;
        RECT 133.580 62.560 135.580 62.600 ;
        RECT 133.230 62.320 135.930 62.560 ;
        RECT 133.190 61.560 135.970 62.320 ;
        RECT 133.190 61.360 133.420 61.560 ;
        RECT 135.740 61.360 135.970 61.560 ;
        RECT 133.580 61.080 135.580 61.310 ;
        RECT 134.030 60.760 135.530 61.080 ;
        RECT 136.230 61.010 139.030 62.960 ;
        RECT 139.730 62.940 141.230 63.260 ;
        RECT 139.680 62.710 141.680 62.940 ;
        RECT 139.730 62.660 141.230 62.710 ;
        RECT 139.290 62.460 139.520 62.660 ;
        RECT 141.840 62.460 142.070 62.660 ;
        RECT 139.290 61.860 142.070 62.460 ;
        RECT 139.290 61.700 139.520 61.860 ;
        RECT 141.840 61.700 142.070 61.860 ;
        RECT 142.230 61.760 143.030 63.260 ;
        RECT 143.730 68.060 150.630 69.260 ;
        RECT 143.730 66.260 144.030 68.060 ;
        RECT 144.930 67.740 146.730 67.910 ;
        RECT 144.725 67.510 148.725 67.740 ;
        RECT 144.290 67.260 144.520 67.460 ;
        RECT 144.930 67.410 146.730 67.510 ;
        RECT 144.290 67.160 144.530 67.260 ;
        RECT 147.730 67.160 148.030 67.310 ;
        RECT 148.930 67.260 149.160 67.460 ;
        RECT 148.830 67.160 149.160 67.260 ;
        RECT 144.290 66.660 149.160 67.160 ;
        RECT 144.290 66.500 144.520 66.660 ;
        RECT 148.930 66.500 149.160 66.660 ;
        RECT 144.725 66.360 148.725 66.450 ;
        RECT 149.330 66.360 150.630 68.060 ;
        RECT 144.725 66.260 150.630 66.360 ;
        RECT 143.730 64.660 150.630 66.260 ;
        RECT 143.730 62.960 144.030 64.660 ;
        RECT 144.725 64.510 148.725 64.660 ;
        RECT 144.290 64.360 144.520 64.460 ;
        RECT 148.930 64.360 149.160 64.460 ;
        RECT 144.290 63.500 149.160 64.360 ;
        RECT 144.330 63.260 149.130 63.500 ;
        RECT 144.725 63.220 148.725 63.260 ;
        RECT 143.730 62.930 144.050 62.960 ;
        RECT 149.330 62.930 150.630 64.660 ;
        RECT 143.730 62.360 150.630 62.930 ;
        RECT 139.680 61.160 141.680 61.650 ;
        RECT 142.230 61.260 147.130 61.760 ;
        RECT 141.130 61.110 141.630 61.160 ;
        RECT 136.230 60.960 139.080 61.010 ;
        RECT 142.230 60.960 143.530 61.260 ;
        RECT 136.230 60.760 143.530 60.960 ;
        RECT 144.180 60.940 145.830 61.110 ;
        RECT 132.230 60.360 143.530 60.760 ;
        RECT 144.130 60.710 146.130 60.940 ;
        RECT 144.230 60.660 145.830 60.710 ;
        RECT 143.740 60.560 143.970 60.660 ;
        RECT 146.290 60.610 146.520 60.660 ;
        RECT 146.230 60.560 146.530 60.610 ;
        RECT 132.230 60.060 139.030 60.360 ;
        RECT 132.230 57.960 132.930 60.060 ;
        RECT 133.580 59.660 135.580 59.700 ;
        RECT 133.230 59.610 135.930 59.660 ;
        RECT 133.130 59.420 135.930 59.610 ;
        RECT 133.130 58.660 135.970 59.420 ;
        RECT 133.130 58.610 133.530 58.660 ;
        RECT 133.130 58.470 133.420 58.610 ;
        RECT 133.190 58.460 133.420 58.470 ;
        RECT 135.740 58.460 135.970 58.660 ;
        RECT 133.580 58.180 135.580 58.410 ;
        RECT 136.230 58.210 139.030 60.060 ;
        RECT 139.730 60.040 141.230 60.360 ;
        RECT 139.680 59.810 141.680 60.040 ;
        RECT 139.730 59.760 141.230 59.810 ;
        RECT 139.290 59.560 139.520 59.760 ;
        RECT 141.840 59.560 142.070 59.760 ;
        RECT 139.290 58.960 142.070 59.560 ;
        RECT 139.290 58.800 139.520 58.960 ;
        RECT 141.840 58.800 142.070 58.960 ;
        RECT 142.230 59.060 143.530 60.360 ;
        RECT 143.730 60.410 144.080 60.560 ;
        RECT 146.130 60.410 146.530 60.560 ;
        RECT 143.730 59.960 146.530 60.410 ;
        RECT 143.730 59.860 144.130 59.960 ;
        RECT 146.130 59.860 146.530 59.960 ;
        RECT 143.740 59.700 143.970 59.860 ;
        RECT 146.230 59.810 146.530 59.860 ;
        RECT 144.380 59.710 145.930 59.810 ;
        RECT 144.130 59.650 145.930 59.710 ;
        RECT 146.290 59.700 146.520 59.810 ;
        RECT 144.130 59.420 146.130 59.650 ;
        RECT 144.130 59.260 145.930 59.420 ;
        RECT 146.830 59.060 147.130 61.260 ;
        RECT 139.680 58.520 141.680 58.750 ;
        RECT 139.680 58.410 141.630 58.520 ;
        RECT 142.230 58.460 147.130 59.060 ;
        RECT 147.510 58.530 150.630 62.360 ;
        RECT 142.230 58.260 143.130 58.460 ;
        RECT 142.180 58.210 143.130 58.260 ;
        RECT 134.030 57.960 135.530 58.180 ;
        RECT 136.230 57.960 143.130 58.210 ;
        RECT 124.630 56.390 126.380 57.660 ;
        RECT 132.230 57.460 143.130 57.960 ;
        RECT 132.130 56.960 143.030 57.460 ;
        RECT 148.880 57.260 150.630 58.530 ;
        RECT 132.130 56.710 139.030 56.960 ;
        RECT 139.730 56.740 141.230 56.960 ;
        RECT 132.130 56.660 133.080 56.710 ;
        RECT 132.130 56.460 133.030 56.660 ;
        RECT 124.630 52.560 127.750 56.390 ;
        RECT 128.130 55.860 133.030 56.460 ;
        RECT 133.630 56.400 135.580 56.510 ;
        RECT 133.580 56.170 135.580 56.400 ;
        RECT 128.130 53.660 128.430 55.860 ;
        RECT 129.330 55.500 131.130 55.660 ;
        RECT 129.130 55.270 131.130 55.500 ;
        RECT 128.740 55.110 128.970 55.220 ;
        RECT 129.330 55.210 131.130 55.270 ;
        RECT 129.330 55.110 130.880 55.210 ;
        RECT 128.730 55.060 129.030 55.110 ;
        RECT 131.290 55.060 131.520 55.220 ;
        RECT 128.730 54.960 129.130 55.060 ;
        RECT 131.130 54.960 131.530 55.060 ;
        RECT 128.730 54.510 131.530 54.960 ;
        RECT 128.730 54.360 129.130 54.510 ;
        RECT 131.180 54.360 131.530 54.510 ;
        RECT 131.730 54.560 133.030 55.860 ;
        RECT 133.190 55.960 133.420 56.120 ;
        RECT 135.740 55.960 135.970 56.120 ;
        RECT 133.190 55.360 135.970 55.960 ;
        RECT 133.190 55.160 133.420 55.360 ;
        RECT 135.740 55.160 135.970 55.360 ;
        RECT 134.030 55.110 135.530 55.160 ;
        RECT 133.580 54.880 135.580 55.110 ;
        RECT 134.030 54.560 135.530 54.880 ;
        RECT 136.230 54.860 139.030 56.710 ;
        RECT 139.680 56.510 141.680 56.740 ;
        RECT 139.290 56.260 139.520 56.460 ;
        RECT 141.840 56.450 142.070 56.460 ;
        RECT 141.840 56.310 142.130 56.450 ;
        RECT 141.730 56.260 142.130 56.310 ;
        RECT 139.290 55.500 142.130 56.260 ;
        RECT 139.330 55.310 142.130 55.500 ;
        RECT 139.330 55.260 142.030 55.310 ;
        RECT 139.680 55.220 141.680 55.260 ;
        RECT 142.330 54.860 143.030 56.960 ;
        RECT 136.230 54.560 143.030 54.860 ;
        RECT 128.730 54.310 129.030 54.360 ;
        RECT 128.740 54.260 128.970 54.310 ;
        RECT 131.290 54.260 131.520 54.360 ;
        RECT 129.430 54.210 131.030 54.260 ;
        RECT 129.130 53.980 131.130 54.210 ;
        RECT 131.730 54.160 143.030 54.560 ;
        RECT 129.430 53.810 131.080 53.980 ;
        RECT 131.730 53.960 139.030 54.160 ;
        RECT 131.730 53.660 133.030 53.960 ;
        RECT 136.180 53.910 139.030 53.960 ;
        RECT 133.630 53.760 134.130 53.810 ;
        RECT 128.130 53.160 133.030 53.660 ;
        RECT 133.580 53.270 135.580 53.760 ;
        RECT 124.630 51.990 131.530 52.560 ;
        RECT 124.630 50.260 125.930 51.990 ;
        RECT 131.210 51.960 131.530 51.990 ;
        RECT 126.535 51.660 130.535 51.700 ;
        RECT 126.130 51.420 130.930 51.660 ;
        RECT 126.100 50.560 130.970 51.420 ;
        RECT 126.100 50.460 126.330 50.560 ;
        RECT 130.740 50.460 130.970 50.560 ;
        RECT 126.535 50.260 130.535 50.410 ;
        RECT 131.230 50.260 131.530 51.960 ;
        RECT 124.630 48.660 131.530 50.260 ;
        RECT 124.630 48.560 130.535 48.660 ;
        RECT 124.630 46.860 125.930 48.560 ;
        RECT 126.535 48.470 130.535 48.560 ;
        RECT 126.100 48.260 126.330 48.420 ;
        RECT 130.740 48.260 130.970 48.420 ;
        RECT 126.100 47.760 130.970 48.260 ;
        RECT 126.100 47.660 126.430 47.760 ;
        RECT 126.100 47.460 126.330 47.660 ;
        RECT 127.230 47.610 127.530 47.760 ;
        RECT 130.730 47.660 130.970 47.760 ;
        RECT 128.530 47.410 130.330 47.510 ;
        RECT 130.740 47.460 130.970 47.660 ;
        RECT 126.535 47.180 130.535 47.410 ;
        RECT 128.530 47.010 130.330 47.180 ;
        RECT 131.230 46.860 131.530 48.660 ;
        RECT 124.630 45.660 131.530 46.860 ;
        RECT 132.230 51.660 133.030 53.160 ;
        RECT 133.190 53.060 133.420 53.220 ;
        RECT 135.740 53.060 135.970 53.220 ;
        RECT 133.190 52.460 135.970 53.060 ;
        RECT 133.190 52.260 133.420 52.460 ;
        RECT 135.740 52.260 135.970 52.460 ;
        RECT 134.030 52.210 135.530 52.260 ;
        RECT 133.580 51.980 135.580 52.210 ;
        RECT 134.030 51.660 135.530 51.980 ;
        RECT 136.230 51.960 139.030 53.910 ;
        RECT 139.730 53.840 141.230 54.160 ;
        RECT 139.680 53.610 141.680 53.840 ;
        RECT 139.290 53.360 139.520 53.560 ;
        RECT 141.840 53.360 142.070 53.560 ;
        RECT 139.290 52.600 142.070 53.360 ;
        RECT 139.330 52.360 142.030 52.600 ;
        RECT 139.680 52.320 141.680 52.360 ;
        RECT 142.230 51.960 143.030 54.160 ;
        RECT 136.230 51.660 143.030 51.960 ;
        RECT 132.230 51.260 143.030 51.660 ;
        RECT 132.230 50.960 139.030 51.260 ;
        RECT 132.230 48.760 133.030 50.960 ;
        RECT 133.580 50.560 135.580 50.600 ;
        RECT 133.230 50.320 135.930 50.560 ;
        RECT 133.190 49.560 135.970 50.320 ;
        RECT 133.190 49.360 133.420 49.560 ;
        RECT 135.740 49.360 135.970 49.560 ;
        RECT 133.580 49.080 135.580 49.310 ;
        RECT 134.030 48.760 135.530 49.080 ;
        RECT 136.230 49.010 139.030 50.960 ;
        RECT 139.730 50.940 141.230 51.260 ;
        RECT 139.680 50.710 141.680 50.940 ;
        RECT 139.730 50.660 141.230 50.710 ;
        RECT 139.290 50.460 139.520 50.660 ;
        RECT 141.840 50.460 142.070 50.660 ;
        RECT 139.290 49.860 142.070 50.460 ;
        RECT 139.290 49.700 139.520 49.860 ;
        RECT 141.840 49.700 142.070 49.860 ;
        RECT 142.230 49.760 143.030 51.260 ;
        RECT 143.730 56.060 150.630 57.260 ;
        RECT 143.730 54.260 144.030 56.060 ;
        RECT 144.930 55.740 146.730 55.910 ;
        RECT 144.725 55.510 148.725 55.740 ;
        RECT 144.290 55.260 144.520 55.460 ;
        RECT 144.930 55.410 146.730 55.510 ;
        RECT 144.290 55.160 144.530 55.260 ;
        RECT 147.730 55.160 148.030 55.310 ;
        RECT 148.930 55.260 149.160 55.460 ;
        RECT 148.830 55.160 149.160 55.260 ;
        RECT 144.290 54.660 149.160 55.160 ;
        RECT 144.290 54.500 144.520 54.660 ;
        RECT 148.930 54.500 149.160 54.660 ;
        RECT 144.725 54.360 148.725 54.450 ;
        RECT 149.330 54.360 150.630 56.060 ;
        RECT 144.725 54.260 150.630 54.360 ;
        RECT 143.730 52.660 150.630 54.260 ;
        RECT 143.730 50.960 144.030 52.660 ;
        RECT 144.725 52.510 148.725 52.660 ;
        RECT 144.290 52.360 144.520 52.460 ;
        RECT 148.930 52.360 149.160 52.460 ;
        RECT 144.290 51.500 149.160 52.360 ;
        RECT 144.330 51.260 149.130 51.500 ;
        RECT 144.725 51.220 148.725 51.260 ;
        RECT 143.730 50.930 144.050 50.960 ;
        RECT 149.330 50.930 150.630 52.660 ;
        RECT 143.730 50.360 150.630 50.930 ;
        RECT 139.680 49.160 141.680 49.650 ;
        RECT 142.230 49.260 147.130 49.760 ;
        RECT 141.130 49.110 141.630 49.160 ;
        RECT 136.230 48.960 139.080 49.010 ;
        RECT 142.230 48.960 143.530 49.260 ;
        RECT 136.230 48.760 143.530 48.960 ;
        RECT 144.180 48.940 145.830 49.110 ;
        RECT 132.230 48.360 143.530 48.760 ;
        RECT 144.130 48.710 146.130 48.940 ;
        RECT 144.230 48.660 145.830 48.710 ;
        RECT 143.740 48.560 143.970 48.660 ;
        RECT 146.290 48.610 146.520 48.660 ;
        RECT 146.230 48.560 146.530 48.610 ;
        RECT 132.230 48.060 139.030 48.360 ;
        RECT 132.230 45.960 132.930 48.060 ;
        RECT 133.580 47.660 135.580 47.700 ;
        RECT 133.230 47.610 135.930 47.660 ;
        RECT 133.130 47.420 135.930 47.610 ;
        RECT 133.130 46.660 135.970 47.420 ;
        RECT 133.130 46.610 133.530 46.660 ;
        RECT 133.130 46.470 133.420 46.610 ;
        RECT 133.190 46.460 133.420 46.470 ;
        RECT 135.740 46.460 135.970 46.660 ;
        RECT 133.580 46.180 135.580 46.410 ;
        RECT 136.230 46.210 139.030 48.060 ;
        RECT 139.730 48.040 141.230 48.360 ;
        RECT 139.680 47.810 141.680 48.040 ;
        RECT 139.730 47.760 141.230 47.810 ;
        RECT 139.290 47.560 139.520 47.760 ;
        RECT 141.840 47.560 142.070 47.760 ;
        RECT 139.290 46.960 142.070 47.560 ;
        RECT 139.290 46.800 139.520 46.960 ;
        RECT 141.840 46.800 142.070 46.960 ;
        RECT 142.230 47.060 143.530 48.360 ;
        RECT 143.730 48.410 144.080 48.560 ;
        RECT 146.130 48.410 146.530 48.560 ;
        RECT 143.730 47.960 146.530 48.410 ;
        RECT 143.730 47.860 144.130 47.960 ;
        RECT 146.130 47.860 146.530 47.960 ;
        RECT 143.740 47.700 143.970 47.860 ;
        RECT 146.230 47.810 146.530 47.860 ;
        RECT 144.380 47.710 145.930 47.810 ;
        RECT 144.130 47.650 145.930 47.710 ;
        RECT 146.290 47.700 146.520 47.810 ;
        RECT 144.130 47.420 146.130 47.650 ;
        RECT 144.130 47.260 145.930 47.420 ;
        RECT 146.830 47.060 147.130 49.260 ;
        RECT 139.680 46.520 141.680 46.750 ;
        RECT 139.680 46.410 141.630 46.520 ;
        RECT 142.230 46.460 147.130 47.060 ;
        RECT 147.510 46.530 150.630 50.360 ;
        RECT 142.230 46.260 143.130 46.460 ;
        RECT 142.180 46.210 143.130 46.260 ;
        RECT 134.030 45.960 135.530 46.180 ;
        RECT 136.230 45.960 143.130 46.210 ;
        RECT 124.630 44.390 126.380 45.660 ;
        RECT 132.230 45.460 143.130 45.960 ;
        RECT 132.130 44.960 143.030 45.460 ;
        RECT 148.880 45.260 150.630 46.530 ;
        RECT 132.130 44.710 139.030 44.960 ;
        RECT 139.730 44.740 141.230 44.960 ;
        RECT 132.130 44.660 133.080 44.710 ;
        RECT 132.130 44.460 133.030 44.660 ;
        RECT 124.630 40.560 127.750 44.390 ;
        RECT 128.130 43.860 133.030 44.460 ;
        RECT 133.630 44.400 135.580 44.510 ;
        RECT 133.580 44.170 135.580 44.400 ;
        RECT 128.130 41.660 128.430 43.860 ;
        RECT 129.330 43.500 131.130 43.660 ;
        RECT 129.130 43.270 131.130 43.500 ;
        RECT 128.740 43.110 128.970 43.220 ;
        RECT 129.330 43.210 131.130 43.270 ;
        RECT 129.330 43.110 130.880 43.210 ;
        RECT 128.730 43.060 129.030 43.110 ;
        RECT 131.290 43.060 131.520 43.220 ;
        RECT 128.730 42.960 129.130 43.060 ;
        RECT 131.130 42.960 131.530 43.060 ;
        RECT 128.730 42.510 131.530 42.960 ;
        RECT 128.730 42.360 129.130 42.510 ;
        RECT 131.180 42.360 131.530 42.510 ;
        RECT 131.730 42.560 133.030 43.860 ;
        RECT 133.190 43.960 133.420 44.120 ;
        RECT 135.740 43.960 135.970 44.120 ;
        RECT 133.190 43.360 135.970 43.960 ;
        RECT 133.190 43.160 133.420 43.360 ;
        RECT 135.740 43.160 135.970 43.360 ;
        RECT 134.030 43.110 135.530 43.160 ;
        RECT 133.580 42.880 135.580 43.110 ;
        RECT 134.030 42.560 135.530 42.880 ;
        RECT 136.230 42.860 139.030 44.710 ;
        RECT 139.680 44.510 141.680 44.740 ;
        RECT 139.290 44.260 139.520 44.460 ;
        RECT 141.840 44.450 142.070 44.460 ;
        RECT 141.840 44.310 142.130 44.450 ;
        RECT 141.730 44.260 142.130 44.310 ;
        RECT 139.290 43.500 142.130 44.260 ;
        RECT 139.330 43.310 142.130 43.500 ;
        RECT 139.330 43.260 142.030 43.310 ;
        RECT 139.680 43.220 141.680 43.260 ;
        RECT 142.330 42.860 143.030 44.960 ;
        RECT 136.230 42.560 143.030 42.860 ;
        RECT 128.730 42.310 129.030 42.360 ;
        RECT 128.740 42.260 128.970 42.310 ;
        RECT 131.290 42.260 131.520 42.360 ;
        RECT 129.430 42.210 131.030 42.260 ;
        RECT 129.130 41.980 131.130 42.210 ;
        RECT 131.730 42.160 143.030 42.560 ;
        RECT 129.430 41.810 131.080 41.980 ;
        RECT 131.730 41.960 139.030 42.160 ;
        RECT 131.730 41.660 133.030 41.960 ;
        RECT 136.180 41.910 139.030 41.960 ;
        RECT 133.630 41.760 134.130 41.810 ;
        RECT 128.130 41.160 133.030 41.660 ;
        RECT 133.580 41.270 135.580 41.760 ;
        RECT 124.630 39.990 131.530 40.560 ;
        RECT 124.630 38.260 125.930 39.990 ;
        RECT 131.210 39.960 131.530 39.990 ;
        RECT 126.535 39.660 130.535 39.700 ;
        RECT 126.130 39.420 130.930 39.660 ;
        RECT 126.100 38.560 130.970 39.420 ;
        RECT 126.100 38.460 126.330 38.560 ;
        RECT 130.740 38.460 130.970 38.560 ;
        RECT 126.535 38.260 130.535 38.410 ;
        RECT 131.230 38.260 131.530 39.960 ;
        RECT 124.630 36.660 131.530 38.260 ;
        RECT 124.630 36.560 130.535 36.660 ;
        RECT 124.630 34.860 125.930 36.560 ;
        RECT 126.535 36.470 130.535 36.560 ;
        RECT 126.100 36.260 126.330 36.420 ;
        RECT 130.740 36.260 130.970 36.420 ;
        RECT 126.100 35.760 130.970 36.260 ;
        RECT 126.100 35.660 126.430 35.760 ;
        RECT 126.100 35.460 126.330 35.660 ;
        RECT 127.230 35.610 127.530 35.760 ;
        RECT 130.730 35.660 130.970 35.760 ;
        RECT 128.530 35.410 130.330 35.510 ;
        RECT 130.740 35.460 130.970 35.660 ;
        RECT 126.535 35.180 130.535 35.410 ;
        RECT 128.530 35.010 130.330 35.180 ;
        RECT 131.230 34.860 131.530 36.660 ;
        RECT 124.630 33.660 131.530 34.860 ;
        RECT 132.230 39.660 133.030 41.160 ;
        RECT 133.190 41.060 133.420 41.220 ;
        RECT 135.740 41.060 135.970 41.220 ;
        RECT 133.190 40.460 135.970 41.060 ;
        RECT 133.190 40.260 133.420 40.460 ;
        RECT 135.740 40.260 135.970 40.460 ;
        RECT 134.030 40.210 135.530 40.260 ;
        RECT 133.580 39.980 135.580 40.210 ;
        RECT 134.030 39.660 135.530 39.980 ;
        RECT 136.230 39.960 139.030 41.910 ;
        RECT 139.730 41.840 141.230 42.160 ;
        RECT 139.680 41.610 141.680 41.840 ;
        RECT 139.290 41.360 139.520 41.560 ;
        RECT 141.840 41.360 142.070 41.560 ;
        RECT 139.290 40.600 142.070 41.360 ;
        RECT 139.330 40.360 142.030 40.600 ;
        RECT 139.680 40.320 141.680 40.360 ;
        RECT 142.230 39.960 143.030 42.160 ;
        RECT 136.230 39.660 143.030 39.960 ;
        RECT 132.230 39.260 143.030 39.660 ;
        RECT 132.230 38.960 139.030 39.260 ;
        RECT 132.230 36.760 133.030 38.960 ;
        RECT 133.580 38.560 135.580 38.600 ;
        RECT 133.230 38.320 135.930 38.560 ;
        RECT 133.190 37.560 135.970 38.320 ;
        RECT 133.190 37.360 133.420 37.560 ;
        RECT 135.740 37.360 135.970 37.560 ;
        RECT 133.580 37.080 135.580 37.310 ;
        RECT 134.030 36.760 135.530 37.080 ;
        RECT 136.230 37.010 139.030 38.960 ;
        RECT 139.730 38.940 141.230 39.260 ;
        RECT 139.680 38.710 141.680 38.940 ;
        RECT 139.730 38.660 141.230 38.710 ;
        RECT 139.290 38.460 139.520 38.660 ;
        RECT 141.840 38.460 142.070 38.660 ;
        RECT 139.290 37.860 142.070 38.460 ;
        RECT 139.290 37.700 139.520 37.860 ;
        RECT 141.840 37.700 142.070 37.860 ;
        RECT 142.230 37.760 143.030 39.260 ;
        RECT 143.730 44.060 150.630 45.260 ;
        RECT 143.730 42.260 144.030 44.060 ;
        RECT 144.930 43.740 146.730 43.910 ;
        RECT 144.725 43.510 148.725 43.740 ;
        RECT 144.290 43.260 144.520 43.460 ;
        RECT 144.930 43.410 146.730 43.510 ;
        RECT 144.290 43.160 144.530 43.260 ;
        RECT 147.730 43.160 148.030 43.310 ;
        RECT 148.930 43.260 149.160 43.460 ;
        RECT 148.830 43.160 149.160 43.260 ;
        RECT 144.290 42.660 149.160 43.160 ;
        RECT 144.290 42.500 144.520 42.660 ;
        RECT 148.930 42.500 149.160 42.660 ;
        RECT 144.725 42.360 148.725 42.450 ;
        RECT 149.330 42.360 150.630 44.060 ;
        RECT 144.725 42.260 150.630 42.360 ;
        RECT 143.730 40.660 150.630 42.260 ;
        RECT 143.730 38.960 144.030 40.660 ;
        RECT 144.725 40.510 148.725 40.660 ;
        RECT 144.290 40.360 144.520 40.460 ;
        RECT 148.930 40.360 149.160 40.460 ;
        RECT 144.290 39.500 149.160 40.360 ;
        RECT 144.330 39.260 149.130 39.500 ;
        RECT 144.725 39.220 148.725 39.260 ;
        RECT 143.730 38.930 144.050 38.960 ;
        RECT 149.330 38.930 150.630 40.660 ;
        RECT 143.730 38.360 150.630 38.930 ;
        RECT 139.680 37.160 141.680 37.650 ;
        RECT 142.230 37.260 147.130 37.760 ;
        RECT 141.130 37.110 141.630 37.160 ;
        RECT 136.230 36.960 139.080 37.010 ;
        RECT 142.230 36.960 143.530 37.260 ;
        RECT 136.230 36.760 143.530 36.960 ;
        RECT 144.180 36.940 145.830 37.110 ;
        RECT 132.230 36.360 143.530 36.760 ;
        RECT 144.130 36.710 146.130 36.940 ;
        RECT 144.230 36.660 145.830 36.710 ;
        RECT 143.740 36.560 143.970 36.660 ;
        RECT 146.290 36.610 146.520 36.660 ;
        RECT 146.230 36.560 146.530 36.610 ;
        RECT 132.230 36.060 139.030 36.360 ;
        RECT 132.230 33.960 132.930 36.060 ;
        RECT 133.580 35.660 135.580 35.700 ;
        RECT 133.230 35.610 135.930 35.660 ;
        RECT 133.130 35.420 135.930 35.610 ;
        RECT 133.130 34.660 135.970 35.420 ;
        RECT 133.130 34.610 133.530 34.660 ;
        RECT 133.130 34.470 133.420 34.610 ;
        RECT 133.190 34.460 133.420 34.470 ;
        RECT 135.740 34.460 135.970 34.660 ;
        RECT 133.580 34.180 135.580 34.410 ;
        RECT 136.230 34.210 139.030 36.060 ;
        RECT 139.730 36.040 141.230 36.360 ;
        RECT 139.680 35.810 141.680 36.040 ;
        RECT 139.730 35.760 141.230 35.810 ;
        RECT 139.290 35.560 139.520 35.760 ;
        RECT 141.840 35.560 142.070 35.760 ;
        RECT 139.290 34.960 142.070 35.560 ;
        RECT 139.290 34.800 139.520 34.960 ;
        RECT 141.840 34.800 142.070 34.960 ;
        RECT 142.230 35.060 143.530 36.360 ;
        RECT 143.730 36.410 144.080 36.560 ;
        RECT 146.130 36.410 146.530 36.560 ;
        RECT 143.730 35.960 146.530 36.410 ;
        RECT 143.730 35.860 144.130 35.960 ;
        RECT 146.130 35.860 146.530 35.960 ;
        RECT 143.740 35.700 143.970 35.860 ;
        RECT 146.230 35.810 146.530 35.860 ;
        RECT 144.380 35.710 145.930 35.810 ;
        RECT 144.130 35.650 145.930 35.710 ;
        RECT 146.290 35.700 146.520 35.810 ;
        RECT 144.130 35.420 146.130 35.650 ;
        RECT 144.130 35.260 145.930 35.420 ;
        RECT 146.830 35.060 147.130 37.260 ;
        RECT 139.680 34.520 141.680 34.750 ;
        RECT 139.680 34.410 141.630 34.520 ;
        RECT 142.230 34.460 147.130 35.060 ;
        RECT 147.510 34.530 150.630 38.360 ;
        RECT 142.230 34.260 143.130 34.460 ;
        RECT 142.180 34.210 143.130 34.260 ;
        RECT 134.030 33.960 135.530 34.180 ;
        RECT 136.230 33.960 143.130 34.210 ;
        RECT 124.630 32.390 126.380 33.660 ;
        RECT 132.230 33.460 143.130 33.960 ;
        RECT 132.130 32.960 143.030 33.460 ;
        RECT 148.880 33.260 150.630 34.530 ;
        RECT 132.130 32.710 139.030 32.960 ;
        RECT 139.730 32.740 141.230 32.960 ;
        RECT 132.130 32.660 133.080 32.710 ;
        RECT 132.130 32.460 133.030 32.660 ;
        RECT 124.630 28.560 127.750 32.390 ;
        RECT 128.130 31.860 133.030 32.460 ;
        RECT 133.630 32.400 135.580 32.510 ;
        RECT 133.580 32.170 135.580 32.400 ;
        RECT 128.130 29.660 128.430 31.860 ;
        RECT 129.330 31.500 131.130 31.660 ;
        RECT 129.130 31.270 131.130 31.500 ;
        RECT 128.740 31.110 128.970 31.220 ;
        RECT 129.330 31.210 131.130 31.270 ;
        RECT 129.330 31.110 130.880 31.210 ;
        RECT 128.730 31.060 129.030 31.110 ;
        RECT 131.290 31.060 131.520 31.220 ;
        RECT 128.730 30.960 129.130 31.060 ;
        RECT 131.130 30.960 131.530 31.060 ;
        RECT 128.730 30.510 131.530 30.960 ;
        RECT 128.730 30.360 129.130 30.510 ;
        RECT 131.180 30.360 131.530 30.510 ;
        RECT 131.730 30.560 133.030 31.860 ;
        RECT 133.190 31.960 133.420 32.120 ;
        RECT 135.740 31.960 135.970 32.120 ;
        RECT 133.190 31.360 135.970 31.960 ;
        RECT 133.190 31.160 133.420 31.360 ;
        RECT 135.740 31.160 135.970 31.360 ;
        RECT 134.030 31.110 135.530 31.160 ;
        RECT 133.580 30.880 135.580 31.110 ;
        RECT 134.030 30.560 135.530 30.880 ;
        RECT 136.230 30.860 139.030 32.710 ;
        RECT 139.680 32.510 141.680 32.740 ;
        RECT 139.290 32.260 139.520 32.460 ;
        RECT 141.840 32.450 142.070 32.460 ;
        RECT 141.840 32.310 142.130 32.450 ;
        RECT 141.730 32.260 142.130 32.310 ;
        RECT 139.290 31.500 142.130 32.260 ;
        RECT 139.330 31.310 142.130 31.500 ;
        RECT 139.330 31.260 142.030 31.310 ;
        RECT 139.680 31.220 141.680 31.260 ;
        RECT 142.330 30.860 143.030 32.960 ;
        RECT 136.230 30.560 143.030 30.860 ;
        RECT 128.730 30.310 129.030 30.360 ;
        RECT 128.740 30.260 128.970 30.310 ;
        RECT 131.290 30.260 131.520 30.360 ;
        RECT 129.430 30.210 131.030 30.260 ;
        RECT 129.130 29.980 131.130 30.210 ;
        RECT 131.730 30.160 143.030 30.560 ;
        RECT 129.430 29.810 131.080 29.980 ;
        RECT 131.730 29.960 139.030 30.160 ;
        RECT 131.730 29.660 133.030 29.960 ;
        RECT 136.180 29.910 139.030 29.960 ;
        RECT 133.630 29.760 134.130 29.810 ;
        RECT 128.130 29.160 133.030 29.660 ;
        RECT 133.580 29.270 135.580 29.760 ;
        RECT 124.630 27.990 131.530 28.560 ;
        RECT 124.630 26.260 125.930 27.990 ;
        RECT 131.210 27.960 131.530 27.990 ;
        RECT 126.535 27.660 130.535 27.700 ;
        RECT 126.130 27.420 130.930 27.660 ;
        RECT 126.100 26.560 130.970 27.420 ;
        RECT 126.100 26.460 126.330 26.560 ;
        RECT 130.740 26.460 130.970 26.560 ;
        RECT 126.535 26.260 130.535 26.410 ;
        RECT 131.230 26.260 131.530 27.960 ;
        RECT 124.630 24.660 131.530 26.260 ;
        RECT 124.630 24.560 130.535 24.660 ;
        RECT 124.630 22.860 125.930 24.560 ;
        RECT 126.535 24.470 130.535 24.560 ;
        RECT 126.100 24.260 126.330 24.420 ;
        RECT 130.740 24.260 130.970 24.420 ;
        RECT 126.100 23.760 130.970 24.260 ;
        RECT 126.100 23.660 126.430 23.760 ;
        RECT 126.100 23.460 126.330 23.660 ;
        RECT 127.230 23.610 127.530 23.760 ;
        RECT 130.730 23.660 130.970 23.760 ;
        RECT 128.530 23.410 130.330 23.510 ;
        RECT 130.740 23.460 130.970 23.660 ;
        RECT 126.535 23.180 130.535 23.410 ;
        RECT 128.530 23.010 130.330 23.180 ;
        RECT 131.230 22.860 131.530 24.660 ;
        RECT 124.630 21.660 131.530 22.860 ;
        RECT 132.230 27.660 133.030 29.160 ;
        RECT 133.190 29.060 133.420 29.220 ;
        RECT 135.740 29.060 135.970 29.220 ;
        RECT 133.190 28.460 135.970 29.060 ;
        RECT 133.190 28.260 133.420 28.460 ;
        RECT 135.740 28.260 135.970 28.460 ;
        RECT 134.030 28.210 135.530 28.260 ;
        RECT 133.580 27.980 135.580 28.210 ;
        RECT 134.030 27.660 135.530 27.980 ;
        RECT 136.230 27.960 139.030 29.910 ;
        RECT 139.730 29.840 141.230 30.160 ;
        RECT 139.680 29.610 141.680 29.840 ;
        RECT 139.290 29.360 139.520 29.560 ;
        RECT 141.840 29.360 142.070 29.560 ;
        RECT 139.290 28.600 142.070 29.360 ;
        RECT 139.330 28.360 142.030 28.600 ;
        RECT 139.680 28.320 141.680 28.360 ;
        RECT 142.230 27.960 143.030 30.160 ;
        RECT 136.230 27.660 143.030 27.960 ;
        RECT 132.230 27.260 143.030 27.660 ;
        RECT 132.230 26.960 139.030 27.260 ;
        RECT 132.230 24.760 133.030 26.960 ;
        RECT 133.580 26.560 135.580 26.600 ;
        RECT 133.230 26.320 135.930 26.560 ;
        RECT 133.190 25.560 135.970 26.320 ;
        RECT 133.190 25.360 133.420 25.560 ;
        RECT 135.740 25.360 135.970 25.560 ;
        RECT 133.580 25.080 135.580 25.310 ;
        RECT 134.030 24.760 135.530 25.080 ;
        RECT 136.230 25.010 139.030 26.960 ;
        RECT 139.730 26.940 141.230 27.260 ;
        RECT 139.680 26.710 141.680 26.940 ;
        RECT 139.730 26.660 141.230 26.710 ;
        RECT 139.290 26.460 139.520 26.660 ;
        RECT 141.840 26.460 142.070 26.660 ;
        RECT 139.290 25.860 142.070 26.460 ;
        RECT 139.290 25.700 139.520 25.860 ;
        RECT 141.840 25.700 142.070 25.860 ;
        RECT 142.230 25.760 143.030 27.260 ;
        RECT 143.730 32.060 150.630 33.260 ;
        RECT 143.730 30.260 144.030 32.060 ;
        RECT 144.930 31.740 146.730 31.910 ;
        RECT 144.725 31.510 148.725 31.740 ;
        RECT 144.290 31.260 144.520 31.460 ;
        RECT 144.930 31.410 146.730 31.510 ;
        RECT 144.290 31.160 144.530 31.260 ;
        RECT 147.730 31.160 148.030 31.310 ;
        RECT 148.930 31.260 149.160 31.460 ;
        RECT 148.830 31.160 149.160 31.260 ;
        RECT 144.290 30.660 149.160 31.160 ;
        RECT 144.290 30.500 144.520 30.660 ;
        RECT 148.930 30.500 149.160 30.660 ;
        RECT 144.725 30.360 148.725 30.450 ;
        RECT 149.330 30.360 150.630 32.060 ;
        RECT 144.725 30.260 150.630 30.360 ;
        RECT 143.730 28.660 150.630 30.260 ;
        RECT 143.730 26.960 144.030 28.660 ;
        RECT 144.725 28.510 148.725 28.660 ;
        RECT 144.290 28.360 144.520 28.460 ;
        RECT 148.930 28.360 149.160 28.460 ;
        RECT 144.290 27.500 149.160 28.360 ;
        RECT 144.330 27.260 149.130 27.500 ;
        RECT 144.725 27.220 148.725 27.260 ;
        RECT 143.730 26.930 144.050 26.960 ;
        RECT 149.330 26.930 150.630 28.660 ;
        RECT 143.730 26.360 150.630 26.930 ;
        RECT 139.680 25.160 141.680 25.650 ;
        RECT 142.230 25.260 147.130 25.760 ;
        RECT 141.130 25.110 141.630 25.160 ;
        RECT 136.230 24.960 139.080 25.010 ;
        RECT 142.230 24.960 143.530 25.260 ;
        RECT 136.230 24.760 143.530 24.960 ;
        RECT 144.180 24.940 145.830 25.110 ;
        RECT 132.230 24.360 143.530 24.760 ;
        RECT 144.130 24.710 146.130 24.940 ;
        RECT 144.230 24.660 145.830 24.710 ;
        RECT 143.740 24.560 143.970 24.660 ;
        RECT 146.290 24.610 146.520 24.660 ;
        RECT 146.230 24.560 146.530 24.610 ;
        RECT 132.230 24.060 139.030 24.360 ;
        RECT 132.230 21.960 132.930 24.060 ;
        RECT 133.580 23.660 135.580 23.700 ;
        RECT 133.230 23.610 135.930 23.660 ;
        RECT 133.130 23.420 135.930 23.610 ;
        RECT 133.130 22.660 135.970 23.420 ;
        RECT 133.130 22.610 133.530 22.660 ;
        RECT 133.130 22.470 133.420 22.610 ;
        RECT 133.190 22.460 133.420 22.470 ;
        RECT 135.740 22.460 135.970 22.660 ;
        RECT 133.580 22.180 135.580 22.410 ;
        RECT 136.230 22.210 139.030 24.060 ;
        RECT 139.730 24.040 141.230 24.360 ;
        RECT 139.680 23.810 141.680 24.040 ;
        RECT 139.730 23.760 141.230 23.810 ;
        RECT 139.290 23.560 139.520 23.760 ;
        RECT 141.840 23.560 142.070 23.760 ;
        RECT 139.290 22.960 142.070 23.560 ;
        RECT 139.290 22.800 139.520 22.960 ;
        RECT 141.840 22.800 142.070 22.960 ;
        RECT 142.230 23.060 143.530 24.360 ;
        RECT 143.730 24.410 144.080 24.560 ;
        RECT 146.130 24.410 146.530 24.560 ;
        RECT 143.730 23.960 146.530 24.410 ;
        RECT 143.730 23.860 144.130 23.960 ;
        RECT 146.130 23.860 146.530 23.960 ;
        RECT 143.740 23.700 143.970 23.860 ;
        RECT 146.230 23.810 146.530 23.860 ;
        RECT 144.380 23.710 145.930 23.810 ;
        RECT 144.130 23.650 145.930 23.710 ;
        RECT 146.290 23.700 146.520 23.810 ;
        RECT 144.130 23.420 146.130 23.650 ;
        RECT 144.130 23.260 145.930 23.420 ;
        RECT 146.830 23.060 147.130 25.260 ;
        RECT 139.680 22.520 141.680 22.750 ;
        RECT 139.680 22.410 141.630 22.520 ;
        RECT 142.230 22.460 147.130 23.060 ;
        RECT 147.510 22.530 150.630 26.360 ;
        RECT 142.230 22.260 143.130 22.460 ;
        RECT 142.180 22.210 143.130 22.260 ;
        RECT 134.030 21.960 135.530 22.180 ;
        RECT 136.230 21.960 143.130 22.210 ;
        RECT 124.630 21.460 126.380 21.660 ;
        RECT 132.230 21.460 143.130 21.960 ;
        RECT 148.880 21.460 150.630 22.530 ;
        RECT 124.630 20.460 126.130 21.460 ;
        RECT 132.130 20.960 143.130 21.460 ;
        RECT 148.885 20.960 150.630 21.460 ;
        RECT 151.130 20.960 154.130 72.160 ;
        RECT 124.630 20.060 131.130 20.460 ;
        RECT 121.730 19.960 131.130 20.060 ;
        RECT 132.130 19.960 146.930 20.960 ;
        RECT 121.730 19.880 131.530 19.960 ;
        RECT 119.360 19.760 131.530 19.880 ;
        RECT 116.780 19.560 131.530 19.760 ;
        RECT 116.780 19.360 143.330 19.560 ;
        RECT 116.780 19.160 143.430 19.360 ;
        RECT 116.780 18.760 132.030 19.160 ;
        RECT 132.480 19.090 143.430 19.160 ;
        RECT 135.130 19.060 143.430 19.090 ;
        RECT 116.780 17.360 131.930 18.760 ;
        RECT 132.730 18.750 136.630 18.760 ;
        RECT 132.730 18.520 136.735 18.750 ;
        RECT 132.300 18.160 132.530 18.470 ;
        RECT 132.730 18.160 136.630 18.520 ;
        RECT 136.940 18.360 137.170 18.470 ;
        RECT 137.850 18.360 138.080 18.470 ;
        RECT 136.940 18.160 138.080 18.360 ;
        RECT 138.230 18.310 142.330 18.860 ;
        RECT 142.490 18.160 142.720 18.470 ;
        RECT 132.300 17.760 142.720 18.160 ;
        RECT 132.300 17.510 132.530 17.760 ;
        RECT 136.940 17.660 142.720 17.760 ;
        RECT 136.940 17.560 138.080 17.660 ;
        RECT 136.940 17.510 137.170 17.560 ;
        RECT 137.850 17.510 138.080 17.560 ;
        RECT 142.490 17.510 142.720 17.660 ;
        RECT 116.780 16.960 132.030 17.360 ;
        RECT 132.735 17.230 136.735 17.460 ;
        RECT 138.285 17.230 142.285 17.460 ;
        RECT 133.230 16.960 136.330 17.230 ;
        RECT 138.430 16.960 142.130 17.230 ;
        RECT 142.930 16.960 143.430 19.060 ;
        RECT 144.030 17.760 146.930 19.960 ;
        RECT 148.885 19.460 154.130 20.960 ;
        RECT 149.130 16.960 154.130 19.460 ;
        RECT 116.780 15.160 154.130 16.960 ;
        RECT 116.780 14.460 138.030 15.160 ;
        RECT 141.930 14.460 154.130 15.160 ;
        RECT 116.780 12.380 124.050 14.460 ;
        RECT 134.030 2.240 136.270 6.900 ;
      LAYER met2 ;
        RECT 133.535 95.190 134.125 95.690 ;
        RECT 133.580 74.110 134.080 95.190 ;
        RECT 121.680 73.610 134.080 74.110 ;
        RECT 121.680 30.960 122.180 73.610 ;
        RECT 135.180 73.110 135.680 94.685 ;
        RECT 136.035 93.010 136.625 93.510 ;
        RECT 122.680 72.610 135.680 73.110 ;
        RECT 136.080 91.300 136.580 93.010 ;
        RECT 136.080 90.690 136.560 91.300 ;
        RECT 122.680 42.960 123.180 72.610 ;
        RECT 136.080 71.910 136.580 90.690 ;
        RECT 136.960 89.920 137.870 91.680 ;
        RECT 123.680 71.410 136.580 71.910 ;
        RECT 123.680 54.960 124.180 71.410 ;
        RECT 137.080 71.110 137.580 89.920 ;
        RECT 138.235 88.820 138.825 89.320 ;
        RECT 124.780 70.610 137.580 71.110 ;
        RECT 138.280 71.210 138.780 88.820 ;
        RECT 139.280 72.210 139.780 87.020 ;
        RECT 140.280 73.410 140.780 84.535 ;
        RECT 141.335 78.660 141.925 79.160 ;
        RECT 141.380 74.210 141.880 78.660 ;
        RECT 143.430 74.210 146.830 74.220 ;
        RECT 141.380 73.710 154.130 74.210 ;
        RECT 143.430 73.410 146.830 73.420 ;
        RECT 140.280 72.910 153.180 73.410 ;
        RECT 143.430 72.900 146.830 72.910 ;
        RECT 139.280 71.710 152.280 72.210 ;
        RECT 138.280 70.710 151.180 71.210 ;
        RECT 124.780 67.060 125.280 70.610 ;
        RECT 126.825 70.260 147.535 70.265 ;
        RECT 126.825 69.860 148.430 70.260 ;
        RECT 150.180 69.910 151.180 70.710 ;
        RECT 126.825 69.855 147.535 69.860 ;
        RECT 126.930 69.460 127.730 69.855 ;
        RECT 147.800 69.460 148.430 69.860 ;
        RECT 126.830 68.460 127.830 69.460 ;
        RECT 124.630 66.360 125.330 67.060 ;
        RECT 127.130 63.360 127.630 68.460 ;
        RECT 129.830 67.560 131.130 69.460 ;
        RECT 129.430 67.260 131.130 67.560 ;
        RECT 131.730 68.110 135.030 68.560 ;
        RECT 129.430 67.210 130.730 67.260 ;
        RECT 128.680 66.360 129.080 67.060 ;
        RECT 131.730 66.260 132.230 68.110 ;
        RECT 129.330 65.660 132.230 66.260 ;
        RECT 132.480 65.260 134.280 65.860 ;
        RECT 132.480 63.360 132.980 65.260 ;
        RECT 134.430 65.060 134.830 67.960 ;
        RECT 133.630 64.460 135.730 65.060 ;
        RECT 127.130 62.760 132.980 63.360 ;
        RECT 127.130 62.660 127.630 62.760 ;
        RECT 134.430 62.260 134.830 64.460 ;
        RECT 133.730 61.660 135.730 62.260 ;
        RECT 127.130 58.460 127.630 60.260 ;
        RECT 128.130 59.360 133.730 59.860 ;
        RECT 134.430 59.360 134.830 61.660 ;
        RECT 128.130 58.760 135.630 59.360 ;
        RECT 128.130 58.660 133.730 58.760 ;
        RECT 132.330 58.460 133.730 58.660 ;
        RECT 126.830 56.460 127.830 58.460 ;
        RECT 124.630 54.960 125.230 55.060 ;
        RECT 123.680 54.460 125.230 54.960 ;
        RECT 124.630 54.360 125.230 54.460 ;
        RECT 127.130 51.360 127.630 56.460 ;
        RECT 129.830 55.560 131.130 57.460 ;
        RECT 129.430 55.260 131.130 55.560 ;
        RECT 131.730 56.110 135.030 56.560 ;
        RECT 129.430 55.210 130.730 55.260 ;
        RECT 128.680 54.360 129.080 55.060 ;
        RECT 131.730 54.260 132.230 56.110 ;
        RECT 129.330 53.660 132.230 54.260 ;
        RECT 132.480 53.260 134.280 53.860 ;
        RECT 132.480 51.360 132.980 53.260 ;
        RECT 134.430 53.060 134.830 55.960 ;
        RECT 133.630 52.460 135.730 53.060 ;
        RECT 127.130 50.760 132.980 51.360 ;
        RECT 127.130 50.660 127.630 50.760 ;
        RECT 134.430 50.260 134.830 52.460 ;
        RECT 133.730 49.660 135.730 50.260 ;
        RECT 127.130 46.460 127.630 48.260 ;
        RECT 128.130 47.360 133.730 47.860 ;
        RECT 134.430 47.360 134.830 49.660 ;
        RECT 128.130 46.760 135.630 47.360 ;
        RECT 128.130 46.660 133.730 46.760 ;
        RECT 132.330 46.460 133.730 46.660 ;
        RECT 126.830 44.460 127.830 46.460 ;
        RECT 124.705 42.960 125.155 42.980 ;
        RECT 122.680 42.460 125.180 42.960 ;
        RECT 124.705 42.440 125.155 42.460 ;
        RECT 127.130 39.360 127.630 44.460 ;
        RECT 129.830 43.560 131.130 45.460 ;
        RECT 129.430 43.260 131.130 43.560 ;
        RECT 131.730 44.110 135.030 44.560 ;
        RECT 129.430 43.210 130.730 43.260 ;
        RECT 128.680 42.360 129.080 43.060 ;
        RECT 131.730 42.260 132.230 44.110 ;
        RECT 129.330 41.660 132.230 42.260 ;
        RECT 132.480 41.260 134.280 41.860 ;
        RECT 132.480 39.360 132.980 41.260 ;
        RECT 134.430 41.060 134.830 43.960 ;
        RECT 133.630 40.460 135.730 41.060 ;
        RECT 127.130 38.760 132.980 39.360 ;
        RECT 127.130 38.660 127.630 38.760 ;
        RECT 134.430 38.260 134.830 40.460 ;
        RECT 133.730 37.660 135.730 38.260 ;
        RECT 127.130 34.460 127.630 36.260 ;
        RECT 128.130 35.360 133.730 35.860 ;
        RECT 134.430 35.360 134.830 37.660 ;
        RECT 128.130 34.760 135.630 35.360 ;
        RECT 128.130 34.660 133.730 34.760 ;
        RECT 132.330 34.460 133.730 34.660 ;
        RECT 126.830 32.460 127.830 34.460 ;
        RECT 124.805 30.960 125.255 30.980 ;
        RECT 121.680 30.460 125.280 30.960 ;
        RECT 124.805 30.440 125.255 30.460 ;
        RECT 127.130 27.360 127.630 32.460 ;
        RECT 129.830 31.560 131.130 33.460 ;
        RECT 129.430 31.260 131.130 31.560 ;
        RECT 131.730 32.110 135.030 32.560 ;
        RECT 129.430 31.210 130.730 31.260 ;
        RECT 128.680 30.360 129.080 31.060 ;
        RECT 131.730 30.260 132.230 32.110 ;
        RECT 129.330 29.660 132.230 30.260 ;
        RECT 132.480 29.260 134.280 29.860 ;
        RECT 132.480 27.360 132.980 29.260 ;
        RECT 134.430 29.060 134.830 31.960 ;
        RECT 133.630 28.460 135.730 29.060 ;
        RECT 127.130 26.760 132.980 27.360 ;
        RECT 127.130 26.660 127.630 26.760 ;
        RECT 134.430 26.260 134.830 28.460 ;
        RECT 133.730 25.660 135.730 26.260 ;
        RECT 127.130 22.460 127.630 24.260 ;
        RECT 128.130 23.360 133.730 23.860 ;
        RECT 134.430 23.360 134.830 25.660 ;
        RECT 128.130 22.760 135.630 23.360 ;
        RECT 128.130 22.660 133.730 22.760 ;
        RECT 132.330 22.460 133.730 22.660 ;
        RECT 126.630 20.960 128.130 22.460 ;
        RECT 119.360 19.760 123.700 19.880 ;
        RECT 116.780 12.380 124.050 19.760 ;
        RECT 126.870 8.205 128.040 20.960 ;
        RECT 136.630 19.960 138.630 69.460 ;
        RECT 147.430 68.460 148.430 69.460 ;
        RECT 141.530 68.260 142.930 68.460 ;
        RECT 141.530 68.160 147.130 68.260 ;
        RECT 139.630 67.560 147.130 68.160 ;
        RECT 140.430 65.260 140.830 67.560 ;
        RECT 141.530 67.060 147.130 67.560 ;
        RECT 147.630 66.660 148.130 68.460 ;
        RECT 139.530 64.660 141.530 65.260 ;
        RECT 140.430 62.460 140.830 64.660 ;
        RECT 147.630 64.160 148.130 64.260 ;
        RECT 142.280 63.560 148.130 64.160 ;
        RECT 139.530 61.860 141.630 62.460 ;
        RECT 140.430 58.960 140.830 61.860 ;
        RECT 142.280 61.660 142.780 63.560 ;
        RECT 140.980 61.060 142.780 61.660 ;
        RECT 143.030 60.660 145.930 61.260 ;
        RECT 143.030 58.810 143.530 60.660 ;
        RECT 146.180 59.860 146.580 60.560 ;
        RECT 144.530 59.660 145.830 59.710 ;
        RECT 140.230 58.360 143.530 58.810 ;
        RECT 144.130 59.360 145.830 59.660 ;
        RECT 144.130 57.460 145.430 59.360 ;
        RECT 147.630 58.460 148.130 63.560 ;
        RECT 150.680 60.560 151.180 69.910 ;
        RECT 150.130 59.760 151.230 60.560 ;
        RECT 147.430 56.460 148.430 58.460 ;
        RECT 141.530 56.260 142.930 56.460 ;
        RECT 141.530 56.160 147.130 56.260 ;
        RECT 139.630 55.560 147.130 56.160 ;
        RECT 140.430 53.260 140.830 55.560 ;
        RECT 141.530 55.060 147.130 55.560 ;
        RECT 147.630 54.660 148.130 56.460 ;
        RECT 139.530 52.660 141.530 53.260 ;
        RECT 140.430 50.460 140.830 52.660 ;
        RECT 147.630 52.160 148.130 52.260 ;
        RECT 142.280 51.560 148.130 52.160 ;
        RECT 139.530 49.860 141.630 50.460 ;
        RECT 140.430 46.960 140.830 49.860 ;
        RECT 142.280 49.660 142.780 51.560 ;
        RECT 140.980 49.060 142.780 49.660 ;
        RECT 143.030 48.660 145.930 49.260 ;
        RECT 143.030 46.810 143.530 48.660 ;
        RECT 146.180 47.860 146.580 48.560 ;
        RECT 144.530 47.660 145.830 47.710 ;
        RECT 140.230 46.360 143.530 46.810 ;
        RECT 144.130 47.360 145.830 47.660 ;
        RECT 144.130 45.460 145.430 47.360 ;
        RECT 147.630 46.460 148.130 51.560 ;
        RECT 151.780 48.410 152.280 71.710 ;
        RECT 150.180 47.910 152.280 48.410 ;
        RECT 147.430 44.460 148.430 46.460 ;
        RECT 141.530 44.260 142.930 44.460 ;
        RECT 141.530 44.160 147.130 44.260 ;
        RECT 139.630 43.560 147.130 44.160 ;
        RECT 140.430 41.260 140.830 43.560 ;
        RECT 141.530 43.060 147.130 43.560 ;
        RECT 147.630 42.660 148.130 44.460 ;
        RECT 139.530 40.660 141.530 41.260 ;
        RECT 140.430 38.460 140.830 40.660 ;
        RECT 147.630 40.160 148.130 40.260 ;
        RECT 142.280 39.560 148.130 40.160 ;
        RECT 139.530 37.860 141.630 38.460 ;
        RECT 140.430 34.960 140.830 37.860 ;
        RECT 142.280 37.660 142.780 39.560 ;
        RECT 140.980 37.060 142.780 37.660 ;
        RECT 143.030 36.660 145.930 37.260 ;
        RECT 143.030 34.810 143.530 36.660 ;
        RECT 146.180 35.860 146.580 36.560 ;
        RECT 144.530 35.660 145.830 35.710 ;
        RECT 140.230 34.360 143.530 34.810 ;
        RECT 144.130 35.360 145.830 35.660 ;
        RECT 144.130 33.460 145.430 35.360 ;
        RECT 147.630 34.460 148.130 39.560 ;
        RECT 152.680 36.410 153.180 72.910 ;
        RECT 150.135 35.910 153.180 36.410 ;
        RECT 152.680 35.860 153.180 35.910 ;
        RECT 147.430 32.460 148.430 34.460 ;
        RECT 141.530 32.260 142.930 32.460 ;
        RECT 141.530 32.160 147.130 32.260 ;
        RECT 139.630 31.560 147.130 32.160 ;
        RECT 140.430 29.260 140.830 31.560 ;
        RECT 141.530 31.060 147.130 31.560 ;
        RECT 147.630 30.660 148.130 32.460 ;
        RECT 139.530 28.660 141.530 29.260 ;
        RECT 140.430 26.460 140.830 28.660 ;
        RECT 147.630 28.160 148.130 28.260 ;
        RECT 142.280 27.560 148.130 28.160 ;
        RECT 139.530 25.860 141.630 26.460 ;
        RECT 140.430 22.960 140.830 25.860 ;
        RECT 142.280 25.660 142.780 27.560 ;
        RECT 140.980 25.060 142.780 25.660 ;
        RECT 143.030 24.660 145.930 25.260 ;
        RECT 143.030 22.810 143.530 24.660 ;
        RECT 146.180 23.860 146.580 24.560 ;
        RECT 144.530 23.660 145.830 23.710 ;
        RECT 140.230 22.360 143.530 22.810 ;
        RECT 144.130 23.360 145.830 23.660 ;
        RECT 144.130 21.460 145.430 23.360 ;
        RECT 147.630 22.460 148.130 27.560 ;
        RECT 150.135 24.260 152.230 24.410 ;
        RECT 153.680 24.285 154.130 73.710 ;
        RECT 153.430 24.260 154.130 24.285 ;
        RECT 150.135 23.910 154.130 24.260 ;
        RECT 150.205 23.860 154.130 23.910 ;
        RECT 150.205 23.835 152.630 23.860 ;
        RECT 147.130 20.960 148.630 22.460 ;
        RECT 137.030 18.660 137.830 19.960 ;
        RECT 138.530 18.760 141.530 18.860 ;
        RECT 136.930 17.360 138.030 18.660 ;
        RECT 138.380 18.360 142.180 18.760 ;
        RECT 138.530 9.940 141.530 18.360 ;
        RECT 144.710 18.350 145.710 19.120 ;
        RECT 147.330 16.760 148.530 20.960 ;
        RECT 147.230 14.460 148.530 16.760 ;
        RECT 111.885 7.035 128.040 8.205 ;
        RECT 138.540 7.725 141.525 9.940 ;
        RECT 147.700 8.780 148.300 14.460 ;
        RECT 147.725 8.760 148.275 8.780 ;
        RECT 111.885 6.645 113.055 7.035 ;
        RECT 111.840 5.475 113.100 6.645 ;
        RECT 133.660 4.740 141.525 7.725 ;
        RECT 133.660 1.620 136.840 4.740 ;
        RECT 133.780 1.080 136.840 1.620 ;
      LAYER met3 ;
        RECT 133.555 95.690 134.105 95.715 ;
        RECT 147.310 95.690 147.810 95.720 ;
        RECT 133.555 95.190 147.810 95.690 ;
        RECT 133.555 95.165 134.105 95.190 ;
        RECT 147.310 95.160 147.810 95.190 ;
        RECT 135.155 94.640 135.705 94.665 ;
        RECT 143.450 94.640 143.950 94.670 ;
        RECT 135.155 94.140 143.950 94.640 ;
        RECT 135.155 94.115 135.705 94.140 ;
        RECT 143.450 94.110 143.950 94.140 ;
        RECT 136.055 93.510 136.605 93.535 ;
        RECT 140.170 93.510 140.670 93.540 ;
        RECT 136.055 93.010 140.670 93.510 ;
        RECT 136.055 92.985 136.605 93.010 ;
        RECT 140.170 92.980 140.670 93.010 ;
        RECT 136.770 90.030 138.100 91.790 ;
        RECT 132.770 89.320 133.270 89.350 ;
        RECT 138.255 89.320 138.805 89.345 ;
        RECT 132.770 88.820 138.805 89.320 ;
        RECT 132.770 88.790 133.270 88.820 ;
        RECT 138.255 88.795 138.805 88.820 ;
        RECT 129.240 86.890 129.740 86.920 ;
        RECT 139.255 86.890 139.805 86.915 ;
        RECT 129.240 86.390 139.805 86.890 ;
        RECT 129.240 86.360 129.740 86.390 ;
        RECT 139.255 86.365 139.805 86.390 ;
        RECT 125.450 84.490 125.950 84.520 ;
        RECT 140.255 84.490 140.805 84.515 ;
        RECT 125.450 83.990 140.805 84.490 ;
        RECT 125.450 83.960 125.950 83.990 ;
        RECT 140.255 83.965 140.805 83.990 ;
        RECT 122.000 79.160 122.500 79.190 ;
        RECT 141.355 79.160 141.905 79.185 ;
        RECT 122.000 78.660 141.905 79.160 ;
        RECT 122.000 78.630 122.500 78.660 ;
        RECT 141.355 78.635 141.905 78.660 ;
        RECT 129.630 67.960 138.630 69.460 ;
        RECT 136.630 67.460 138.630 67.960 ;
        RECT 124.630 66.960 125.130 67.060 ;
        RECT 128.130 66.960 129.130 67.460 ;
        RECT 124.630 66.460 129.130 66.960 ;
        RECT 124.630 66.360 125.130 66.460 ;
        RECT 128.130 65.960 129.130 66.460 ;
        RECT 146.130 60.460 147.130 60.960 ;
        RECT 150.130 60.460 150.630 60.560 ;
        RECT 146.130 60.410 150.630 60.460 ;
        RECT 146.130 59.960 150.655 60.410 ;
        RECT 146.130 59.460 147.130 59.960 ;
        RECT 150.130 59.910 150.655 59.960 ;
        RECT 150.130 59.860 150.630 59.910 ;
        RECT 136.630 57.460 145.630 58.960 ;
        RECT 129.630 55.960 138.630 57.460 ;
        RECT 124.630 54.960 125.130 55.060 ;
        RECT 128.130 54.960 129.130 55.460 ;
        RECT 124.630 54.460 129.130 54.960 ;
        RECT 124.630 54.360 125.130 54.460 ;
        RECT 128.130 53.960 129.130 54.460 ;
        RECT 146.130 48.460 147.130 48.960 ;
        RECT 150.130 48.460 150.630 48.560 ;
        RECT 146.130 48.410 150.630 48.460 ;
        RECT 146.130 47.960 150.655 48.410 ;
        RECT 146.130 47.460 147.130 47.960 ;
        RECT 150.130 47.910 150.655 47.960 ;
        RECT 150.130 47.860 150.630 47.910 ;
        RECT 136.630 45.460 145.630 46.960 ;
        RECT 129.630 43.960 138.630 45.460 ;
        RECT 124.630 42.960 125.130 43.060 ;
        RECT 128.130 42.960 129.130 43.460 ;
        RECT 124.630 42.460 129.130 42.960 ;
        RECT 124.630 42.360 125.130 42.460 ;
        RECT 128.130 41.960 129.130 42.460 ;
        RECT 146.130 36.460 147.130 36.960 ;
        RECT 150.130 36.460 150.630 36.560 ;
        RECT 146.130 36.435 150.630 36.460 ;
        RECT 146.130 35.960 150.705 36.435 ;
        RECT 146.130 35.460 147.130 35.960 ;
        RECT 150.130 35.885 150.705 35.960 ;
        RECT 150.130 35.860 150.630 35.885 ;
        RECT 136.630 33.460 145.630 34.960 ;
        RECT 129.630 31.960 138.630 33.460 ;
        RECT 124.630 30.960 125.130 31.060 ;
        RECT 128.130 30.960 129.130 31.460 ;
        RECT 124.630 30.460 129.130 30.960 ;
        RECT 124.630 30.360 125.130 30.460 ;
        RECT 128.130 29.960 129.130 30.460 ;
        RECT 146.130 24.460 147.130 24.960 ;
        RECT 150.130 24.460 150.630 24.560 ;
        RECT 146.130 24.435 150.630 24.460 ;
        RECT 146.130 23.960 150.705 24.435 ;
        RECT 146.130 23.460 147.130 23.960 ;
        RECT 150.130 23.885 150.705 23.960 ;
        RECT 150.130 23.860 150.630 23.885 ;
        RECT 136.630 22.960 138.630 23.460 ;
        RECT 136.630 21.460 145.630 22.960 ;
        RECT 43.105 19.800 44.595 19.825 ;
        RECT 43.100 19.760 123.360 19.800 ;
        RECT 43.100 18.300 124.050 19.760 ;
        RECT 144.660 18.375 145.760 19.095 ;
        RECT 43.105 18.275 44.595 18.300 ;
        RECT 116.780 12.380 124.050 18.300 ;
        RECT 111.860 5.555 113.080 6.670 ;
        RECT 111.855 4.385 113.085 5.555 ;
        RECT 133.780 1.080 136.840 7.610 ;
        RECT 147.700 6.330 148.300 9.380 ;
        RECT 147.705 6.305 148.295 6.330 ;
      LAYER met4 ;
        RECT 3.980 224.760 3.990 225.060 ;
        RECT 4.290 224.760 7.670 225.060 ;
        RECT 7.970 224.760 11.350 225.060 ;
        RECT 11.650 224.760 15.030 225.060 ;
        RECT 15.330 224.760 18.710 225.060 ;
        RECT 19.010 224.760 22.390 225.060 ;
        RECT 22.690 224.760 26.070 225.060 ;
        RECT 26.370 224.760 29.750 225.060 ;
        RECT 30.050 224.760 33.430 225.060 ;
        RECT 33.730 224.760 37.110 225.060 ;
        RECT 37.410 224.760 40.790 225.060 ;
        RECT 41.090 224.760 44.470 225.060 ;
        RECT 44.770 224.760 48.150 225.060 ;
        RECT 48.450 224.760 51.830 225.060 ;
        RECT 52.130 224.760 55.510 225.060 ;
        RECT 55.810 224.760 59.190 225.060 ;
        RECT 59.490 224.760 62.870 225.060 ;
        RECT 63.170 224.760 66.550 225.060 ;
        RECT 66.850 224.760 70.230 225.060 ;
        RECT 70.530 224.760 73.910 225.060 ;
        RECT 74.210 224.760 77.590 225.060 ;
        RECT 77.890 224.760 81.270 225.060 ;
        RECT 81.570 224.760 84.950 225.060 ;
        RECT 85.250 224.760 88.630 225.060 ;
        RECT 49.000 220.760 50.500 224.760 ;
        RECT 121.750 96.550 122.050 224.760 ;
        RECT 125.430 96.600 125.730 224.760 ;
        RECT 121.730 76.980 122.580 96.550 ;
        RECT 125.320 80.760 126.170 96.600 ;
        RECT 129.110 96.520 129.410 224.760 ;
        RECT 132.790 96.550 133.090 224.760 ;
        RECT 136.470 96.570 136.770 224.760 ;
        RECT 129.020 80.760 129.870 96.520 ;
        RECT 132.630 81.590 133.480 96.550 ;
        RECT 136.280 91.790 137.130 96.570 ;
        RECT 140.150 96.440 140.450 224.760 ;
        RECT 143.830 96.440 144.130 224.760 ;
        RECT 136.280 91.160 138.100 91.790 ;
        RECT 136.280 90.090 138.120 91.160 ;
        RECT 136.280 90.030 138.100 90.090 ;
        RECT 136.280 89.950 137.990 90.030 ;
        RECT 132.630 80.760 133.460 81.590 ;
        RECT 136.280 80.760 137.130 89.950 ;
        RECT 140.110 80.760 140.960 96.440 ;
        RECT 143.510 94.645 144.360 96.440 ;
        RECT 147.510 96.100 147.810 224.760 ;
        RECT 143.445 94.135 144.360 94.645 ;
        RECT 143.450 92.760 144.360 94.135 ;
        RECT 125.320 80.260 126.230 80.760 ;
        RECT 128.910 80.260 129.890 80.760 ;
        RECT 132.570 80.260 133.460 80.760 ;
        RECT 136.140 80.260 137.210 80.760 ;
        RECT 140.000 80.260 141.060 80.760 ;
        RECT 125.320 77.030 126.170 80.260 ;
        RECT 121.750 76.940 122.050 76.980 ;
        RECT 125.430 76.940 125.730 77.030 ;
        RECT 129.020 76.950 129.870 80.260 ;
        RECT 132.630 80.170 133.460 80.260 ;
        RECT 132.630 76.980 133.480 80.170 ;
        RECT 136.280 77.000 137.130 80.260 ;
        RECT 136.470 76.960 136.770 77.000 ;
        RECT 140.110 76.870 140.960 80.260 ;
        RECT 143.510 76.870 144.360 92.760 ;
        RECT 143.830 76.580 144.130 76.870 ;
        RECT 147.180 76.530 148.030 96.100 ;
        RECT 147.510 76.440 147.810 76.530 ;
        RECT 50.500 42.440 108.320 43.940 ;
        RECT 2.500 18.300 44.600 19.800 ;
        RECT 106.630 11.360 108.130 42.440 ;
        RECT 119.360 19.760 123.700 19.880 ;
        RECT 116.780 12.380 124.050 19.760 ;
        RECT 144.220 17.880 146.850 20.230 ;
        RECT 144.590 11.360 146.090 17.880 ;
        RECT 106.630 9.860 146.090 11.360 ;
        RECT 111.880 4.380 113.060 5.560 ;
        RECT 111.885 2.495 113.055 4.380 ;
        RECT 112.400 1.000 113.000 2.495 ;
        RECT 133.780 1.080 136.840 7.610 ;
        RECT 147.700 3.200 148.300 6.930 ;
        RECT 147.700 2.600 157.160 3.200 ;
        RECT 134.480 1.000 135.080 1.080 ;
        RECT 156.560 1.000 157.160 2.600 ;
  END
END tt_um_emilian_rf_playground
END LIBRARY

