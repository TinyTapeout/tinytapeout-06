VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_obriensp_be8
  CLASS BLOCK ;
  FOREIGN tt_um_obriensp_be8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 111.520 ;
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 146.280 2.480 147.880 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 95.080 10.000 96.680 107.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 43.880 10.000 45.480 107.700 ;
    END
  END VGND
  PIN VPWR
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 143.180 10.000 144.780 107.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 120.680 10.000 122.280 107.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 69.480 10.000 71.080 107.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 18.280 10.000 19.880 107.700 ;
    END
  END VPWR
  PIN clk
    ANTENNAGATEAREA 0.852000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 154.870 90.940 155.170 111.520 ;
    END
  END clk
  PIN ena
    PORT
      LAYER met4 ;
        RECT 158.550 110.520 158.850 111.520 ;
    END
  END ena
  PIN rst_n
    ANTENNAGATEAREA 0.372000 ;
    ANTENNADIFFAREA 1.738800 ;
    PORT
      LAYER met4 ;
        RECT 151.190 91.620 151.490 111.520 ;
    END
  END rst_n
  PIN ui_in[0]
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 147.510 110.350 147.810 111.520 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 1.304100 ;
    PORT
      LAYER met4 ;
        RECT 143.830 110.350 144.130 111.520 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 140.150 80.060 140.450 111.520 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 136.470 110.350 136.770 111.520 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 132.790 102.500 133.090 111.520 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 129.110 110.350 129.410 111.520 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 125.430 110.350 125.730 111.520 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met4 ;
        RECT 121.750 110.520 122.050 111.520 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    PORT
      LAYER met4 ;
        RECT 118.070 110.520 118.370 111.520 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    PORT
      LAYER met4 ;
        RECT 114.390 110.520 114.690 111.520 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 110.710 108.620 111.010 111.520 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 107.030 96.380 107.330 111.520 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    PORT
      LAYER met4 ;
        RECT 103.350 110.520 103.650 111.520 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    PORT
      LAYER met4 ;
        RECT 99.670 110.520 99.970 111.520 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    PORT
      LAYER met4 ;
        RECT 95.990 110.520 96.290 111.520 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    PORT
      LAYER met4 ;
        RECT 92.310 110.520 92.610 111.520 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 29.750 84.140 30.050 111.520 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 26.070 90.260 26.370 111.520 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 22.390 105.900 22.690 111.520 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 18.710 110.350 19.010 111.520 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 15.030 58.980 15.330 111.520 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 11.350 96.380 11.650 111.520 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 7.670 96.380 7.970 111.520 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 3.990 94.340 4.290 111.520 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 59.190 96.380 59.490 111.520 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 55.510 109.300 55.810 111.520 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met4 ;
        RECT 51.830 109.300 52.130 111.520 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 48.150 107.940 48.450 111.520 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met4 ;
        RECT 44.470 110.520 44.770 111.520 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 40.790 102.500 41.090 111.520 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 37.110 90.260 37.410 111.520 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 33.430 106.950 33.730 111.520 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    ANTENNAGATEAREA 0.252000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met4 ;
        RECT 88.630 90.260 88.930 111.520 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    ANTENNAGATEAREA 0.373500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met4 ;
        RECT 84.950 92.300 85.250 111.520 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    ANTENNAGATEAREA 0.252000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met4 ;
        RECT 81.270 93.660 81.570 111.520 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    ANTENNAGATEAREA 0.252000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met4 ;
        RECT 77.590 87.540 77.890 111.520 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    ANTENNAGATEAREA 0.252000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met4 ;
        RECT 73.910 91.620 74.210 111.520 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    ANTENNAGATEAREA 0.252000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met4 ;
        RECT 70.230 110.350 70.530 111.520 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    ANTENNAGATEAREA 0.252000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met4 ;
        RECT 66.550 99.470 66.850 111.520 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    ANTENNAGATEAREA 0.252000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met4 ;
        RECT 62.870 96.380 63.170 111.520 ;
    END
  END uo_out[7]
  OBS
      LAYER li1 ;
        RECT 2.760 2.635 158.240 108.885 ;
      LAYER met1 ;
        RECT 0.530 0.040 160.930 111.480 ;
      LAYER met2 ;
        RECT 0.560 0.010 160.910 111.510 ;
      LAYER met3 ;
        RECT 2.365 0.175 160.935 111.345 ;
      LAYER met4 ;
        RECT 4.690 95.980 7.270 111.345 ;
        RECT 8.370 95.980 10.950 111.345 ;
        RECT 12.050 95.980 14.630 111.345 ;
        RECT 4.690 93.940 14.630 95.980 ;
        RECT 3.975 58.580 14.630 93.940 ;
        RECT 15.730 109.950 18.310 111.345 ;
        RECT 19.410 109.950 21.990 111.345 ;
        RECT 15.730 108.100 21.990 109.950 ;
        RECT 15.730 58.580 17.880 108.100 ;
        RECT 3.975 9.600 17.880 58.580 ;
        RECT 20.280 105.500 21.990 108.100 ;
        RECT 23.090 105.500 25.670 111.345 ;
        RECT 20.280 89.860 25.670 105.500 ;
        RECT 26.770 89.860 29.350 111.345 ;
        RECT 20.280 83.740 29.350 89.860 ;
        RECT 30.450 106.550 33.030 111.345 ;
        RECT 34.130 106.550 36.710 111.345 ;
        RECT 30.450 89.860 36.710 106.550 ;
        RECT 37.810 102.100 40.390 111.345 ;
        RECT 41.490 110.120 44.070 111.345 ;
        RECT 45.170 110.120 47.750 111.345 ;
        RECT 41.490 108.100 47.750 110.120 ;
        RECT 41.490 102.100 43.480 108.100 ;
        RECT 37.810 89.860 43.480 102.100 ;
        RECT 30.450 83.740 43.480 89.860 ;
        RECT 20.280 9.600 43.480 83.740 ;
        RECT 45.880 107.540 47.750 108.100 ;
        RECT 48.850 108.900 51.430 111.345 ;
        RECT 52.530 108.900 55.110 111.345 ;
        RECT 56.210 108.900 58.790 111.345 ;
        RECT 48.850 107.540 58.790 108.900 ;
        RECT 45.880 95.980 58.790 107.540 ;
        RECT 59.890 95.980 62.470 111.345 ;
        RECT 63.570 99.070 66.150 111.345 ;
        RECT 67.250 109.950 69.830 111.345 ;
        RECT 70.930 109.950 73.510 111.345 ;
        RECT 67.250 108.100 73.510 109.950 ;
        RECT 67.250 99.070 69.080 108.100 ;
        RECT 63.570 95.980 69.080 99.070 ;
        RECT 45.880 9.600 69.080 95.980 ;
        RECT 71.480 91.220 73.510 108.100 ;
        RECT 74.610 91.220 77.190 111.345 ;
        RECT 71.480 87.140 77.190 91.220 ;
        RECT 78.290 93.260 80.870 111.345 ;
        RECT 81.970 93.260 84.550 111.345 ;
        RECT 78.290 91.900 84.550 93.260 ;
        RECT 85.650 91.900 88.230 111.345 ;
        RECT 78.290 89.860 88.230 91.900 ;
        RECT 89.330 110.120 91.910 111.345 ;
        RECT 93.010 110.120 95.590 111.345 ;
        RECT 96.690 110.120 99.270 111.345 ;
        RECT 100.370 110.120 102.950 111.345 ;
        RECT 104.050 110.120 106.630 111.345 ;
        RECT 89.330 108.100 106.630 110.120 ;
        RECT 89.330 89.860 94.680 108.100 ;
        RECT 78.290 87.140 94.680 89.860 ;
        RECT 71.480 9.600 94.680 87.140 ;
        RECT 97.080 95.980 106.630 108.100 ;
        RECT 107.730 108.220 110.310 111.345 ;
        RECT 111.410 110.120 113.990 111.345 ;
        RECT 115.090 110.120 117.670 111.345 ;
        RECT 118.770 110.120 121.350 111.345 ;
        RECT 122.450 110.120 125.030 111.345 ;
        RECT 111.410 109.950 125.030 110.120 ;
        RECT 126.130 109.950 128.710 111.345 ;
        RECT 129.810 109.950 132.390 111.345 ;
        RECT 111.410 108.220 132.390 109.950 ;
        RECT 107.730 108.100 132.390 108.220 ;
        RECT 107.730 95.980 120.280 108.100 ;
        RECT 97.080 9.600 120.280 95.980 ;
        RECT 122.680 102.100 132.390 108.100 ;
        RECT 133.490 109.950 136.070 111.345 ;
        RECT 137.170 109.950 139.750 111.345 ;
        RECT 133.490 102.100 139.750 109.950 ;
        RECT 122.680 79.660 139.750 102.100 ;
        RECT 140.850 109.950 143.430 111.345 ;
        RECT 144.530 109.950 147.110 111.345 ;
        RECT 148.210 109.950 150.790 111.345 ;
        RECT 140.850 109.440 150.790 109.950 ;
        RECT 140.850 108.100 145.880 109.440 ;
        RECT 140.850 79.660 142.780 108.100 ;
        RECT 122.680 9.600 142.780 79.660 ;
        RECT 145.180 9.600 145.880 108.100 ;
        RECT 3.975 2.080 145.880 9.600 ;
        RECT 148.280 91.220 150.790 109.440 ;
        RECT 151.890 91.220 154.470 111.345 ;
        RECT 148.280 90.540 154.470 91.220 ;
        RECT 155.570 110.120 158.150 111.345 ;
        RECT 159.250 110.120 160.705 111.345 ;
        RECT 155.570 90.540 160.705 110.120 ;
        RECT 148.280 2.080 160.705 90.540 ;
        RECT 3.975 0.855 160.705 2.080 ;
  END
END tt_um_obriensp_be8
END LIBRARY

