VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_mattvenn_inverter
  CLASS BLOCK ;
  FOREIGN tt_um_mattvenn_inverter ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 154.870 224.760 155.170 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 158.550 224.760 158.850 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 151.190 224.760 151.490 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.180000 ;
    PORT
      LAYER met4 ;
        RECT 156.560 0.000 157.160 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.300000 ;
    PORT
      LAYER met4 ;
        RECT 134.480 0.000 135.080 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 112.400 0.000 113.000 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 90.320 0.000 90.920 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 68.240 0.000 68.840 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 46.160 0.000 46.760 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 24.080 0.000 24.680 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 2.000 0.000 2.600 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 147.510 224.760 147.810 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 140.150 224.760 140.450 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 136.470 224.760 136.770 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 129.110 224.760 129.410 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 125.430 224.760 125.730 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.070 224.760 118.370 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 114.390 224.760 114.690 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.030 224.760 107.330 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 103.350 224.760 103.650 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 95.990 224.760 96.290 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 92.310 224.760 92.610 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 9.526400 ;
    PORT
      LAYER met4 ;
        RECT 29.750 224.760 30.050 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 9.526400 ;
    PORT
      LAYER met4 ;
        RECT 26.070 224.760 26.370 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 9.526400 ;
    PORT
      LAYER met4 ;
        RECT 22.390 224.760 22.690 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 9.526400 ;
    PORT
      LAYER met4 ;
        RECT 18.710 224.760 19.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 9.526400 ;
    PORT
      LAYER met4 ;
        RECT 15.030 224.760 15.330 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 9.526400 ;
    PORT
      LAYER met4 ;
        RECT 11.350 224.760 11.650 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 9.526400 ;
    PORT
      LAYER met4 ;
        RECT 7.670 224.760 7.970 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 9.526400 ;
    PORT
      LAYER met4 ;
        RECT 3.990 224.760 4.290 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 9.526400 ;
    PORT
      LAYER met4 ;
        RECT 59.190 224.760 59.490 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 9.526400 ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 9.526400 ;
    PORT
      LAYER met4 ;
        RECT 51.830 224.760 52.130 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 9.526400 ;
    PORT
      LAYER met4 ;
        RECT 48.150 224.760 48.450 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 9.526400 ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 9.526400 ;
    PORT
      LAYER met4 ;
        RECT 40.790 224.760 41.090 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 9.526400 ;
    PORT
      LAYER met4 ;
        RECT 37.110 224.760 37.410 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 9.526400 ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 9.526400 ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 9.526400 ;
    PORT
      LAYER met4 ;
        RECT 84.950 224.760 85.250 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 9.526400 ;
    PORT
      LAYER met4 ;
        RECT 81.270 224.760 81.570 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 9.526400 ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 9.526400 ;
    PORT
      LAYER met4 ;
        RECT 73.910 224.760 74.210 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 9.526400 ;
    PORT
      LAYER met4 ;
        RECT 70.230 224.760 70.530 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 9.526400 ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 9.526400 ;
    PORT
      LAYER met4 ;
        RECT 62.870 224.760 63.170 225.760 ;
    END
  END uo_out[7]
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 2.500 220.760 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 49.000 5.000 50.500 220.760 ;
    END
  END VGND
  OBS
      LAYER nwell ;
        RECT 138.250 18.030 140.360 21.220 ;
        RECT 142.520 17.980 153.790 21.170 ;
      LAYER pwell ;
        RECT 138.230 14.030 140.340 17.130 ;
        RECT 142.490 13.990 153.760 17.090 ;
      LAYER li1 ;
        RECT 138.990 21.040 139.590 21.080 ;
        RECT 138.430 20.870 140.180 21.040 ;
        RECT 144.910 20.990 150.680 21.030 ;
        RECT 138.430 18.380 138.600 20.870 ;
        RECT 138.990 20.860 139.590 20.870 ;
        RECT 139.140 20.360 139.470 20.530 ;
        RECT 139.000 19.105 139.170 20.145 ;
        RECT 139.440 19.105 139.610 20.145 ;
        RECT 139.140 18.720 139.470 18.890 ;
        RECT 140.010 18.380 140.180 20.870 ;
        RECT 138.430 18.210 140.180 18.380 ;
        RECT 142.700 20.820 153.610 20.990 ;
        RECT 142.700 18.330 142.870 20.820 ;
        RECT 144.910 20.790 150.680 20.820 ;
        RECT 143.910 20.310 144.240 20.480 ;
        RECT 144.870 20.310 145.200 20.480 ;
        RECT 145.830 20.310 146.160 20.480 ;
        RECT 146.790 20.310 147.120 20.480 ;
        RECT 147.750 20.310 148.080 20.480 ;
        RECT 148.710 20.310 149.040 20.480 ;
        RECT 149.670 20.310 150.000 20.480 ;
        RECT 150.630 20.310 150.960 20.480 ;
        RECT 151.590 20.310 151.920 20.480 ;
        RECT 152.550 20.310 152.880 20.480 ;
        RECT 143.270 19.055 143.440 20.095 ;
        RECT 143.750 19.055 143.920 20.095 ;
        RECT 144.230 19.055 144.400 20.095 ;
        RECT 144.710 19.055 144.880 20.095 ;
        RECT 145.190 19.055 145.360 20.095 ;
        RECT 145.670 19.055 145.840 20.095 ;
        RECT 146.150 19.055 146.320 20.095 ;
        RECT 146.630 19.055 146.800 20.095 ;
        RECT 147.110 19.055 147.280 20.095 ;
        RECT 147.590 19.055 147.760 20.095 ;
        RECT 148.070 19.055 148.240 20.095 ;
        RECT 148.550 19.055 148.720 20.095 ;
        RECT 149.030 19.055 149.200 20.095 ;
        RECT 149.510 19.055 149.680 20.095 ;
        RECT 149.990 19.055 150.160 20.095 ;
        RECT 150.470 19.055 150.640 20.095 ;
        RECT 150.950 19.055 151.120 20.095 ;
        RECT 151.430 19.055 151.600 20.095 ;
        RECT 151.910 19.055 152.080 20.095 ;
        RECT 152.390 19.055 152.560 20.095 ;
        RECT 152.870 19.055 153.040 20.095 ;
        RECT 143.430 18.670 143.760 18.840 ;
        RECT 144.390 18.670 144.720 18.840 ;
        RECT 145.350 18.670 145.680 18.840 ;
        RECT 146.310 18.670 146.640 18.840 ;
        RECT 147.270 18.670 147.600 18.840 ;
        RECT 148.230 18.670 148.560 18.840 ;
        RECT 149.190 18.670 149.520 18.840 ;
        RECT 150.150 18.670 150.480 18.840 ;
        RECT 151.110 18.670 151.440 18.840 ;
        RECT 152.070 18.670 152.400 18.840 ;
        RECT 153.440 18.330 153.610 20.820 ;
        RECT 142.700 18.160 153.610 18.330 ;
        RECT 138.410 16.780 140.160 16.950 ;
        RECT 138.410 14.380 138.580 16.780 ;
        RECT 139.120 16.270 139.450 16.440 ;
        RECT 138.980 15.060 139.150 16.100 ;
        RECT 139.420 15.060 139.590 16.100 ;
        RECT 139.120 14.720 139.450 14.890 ;
        RECT 139.020 14.380 139.570 14.400 ;
        RECT 139.990 14.380 140.160 16.780 ;
        RECT 138.410 14.210 140.160 14.380 ;
        RECT 142.670 16.740 153.580 16.910 ;
        RECT 142.670 14.340 142.840 16.740 ;
        RECT 143.880 16.230 144.210 16.400 ;
        RECT 144.840 16.230 145.170 16.400 ;
        RECT 145.800 16.230 146.130 16.400 ;
        RECT 146.760 16.230 147.090 16.400 ;
        RECT 147.720 16.230 148.050 16.400 ;
        RECT 148.680 16.230 149.010 16.400 ;
        RECT 149.640 16.230 149.970 16.400 ;
        RECT 150.600 16.230 150.930 16.400 ;
        RECT 151.560 16.230 151.890 16.400 ;
        RECT 152.520 16.230 152.850 16.400 ;
        RECT 143.240 15.020 143.410 16.060 ;
        RECT 143.720 15.020 143.890 16.060 ;
        RECT 144.200 15.020 144.370 16.060 ;
        RECT 144.680 15.020 144.850 16.060 ;
        RECT 145.160 15.020 145.330 16.060 ;
        RECT 145.640 15.020 145.810 16.060 ;
        RECT 146.120 15.020 146.290 16.060 ;
        RECT 146.600 15.020 146.770 16.060 ;
        RECT 147.080 15.020 147.250 16.060 ;
        RECT 147.560 15.020 147.730 16.060 ;
        RECT 148.040 15.020 148.210 16.060 ;
        RECT 148.520 15.020 148.690 16.060 ;
        RECT 149.000 15.020 149.170 16.060 ;
        RECT 149.480 15.020 149.650 16.060 ;
        RECT 149.960 15.020 150.130 16.060 ;
        RECT 150.440 15.020 150.610 16.060 ;
        RECT 150.920 15.020 151.090 16.060 ;
        RECT 151.400 15.020 151.570 16.060 ;
        RECT 151.880 15.020 152.050 16.060 ;
        RECT 152.360 15.020 152.530 16.060 ;
        RECT 152.840 15.020 153.010 16.060 ;
        RECT 143.400 14.680 143.730 14.850 ;
        RECT 144.360 14.680 144.690 14.850 ;
        RECT 145.320 14.680 145.650 14.850 ;
        RECT 146.280 14.680 146.610 14.850 ;
        RECT 147.240 14.680 147.570 14.850 ;
        RECT 148.200 14.680 148.530 14.850 ;
        RECT 149.160 14.680 149.490 14.850 ;
        RECT 150.120 14.680 150.450 14.850 ;
        RECT 151.080 14.680 151.410 14.850 ;
        RECT 152.040 14.680 152.370 14.850 ;
        RECT 145.040 14.340 150.720 14.370 ;
        RECT 153.410 14.340 153.580 16.740 ;
        RECT 139.020 14.190 139.570 14.210 ;
        RECT 142.670 14.170 153.580 14.340 ;
        RECT 145.040 14.110 150.720 14.170 ;
      LAYER mcon ;
        RECT 139.220 20.360 139.390 20.530 ;
        RECT 139.000 19.185 139.170 20.065 ;
        RECT 139.440 19.185 139.610 20.065 ;
        RECT 139.220 18.720 139.390 18.890 ;
        RECT 143.990 20.310 144.160 20.480 ;
        RECT 144.950 20.310 145.120 20.480 ;
        RECT 145.910 20.310 146.080 20.480 ;
        RECT 146.870 20.310 147.040 20.480 ;
        RECT 147.830 20.310 148.000 20.480 ;
        RECT 148.790 20.310 148.960 20.480 ;
        RECT 149.750 20.310 149.920 20.480 ;
        RECT 150.710 20.310 150.880 20.480 ;
        RECT 151.670 20.310 151.840 20.480 ;
        RECT 152.630 20.310 152.800 20.480 ;
        RECT 143.270 19.135 143.440 20.015 ;
        RECT 143.750 19.135 143.920 20.015 ;
        RECT 144.230 19.135 144.400 20.015 ;
        RECT 144.710 19.135 144.880 20.015 ;
        RECT 145.190 19.135 145.360 20.015 ;
        RECT 145.670 19.135 145.840 20.015 ;
        RECT 146.150 19.135 146.320 20.015 ;
        RECT 146.630 19.135 146.800 20.015 ;
        RECT 147.110 19.135 147.280 20.015 ;
        RECT 147.590 19.135 147.760 20.015 ;
        RECT 148.070 19.135 148.240 20.015 ;
        RECT 148.550 19.135 148.720 20.015 ;
        RECT 149.030 19.135 149.200 20.015 ;
        RECT 149.510 19.135 149.680 20.015 ;
        RECT 149.990 19.135 150.160 20.015 ;
        RECT 150.470 19.135 150.640 20.015 ;
        RECT 150.950 19.135 151.120 20.015 ;
        RECT 151.430 19.135 151.600 20.015 ;
        RECT 151.910 19.135 152.080 20.015 ;
        RECT 152.390 19.135 152.560 20.015 ;
        RECT 152.870 19.135 153.040 20.015 ;
        RECT 143.510 18.670 143.680 18.840 ;
        RECT 144.470 18.670 144.640 18.840 ;
        RECT 145.430 18.670 145.600 18.840 ;
        RECT 146.390 18.670 146.560 18.840 ;
        RECT 147.350 18.670 147.520 18.840 ;
        RECT 148.310 18.670 148.480 18.840 ;
        RECT 149.270 18.670 149.440 18.840 ;
        RECT 150.230 18.670 150.400 18.840 ;
        RECT 151.190 18.670 151.360 18.840 ;
        RECT 152.150 18.670 152.320 18.840 ;
        RECT 139.200 16.270 139.370 16.440 ;
        RECT 138.980 15.140 139.150 16.020 ;
        RECT 139.420 15.140 139.590 16.020 ;
        RECT 139.200 14.720 139.370 14.890 ;
        RECT 143.960 16.230 144.130 16.400 ;
        RECT 144.920 16.230 145.090 16.400 ;
        RECT 145.880 16.230 146.050 16.400 ;
        RECT 146.840 16.230 147.010 16.400 ;
        RECT 147.800 16.230 147.970 16.400 ;
        RECT 148.760 16.230 148.930 16.400 ;
        RECT 149.720 16.230 149.890 16.400 ;
        RECT 150.680 16.230 150.850 16.400 ;
        RECT 151.640 16.230 151.810 16.400 ;
        RECT 152.600 16.230 152.770 16.400 ;
        RECT 143.240 15.100 143.410 15.980 ;
        RECT 143.720 15.100 143.890 15.980 ;
        RECT 144.200 15.100 144.370 15.980 ;
        RECT 144.680 15.100 144.850 15.980 ;
        RECT 145.160 15.100 145.330 15.980 ;
        RECT 145.640 15.100 145.810 15.980 ;
        RECT 146.120 15.100 146.290 15.980 ;
        RECT 146.600 15.100 146.770 15.980 ;
        RECT 147.080 15.100 147.250 15.980 ;
        RECT 147.560 15.100 147.730 15.980 ;
        RECT 148.040 15.100 148.210 15.980 ;
        RECT 148.520 15.100 148.690 15.980 ;
        RECT 149.000 15.100 149.170 15.980 ;
        RECT 149.480 15.100 149.650 15.980 ;
        RECT 149.960 15.100 150.130 15.980 ;
        RECT 150.440 15.100 150.610 15.980 ;
        RECT 150.920 15.100 151.090 15.980 ;
        RECT 151.400 15.100 151.570 15.980 ;
        RECT 151.880 15.100 152.050 15.980 ;
        RECT 152.360 15.100 152.530 15.980 ;
        RECT 152.840 15.100 153.010 15.980 ;
        RECT 143.480 14.680 143.650 14.850 ;
        RECT 144.440 14.680 144.610 14.850 ;
        RECT 145.400 14.680 145.570 14.850 ;
        RECT 146.360 14.680 146.530 14.850 ;
        RECT 147.320 14.680 147.490 14.850 ;
        RECT 148.280 14.680 148.450 14.850 ;
        RECT 149.240 14.680 149.410 14.850 ;
        RECT 150.200 14.680 150.370 14.850 ;
        RECT 151.160 14.680 151.330 14.850 ;
        RECT 152.120 14.680 152.290 14.850 ;
      LAYER met1 ;
        RECT 126.950 23.280 128.450 23.310 ;
        RECT 133.190 23.280 156.260 23.380 ;
        RECT 126.950 21.880 156.260 23.280 ;
        RECT 126.950 21.780 134.410 21.880 ;
        RECT 126.950 21.750 128.450 21.780 ;
        RECT 137.540 20.030 138.030 21.880 ;
        RECT 138.870 20.770 139.700 21.880 ;
        RECT 141.870 21.620 142.230 21.880 ;
        RECT 141.840 21.260 142.260 21.620 ;
        RECT 144.830 21.310 150.830 21.880 ;
        RECT 144.820 20.760 150.830 21.310 ;
        RECT 140.425 20.590 141.670 20.595 ;
        RECT 139.110 20.345 141.670 20.590 ;
        RECT 139.110 20.340 140.680 20.345 ;
        RECT 139.160 20.330 139.450 20.340 ;
        RECT 138.970 20.030 139.200 20.125 ;
        RECT 137.540 19.320 139.200 20.030 ;
        RECT 137.970 19.260 139.200 19.320 ;
        RECT 138.970 19.125 139.200 19.260 ;
        RECT 139.410 19.890 139.640 20.125 ;
        RECT 139.410 19.490 141.130 19.890 ;
        RECT 139.410 19.125 139.640 19.490 ;
        RECT 141.425 18.945 141.670 20.345 ;
        RECT 139.125 18.695 141.670 18.945 ;
        RECT 142.140 20.315 153.115 20.565 ;
        RECT 142.140 18.885 142.390 20.315 ;
        RECT 143.930 20.280 144.220 20.315 ;
        RECT 144.890 20.280 145.180 20.315 ;
        RECT 145.850 20.280 146.140 20.315 ;
        RECT 146.810 20.280 147.100 20.315 ;
        RECT 147.770 20.280 148.060 20.315 ;
        RECT 148.730 20.280 149.020 20.315 ;
        RECT 149.690 20.280 149.980 20.315 ;
        RECT 150.650 20.280 150.940 20.315 ;
        RECT 151.610 20.280 151.900 20.315 ;
        RECT 152.570 20.280 152.860 20.315 ;
        RECT 143.240 20.040 143.470 20.075 ;
        RECT 143.180 19.750 143.560 20.040 ;
        RECT 143.240 19.075 143.470 19.750 ;
        RECT 143.720 19.410 143.950 20.075 ;
        RECT 144.200 20.060 144.430 20.075 ;
        RECT 144.140 19.770 144.520 20.060 ;
        RECT 143.660 19.140 144.020 19.410 ;
        RECT 143.720 19.075 143.950 19.140 ;
        RECT 144.200 19.075 144.430 19.770 ;
        RECT 144.680 19.430 144.910 20.075 ;
        RECT 145.160 20.070 145.390 20.075 ;
        RECT 145.070 19.760 145.440 20.070 ;
        RECT 144.620 19.160 144.980 19.430 ;
        RECT 144.680 19.075 144.910 19.160 ;
        RECT 145.160 19.075 145.390 19.760 ;
        RECT 145.640 19.410 145.870 20.075 ;
        RECT 146.120 20.050 146.350 20.075 ;
        RECT 146.080 19.740 146.450 20.050 ;
        RECT 145.570 19.140 145.930 19.410 ;
        RECT 145.640 19.075 145.870 19.140 ;
        RECT 146.120 19.075 146.350 19.740 ;
        RECT 146.600 19.390 146.830 20.075 ;
        RECT 147.080 20.050 147.310 20.075 ;
        RECT 147.020 19.740 147.390 20.050 ;
        RECT 146.510 19.120 146.870 19.390 ;
        RECT 146.600 19.075 146.830 19.120 ;
        RECT 147.080 19.075 147.310 19.740 ;
        RECT 147.560 19.420 147.790 20.075 ;
        RECT 148.040 20.070 148.270 20.075 ;
        RECT 148.000 19.760 148.370 20.070 ;
        RECT 147.490 19.150 147.850 19.420 ;
        RECT 147.560 19.075 147.790 19.150 ;
        RECT 148.040 19.075 148.270 19.760 ;
        RECT 148.520 19.400 148.750 20.075 ;
        RECT 148.920 19.770 149.290 20.080 ;
        RECT 148.460 19.130 148.820 19.400 ;
        RECT 148.520 19.075 148.750 19.130 ;
        RECT 149.000 19.075 149.230 19.770 ;
        RECT 149.480 19.380 149.710 20.075 ;
        RECT 149.960 20.030 150.190 20.075 ;
        RECT 149.900 19.720 150.270 20.030 ;
        RECT 149.420 19.110 149.780 19.380 ;
        RECT 149.480 19.075 149.710 19.110 ;
        RECT 149.960 19.075 150.190 19.720 ;
        RECT 150.440 19.400 150.670 20.075 ;
        RECT 150.920 20.050 151.150 20.075 ;
        RECT 150.860 19.740 151.230 20.050 ;
        RECT 150.400 19.130 150.760 19.400 ;
        RECT 150.440 19.075 150.670 19.130 ;
        RECT 150.920 19.075 151.150 19.740 ;
        RECT 151.400 19.400 151.630 20.075 ;
        RECT 151.820 19.770 152.190 20.080 ;
        RECT 151.360 19.130 151.720 19.400 ;
        RECT 151.400 19.075 151.630 19.130 ;
        RECT 151.880 19.075 152.110 19.770 ;
        RECT 152.360 19.400 152.590 20.075 ;
        RECT 152.780 19.770 153.150 20.080 ;
        RECT 152.280 19.130 152.640 19.400 ;
        RECT 152.360 19.075 152.590 19.130 ;
        RECT 152.840 19.075 153.070 19.770 ;
        RECT 142.085 18.805 142.390 18.885 ;
        RECT 143.450 18.805 143.740 18.870 ;
        RECT 144.410 18.805 144.700 18.870 ;
        RECT 145.370 18.805 145.660 18.870 ;
        RECT 146.330 18.805 146.620 18.870 ;
        RECT 147.290 18.805 147.580 18.870 ;
        RECT 148.250 18.805 148.540 18.870 ;
        RECT 149.210 18.805 149.500 18.870 ;
        RECT 150.170 18.805 150.460 18.870 ;
        RECT 151.130 18.805 151.420 18.870 ;
        RECT 152.090 18.805 152.380 18.870 ;
        RECT 139.160 18.690 139.450 18.695 ;
        RECT 134.750 17.745 135.750 18.000 ;
        RECT 141.105 17.745 141.355 18.695 ;
        RECT 142.085 18.555 152.685 18.805 ;
        RECT 142.085 17.820 142.335 18.555 ;
        RECT 155.080 17.950 156.080 18.240 ;
        RECT 154.240 17.830 156.080 17.950 ;
        RECT 134.750 17.740 141.355 17.745 ;
        RECT 134.480 17.495 141.355 17.740 ;
        RECT 134.480 17.030 135.750 17.495 ;
        RECT 134.450 17.000 135.750 17.030 ;
        RECT 134.450 16.430 135.110 17.000 ;
        RECT 139.130 16.460 139.800 16.490 ;
        RECT 141.105 16.460 141.355 17.495 ;
        RECT 142.080 17.360 142.480 17.820 ;
        RECT 154.240 17.420 157.190 17.830 ;
        RECT 142.085 16.460 142.335 17.360 ;
        RECT 155.080 17.240 157.190 17.420 ;
        RECT 155.210 17.230 157.190 17.240 ;
        RECT 139.130 16.270 141.730 16.460 ;
        RECT 139.140 16.240 139.430 16.270 ;
        RECT 139.580 16.230 141.730 16.270 ;
        RECT 140.600 16.210 141.730 16.230 ;
        RECT 142.085 16.220 153.155 16.460 ;
        RECT 142.085 16.210 150.910 16.220 ;
        RECT 151.200 16.210 153.155 16.220 ;
        RECT 138.950 16.030 139.180 16.080 ;
        RECT 137.880 15.930 139.180 16.030 ;
        RECT 137.540 15.260 139.180 15.930 ;
        RECT 130.820 13.560 132.320 13.590 ;
        RECT 130.820 13.400 134.960 13.560 ;
        RECT 137.540 13.400 138.000 15.260 ;
        RECT 138.950 15.080 139.180 15.260 ;
        RECT 139.390 15.780 139.620 16.080 ;
        RECT 139.390 15.380 141.130 15.780 ;
        RECT 139.390 15.080 139.620 15.380 ;
        RECT 139.140 14.895 139.430 14.920 ;
        RECT 141.475 14.895 141.725 16.210 ;
        RECT 142.085 14.895 142.335 16.210 ;
        RECT 143.900 16.200 144.190 16.210 ;
        RECT 144.860 16.200 145.150 16.210 ;
        RECT 145.820 16.200 146.110 16.210 ;
        RECT 146.780 16.200 147.070 16.210 ;
        RECT 147.740 16.200 148.030 16.210 ;
        RECT 148.700 16.200 148.990 16.210 ;
        RECT 149.660 16.200 149.950 16.210 ;
        RECT 150.620 16.200 150.910 16.210 ;
        RECT 151.580 16.200 151.870 16.210 ;
        RECT 152.540 16.200 152.830 16.210 ;
        RECT 143.210 16.010 143.440 16.040 ;
        RECT 143.150 15.720 143.530 16.010 ;
        RECT 143.210 15.040 143.440 15.720 ;
        RECT 143.690 15.380 143.920 16.040 ;
        RECT 144.170 16.030 144.400 16.040 ;
        RECT 144.110 15.740 144.490 16.030 ;
        RECT 143.630 15.110 143.990 15.380 ;
        RECT 143.690 15.040 143.920 15.110 ;
        RECT 144.170 15.040 144.400 15.740 ;
        RECT 144.650 15.400 144.880 16.040 ;
        RECT 145.040 15.730 145.410 16.040 ;
        RECT 144.590 15.130 144.950 15.400 ;
        RECT 144.650 15.040 144.880 15.130 ;
        RECT 145.130 15.040 145.360 15.730 ;
        RECT 145.610 15.380 145.840 16.040 ;
        RECT 146.090 16.020 146.320 16.040 ;
        RECT 146.050 15.710 146.420 16.020 ;
        RECT 145.540 15.110 145.900 15.380 ;
        RECT 145.610 15.040 145.840 15.110 ;
        RECT 146.090 15.040 146.320 15.710 ;
        RECT 146.570 15.360 146.800 16.040 ;
        RECT 147.050 16.020 147.280 16.040 ;
        RECT 146.990 15.710 147.360 16.020 ;
        RECT 146.480 15.090 146.840 15.360 ;
        RECT 146.570 15.040 146.800 15.090 ;
        RECT 147.050 15.040 147.280 15.710 ;
        RECT 147.530 15.390 147.760 16.040 ;
        RECT 147.970 15.730 148.340 16.040 ;
        RECT 147.460 15.120 147.820 15.390 ;
        RECT 147.530 15.040 147.760 15.120 ;
        RECT 148.010 15.040 148.240 15.730 ;
        RECT 148.490 15.370 148.720 16.040 ;
        RECT 148.890 15.740 149.260 16.050 ;
        RECT 148.430 15.100 148.790 15.370 ;
        RECT 148.490 15.040 148.720 15.100 ;
        RECT 148.970 15.040 149.200 15.740 ;
        RECT 149.450 15.350 149.680 16.040 ;
        RECT 149.930 16.000 150.160 16.040 ;
        RECT 149.870 15.690 150.240 16.000 ;
        RECT 149.390 15.080 149.750 15.350 ;
        RECT 149.450 15.040 149.680 15.080 ;
        RECT 149.930 15.040 150.160 15.690 ;
        RECT 150.410 15.370 150.640 16.040 ;
        RECT 150.890 16.020 151.120 16.040 ;
        RECT 150.830 15.710 151.200 16.020 ;
        RECT 150.370 15.100 150.730 15.370 ;
        RECT 150.410 15.040 150.640 15.100 ;
        RECT 150.890 15.040 151.120 15.710 ;
        RECT 151.370 15.370 151.600 16.040 ;
        RECT 151.790 15.740 152.160 16.050 ;
        RECT 151.330 15.100 151.690 15.370 ;
        RECT 151.370 15.040 151.600 15.100 ;
        RECT 151.850 15.040 152.080 15.740 ;
        RECT 152.330 15.370 152.560 16.040 ;
        RECT 152.750 15.740 153.120 16.050 ;
        RECT 152.250 15.100 152.610 15.370 ;
        RECT 152.330 15.040 152.560 15.100 ;
        RECT 152.810 15.040 153.040 15.740 ;
        RECT 139.105 14.645 141.730 14.895 ;
        RECT 142.085 14.655 152.755 14.895 ;
        RECT 142.240 14.645 152.755 14.655 ;
        RECT 138.910 14.370 139.670 14.440 ;
        RECT 138.900 13.400 139.670 14.370 ;
        RECT 141.820 13.840 142.240 14.200 ;
        RECT 141.850 13.400 142.210 13.840 ;
        RECT 144.830 13.400 150.830 14.400 ;
        RECT 130.820 12.060 156.610 13.400 ;
        RECT 130.820 12.030 132.320 12.060 ;
        RECT 133.540 11.900 156.610 12.060 ;
      LAYER via ;
        RECT 141.870 21.260 142.230 21.620 ;
        RECT 140.700 19.490 141.100 19.890 ;
        RECT 143.230 19.750 143.510 20.040 ;
        RECT 144.190 19.770 144.470 20.060 ;
        RECT 143.710 19.140 143.970 19.410 ;
        RECT 145.120 19.760 145.390 20.070 ;
        RECT 144.670 19.160 144.930 19.430 ;
        RECT 146.130 19.740 146.400 20.050 ;
        RECT 145.620 19.140 145.880 19.410 ;
        RECT 147.070 19.740 147.340 20.050 ;
        RECT 146.560 19.120 146.820 19.390 ;
        RECT 148.050 19.760 148.320 20.070 ;
        RECT 147.540 19.150 147.800 19.420 ;
        RECT 148.970 19.770 149.240 20.080 ;
        RECT 148.510 19.130 148.770 19.400 ;
        RECT 149.950 19.720 150.220 20.030 ;
        RECT 149.470 19.110 149.730 19.380 ;
        RECT 150.910 19.740 151.180 20.050 ;
        RECT 150.450 19.130 150.710 19.400 ;
        RECT 151.870 19.770 152.140 20.080 ;
        RECT 151.410 19.130 151.670 19.400 ;
        RECT 152.830 19.770 153.100 20.080 ;
        RECT 152.330 19.130 152.590 19.400 ;
        RECT 134.480 16.430 135.080 17.030 ;
        RECT 142.080 17.390 142.480 17.790 ;
        RECT 154.450 17.540 154.710 17.800 ;
        RECT 156.560 17.230 157.160 17.830 ;
        RECT 140.700 15.380 141.100 15.780 ;
        RECT 143.200 15.720 143.480 16.010 ;
        RECT 144.160 15.740 144.440 16.030 ;
        RECT 143.680 15.110 143.940 15.380 ;
        RECT 145.090 15.730 145.360 16.040 ;
        RECT 144.640 15.130 144.900 15.400 ;
        RECT 146.100 15.710 146.370 16.020 ;
        RECT 145.590 15.110 145.850 15.380 ;
        RECT 147.040 15.710 147.310 16.020 ;
        RECT 146.530 15.090 146.790 15.360 ;
        RECT 148.020 15.730 148.290 16.040 ;
        RECT 147.510 15.120 147.770 15.390 ;
        RECT 148.940 15.740 149.210 16.050 ;
        RECT 148.480 15.100 148.740 15.370 ;
        RECT 149.920 15.690 150.190 16.000 ;
        RECT 149.440 15.080 149.700 15.350 ;
        RECT 150.880 15.710 151.150 16.020 ;
        RECT 150.420 15.100 150.680 15.370 ;
        RECT 151.840 15.740 152.110 16.050 ;
        RECT 151.380 15.100 151.640 15.370 ;
        RECT 152.800 15.740 153.070 16.050 ;
        RECT 152.300 15.100 152.560 15.370 ;
        RECT 141.850 13.840 142.210 14.200 ;
      LAYER met2 ;
        RECT 121.765 23.280 123.215 23.300 ;
        RECT 121.740 21.780 128.480 23.280 ;
        RECT 121.765 21.760 123.215 21.780 ;
        RECT 140.700 17.790 141.100 19.920 ;
        RECT 141.870 19.460 142.230 21.650 ;
        RECT 143.230 20.040 143.510 20.090 ;
        RECT 144.190 20.040 144.470 20.110 ;
        RECT 145.120 20.040 145.390 20.120 ;
        RECT 146.130 20.040 146.400 20.100 ;
        RECT 147.070 20.040 147.340 20.100 ;
        RECT 148.050 20.040 148.320 20.120 ;
        RECT 148.970 20.040 149.240 20.130 ;
        RECT 149.950 20.040 150.220 20.080 ;
        RECT 150.910 20.040 151.180 20.100 ;
        RECT 151.870 20.040 152.140 20.130 ;
        RECT 152.830 20.040 153.100 20.130 ;
        RECT 143.180 19.780 154.710 20.040 ;
        RECT 143.230 19.700 143.510 19.780 ;
        RECT 144.190 19.720 144.470 19.780 ;
        RECT 145.120 19.710 145.390 19.780 ;
        RECT 146.130 19.690 146.400 19.780 ;
        RECT 147.070 19.690 147.340 19.780 ;
        RECT 148.050 19.710 148.320 19.780 ;
        RECT 148.970 19.720 149.240 19.780 ;
        RECT 149.950 19.670 150.220 19.780 ;
        RECT 150.910 19.690 151.180 19.780 ;
        RECT 151.870 19.720 152.140 19.780 ;
        RECT 152.830 19.720 153.100 19.780 ;
        RECT 144.670 19.460 144.930 19.480 ;
        RECT 147.540 19.460 147.800 19.470 ;
        RECT 141.870 19.100 153.850 19.460 ;
        RECT 143.710 19.090 143.970 19.100 ;
        RECT 145.620 19.090 145.880 19.100 ;
        RECT 146.560 19.070 146.820 19.100 ;
        RECT 148.510 19.080 148.770 19.100 ;
        RECT 149.470 19.060 149.730 19.100 ;
        RECT 150.450 19.080 150.710 19.100 ;
        RECT 151.410 19.080 151.670 19.100 ;
        RECT 152.330 19.080 152.590 19.100 ;
        RECT 154.450 18.140 154.710 19.780 ;
        RECT 140.700 17.390 142.510 17.790 ;
        RECT 134.480 16.215 135.080 17.060 ;
        RECT 134.460 15.665 135.100 16.215 ;
        RECT 134.480 15.640 135.080 15.665 ;
        RECT 140.700 15.350 141.100 17.390 ;
        RECT 154.340 17.175 154.810 18.140 ;
        RECT 154.340 17.040 154.965 17.175 ;
        RECT 154.450 16.590 154.965 17.040 ;
        RECT 143.200 16.010 143.480 16.060 ;
        RECT 144.160 16.010 144.440 16.080 ;
        RECT 145.090 16.010 145.360 16.090 ;
        RECT 146.100 16.010 146.370 16.070 ;
        RECT 147.040 16.010 147.310 16.070 ;
        RECT 148.020 16.010 148.290 16.090 ;
        RECT 148.940 16.010 149.210 16.100 ;
        RECT 149.920 16.010 150.190 16.050 ;
        RECT 150.880 16.010 151.150 16.070 ;
        RECT 151.840 16.010 152.110 16.100 ;
        RECT 152.800 16.010 153.070 16.100 ;
        RECT 154.400 16.010 154.965 16.590 ;
        RECT 156.560 16.585 157.160 17.860 ;
        RECT 156.540 16.035 157.180 16.585 ;
        RECT 156.560 16.010 157.160 16.035 ;
        RECT 143.150 15.750 154.965 16.010 ;
        RECT 143.200 15.670 143.480 15.750 ;
        RECT 144.160 15.690 144.440 15.750 ;
        RECT 145.090 15.680 145.360 15.750 ;
        RECT 146.100 15.660 146.370 15.750 ;
        RECT 147.040 15.660 147.310 15.750 ;
        RECT 148.020 15.680 148.290 15.750 ;
        RECT 148.940 15.690 149.210 15.750 ;
        RECT 149.920 15.640 150.190 15.750 ;
        RECT 150.880 15.660 151.150 15.750 ;
        RECT 151.840 15.690 152.110 15.750 ;
        RECT 152.800 15.690 153.070 15.750 ;
        RECT 154.400 15.555 154.965 15.750 ;
        RECT 154.400 15.530 154.660 15.555 ;
        RECT 144.640 15.430 144.900 15.450 ;
        RECT 147.510 15.430 147.770 15.440 ;
        RECT 141.850 15.070 153.820 15.430 ;
        RECT 141.850 13.810 142.210 15.070 ;
        RECT 143.680 15.060 143.940 15.070 ;
        RECT 145.590 15.060 145.850 15.070 ;
        RECT 146.530 15.040 146.790 15.070 ;
        RECT 148.480 15.050 148.740 15.070 ;
        RECT 149.440 15.030 149.700 15.070 ;
        RECT 150.420 15.050 150.680 15.070 ;
        RECT 151.380 15.050 151.640 15.070 ;
        RECT 152.300 15.050 152.560 15.070 ;
        RECT 129.755 13.560 131.205 13.580 ;
        RECT 129.730 12.060 132.350 13.560 ;
        RECT 129.755 12.040 131.205 12.060 ;
      LAYER via2 ;
        RECT 121.765 21.805 123.215 23.255 ;
        RECT 134.505 15.665 135.055 16.215 ;
        RECT 156.585 16.035 157.135 16.585 ;
        RECT 129.755 12.085 131.205 13.535 ;
      LAYER met3 ;
        RECT 34.055 23.280 35.545 23.305 ;
        RECT 34.050 21.780 123.240 23.280 ;
        RECT 34.055 21.755 35.545 21.780 ;
        RECT 134.480 15.105 135.080 16.240 ;
        RECT 134.455 14.515 135.105 15.105 ;
        RECT 156.560 14.890 157.160 16.610 ;
        RECT 156.565 14.865 157.155 14.890 ;
        RECT 134.480 14.510 135.080 14.515 ;
        RECT 128.595 13.560 130.085 13.585 ;
        RECT 128.590 12.060 131.230 13.560 ;
        RECT 128.595 12.035 130.085 12.060 ;
      LAYER via3 ;
        RECT 34.055 21.785 35.545 23.275 ;
        RECT 134.485 14.515 135.075 15.105 ;
        RECT 156.565 14.895 157.155 15.485 ;
        RECT 128.595 12.065 130.085 13.555 ;
      LAYER met4 ;
        RECT 3.990 223.380 4.290 224.760 ;
        RECT 7.670 223.380 7.970 224.760 ;
        RECT 11.350 223.380 11.650 224.760 ;
        RECT 15.030 223.380 15.330 224.760 ;
        RECT 18.710 223.380 19.010 224.760 ;
        RECT 22.390 223.380 22.690 224.760 ;
        RECT 26.070 223.380 26.370 224.760 ;
        RECT 29.750 223.380 30.050 224.760 ;
        RECT 33.430 223.380 33.730 224.760 ;
        RECT 37.110 223.380 37.410 224.760 ;
        RECT 40.790 223.380 41.090 224.760 ;
        RECT 44.470 223.380 44.770 224.760 ;
        RECT 48.150 223.380 48.450 224.760 ;
        RECT 51.830 223.380 52.130 224.760 ;
        RECT 55.510 223.380 55.810 224.760 ;
        RECT 59.190 223.380 59.490 224.760 ;
        RECT 62.870 223.380 63.170 224.760 ;
        RECT 66.550 223.380 66.850 224.760 ;
        RECT 70.230 223.380 70.530 224.760 ;
        RECT 73.910 223.380 74.210 224.760 ;
        RECT 77.590 223.380 77.890 224.760 ;
        RECT 81.270 223.380 81.570 224.760 ;
        RECT 84.950 223.380 85.250 224.760 ;
        RECT 88.630 223.380 88.930 224.760 ;
        RECT 3.400 222.070 89.640 223.380 ;
        RECT 49.000 220.760 50.500 222.070 ;
        RECT 2.500 21.780 35.550 23.280 ;
        RECT 50.500 12.060 130.090 13.560 ;
        RECT 134.480 1.000 135.080 15.110 ;
        RECT 156.560 1.000 157.160 15.490 ;
  END
END tt_um_mattvenn_inverter
END LIBRARY

