MACRO tt_um_alfiero88_VCII
  CLASS BLOCK ;
  FOREIGN tt_um_alfiero88_VCII ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 154.870 224.760 155.170 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 158.550 224.760 158.850 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 151.190 224.760 151.490 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 7.500000 ;
    ANTENNADIFFAREA 52.199997 ;
    PORT
      LAYER met4 ;
        RECT 156.560 0.000 157.160 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 15.809999 ;
    PORT
      LAYER met4 ;
        RECT 134.480 0.000 135.080 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 15.000000 ;
    ANTENNADIFFAREA 7.830000 ;
    PORT
      LAYER met4 ;
        RECT 112.400 0.000 113.000 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 15.000000 ;
    PORT
      LAYER met4 ;
        RECT 90.320 0.000 90.920 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 68.240 0.000 68.840 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 46.160 0.000 46.760 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 24.080 0.000 24.680 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 2.000 0.000 2.600 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 147.510 224.760 147.810 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 140.150 224.760 140.450 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 136.470 224.760 136.770 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 129.110 224.760 129.410 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 125.430 224.760 125.730 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.070 224.760 118.370 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 114.390 224.760 114.690 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.030 224.760 107.330 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 103.350 224.760 103.650 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 95.990 224.760 96.290 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 92.310 224.760 92.610 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 122.393394 ;
    PORT
      LAYER met4 ;
        RECT 29.750 224.760 30.050 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 122.393394 ;
    PORT
      LAYER met4 ;
        RECT 26.070 224.760 26.370 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 122.393394 ;
    PORT
      LAYER met4 ;
        RECT 22.390 224.760 22.690 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 122.393394 ;
    PORT
      LAYER met4 ;
        RECT 18.710 224.760 19.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 122.393394 ;
    PORT
      LAYER met4 ;
        RECT 15.030 224.760 15.330 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 122.393394 ;
    PORT
      LAYER met4 ;
        RECT 11.350 224.760 11.650 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 122.393394 ;
    PORT
      LAYER met4 ;
        RECT 7.670 224.760 7.970 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 122.393394 ;
    PORT
      LAYER met4 ;
        RECT 3.990 224.760 4.290 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 122.393394 ;
    PORT
      LAYER met4 ;
        RECT 59.190 224.760 59.490 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 122.393394 ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 122.393394 ;
    PORT
      LAYER met4 ;
        RECT 51.830 224.760 52.130 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 122.393394 ;
    PORT
      LAYER met4 ;
        RECT 48.150 224.760 48.450 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 122.393394 ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 122.393394 ;
    PORT
      LAYER met4 ;
        RECT 40.790 224.760 41.090 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 122.393394 ;
    PORT
      LAYER met4 ;
        RECT 37.110 224.760 37.410 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 122.393394 ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 122.393394 ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 122.393394 ;
    PORT
      LAYER met4 ;
        RECT 84.950 224.760 85.250 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 122.393394 ;
    PORT
      LAYER met4 ;
        RECT 81.270 224.760 81.570 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 122.393394 ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 122.393394 ;
    PORT
      LAYER met4 ;
        RECT 73.910 224.760 74.210 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 122.393394 ;
    PORT
      LAYER met4 ;
        RECT 70.230 224.760 70.530 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 122.393394 ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 122.393394 ;
    PORT
      LAYER met4 ;
        RECT 62.870 224.760 63.170 225.760 ;
    END
  END uo_out[7]
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 2.500 220.760 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 49.000 5.000 50.500 220.760 ;
    END
  END VGND
  OBS
      LAYER pwell ;
        RECT 107.510 117.165 110.610 141.735 ;
        RECT 112.820 117.165 115.920 141.735 ;
        RECT 121.860 136.315 135.680 142.235 ;
        RECT 121.860 134.305 137.680 136.315 ;
        RECT 121.860 130.315 137.680 134.295 ;
        RECT 107.500 89.795 110.600 114.365 ;
        RECT 125.300 112.455 136.760 127.565 ;
      LAYER nwell ;
        RECT 144.090 120.705 147.280 128.825 ;
        RECT 144.060 110.925 147.250 119.045 ;
      LAYER pwell ;
        RECT 113.230 94.615 117.330 108.085 ;
        RECT 107.510 63.475 110.610 88.045 ;
      LAYER nwell ;
        RECT 120.600 81.005 147.370 108.475 ;
      LAYER pwell ;
        RECT 107.510 37.665 110.610 62.235 ;
      LAYER nwell ;
        RECT 120.600 50.645 147.370 78.115 ;
      LAYER pwell ;
        RECT 112.620 38.285 115.720 44.535 ;
        RECT 117.660 38.245 128.850 44.715 ;
      LAYER nwell ;
        RECT 130.500 38.185 137.690 44.655 ;
        RECT 139.900 43.785 147.090 46.745 ;
        RECT 139.890 38.325 147.080 41.285 ;
      LAYER pwell ;
        RECT 109.220 36.355 109.570 37.665 ;
      LAYER li1 ;
        RECT 122.040 141.885 135.500 142.055 ;
        RECT 113.730 141.555 115.050 141.695 ;
        RECT 122.040 141.645 122.210 141.885 ;
        RECT 107.690 141.385 110.430 141.555 ;
        RECT 107.690 136.845 107.860 141.385 ;
        RECT 108.540 140.815 109.580 140.985 ;
        RECT 108.200 138.755 108.370 140.755 ;
        RECT 109.750 138.755 109.920 140.755 ;
        RECT 108.540 138.525 109.580 138.695 ;
        RECT 107.480 135.805 107.940 136.845 ;
        RECT 108.200 136.465 108.370 138.465 ;
        RECT 109.750 136.465 109.920 138.465 ;
        RECT 108.540 136.235 109.580 136.405 ;
        RECT 107.690 122.965 107.860 135.805 ;
        RECT 108.200 134.175 108.370 136.175 ;
        RECT 109.750 134.175 109.920 136.175 ;
        RECT 108.540 133.945 109.580 134.115 ;
        RECT 108.200 131.885 108.370 133.885 ;
        RECT 109.750 131.885 109.920 133.885 ;
        RECT 108.540 131.655 109.580 131.825 ;
        RECT 108.200 129.595 108.370 131.595 ;
        RECT 109.750 129.595 109.920 131.595 ;
        RECT 108.540 129.365 109.580 129.535 ;
        RECT 108.200 127.305 108.370 129.305 ;
        RECT 109.750 127.305 109.920 129.305 ;
        RECT 108.540 127.075 109.580 127.245 ;
        RECT 108.200 125.015 108.370 127.015 ;
        RECT 109.750 125.015 109.920 127.015 ;
        RECT 108.540 124.785 109.580 124.955 ;
        RECT 107.500 121.805 107.940 122.965 ;
        RECT 108.200 122.725 108.370 124.725 ;
        RECT 109.750 122.725 109.920 124.725 ;
        RECT 108.540 122.495 109.580 122.665 ;
        RECT 107.690 117.515 107.860 121.805 ;
        RECT 108.200 120.435 108.370 122.435 ;
        RECT 109.750 120.435 109.920 122.435 ;
        RECT 108.540 120.205 109.580 120.375 ;
        RECT 108.200 118.145 108.370 120.145 ;
        RECT 109.750 118.145 109.920 120.145 ;
        RECT 108.540 117.915 109.580 118.085 ;
        RECT 110.260 117.515 110.430 141.385 ;
        RECT 107.690 117.345 110.430 117.515 ;
        RECT 113.000 141.385 115.740 141.555 ;
        RECT 113.000 117.515 113.170 141.385 ;
        RECT 113.730 141.325 115.050 141.385 ;
        RECT 113.850 140.815 114.890 140.985 ;
        RECT 113.510 138.755 113.680 140.755 ;
        RECT 115.060 138.755 115.230 140.755 ;
        RECT 113.850 138.525 114.890 138.695 ;
        RECT 113.510 136.465 113.680 138.465 ;
        RECT 115.060 136.465 115.230 138.465 ;
        RECT 113.850 136.235 114.890 136.405 ;
        RECT 113.510 134.175 113.680 136.175 ;
        RECT 115.060 134.175 115.230 136.175 ;
        RECT 113.850 133.945 114.890 134.115 ;
        RECT 113.510 131.885 113.680 133.885 ;
        RECT 115.060 131.885 115.230 133.885 ;
        RECT 113.850 131.655 114.890 131.825 ;
        RECT 113.510 129.595 113.680 131.595 ;
        RECT 115.060 129.595 115.230 131.595 ;
        RECT 113.850 129.365 114.890 129.535 ;
        RECT 113.510 127.305 113.680 129.305 ;
        RECT 115.060 127.305 115.230 129.305 ;
        RECT 113.850 127.075 114.890 127.245 ;
        RECT 113.510 125.015 113.680 127.015 ;
        RECT 115.060 125.015 115.230 127.015 ;
        RECT 113.850 124.785 114.890 124.955 ;
        RECT 113.510 122.725 113.680 124.725 ;
        RECT 115.060 122.725 115.230 124.725 ;
        RECT 113.850 122.495 114.890 122.665 ;
        RECT 113.510 120.435 113.680 122.435 ;
        RECT 115.060 120.435 115.230 122.435 ;
        RECT 113.850 120.205 114.890 120.375 ;
        RECT 113.510 118.145 113.680 120.145 ;
        RECT 115.060 118.145 115.230 120.145 ;
        RECT 113.850 117.915 114.890 118.085 ;
        RECT 115.570 117.515 115.740 141.385 ;
        RECT 121.980 140.825 122.260 141.645 ;
        RECT 122.690 141.055 124.850 141.405 ;
        RECT 132.690 141.055 134.850 141.405 ;
        RECT 122.040 140.575 122.210 140.825 ;
        RECT 135.330 140.575 135.500 141.885 ;
        RECT 122.040 140.405 135.500 140.575 ;
        RECT 122.040 139.925 135.500 140.095 ;
        RECT 122.040 139.675 122.210 139.925 ;
        RECT 121.980 138.855 122.260 139.675 ;
        RECT 122.690 139.095 124.850 139.445 ;
        RECT 132.690 139.095 134.850 139.445 ;
        RECT 122.040 138.615 122.210 138.855 ;
        RECT 135.330 138.615 135.500 139.925 ;
        RECT 122.040 138.445 135.500 138.615 ;
        RECT 122.040 137.955 135.500 138.125 ;
        RECT 122.040 137.705 122.210 137.955 ;
        RECT 121.980 136.885 122.260 137.705 ;
        RECT 122.690 137.125 124.850 137.475 ;
        RECT 132.690 137.125 134.850 137.475 ;
        RECT 122.040 136.645 122.210 136.885 ;
        RECT 135.330 136.645 135.500 137.955 ;
        RECT 122.040 136.475 135.500 136.645 ;
        RECT 122.040 135.965 137.500 136.135 ;
        RECT 122.040 135.745 122.210 135.965 ;
        RECT 121.980 134.895 122.270 135.745 ;
        RECT 122.690 135.135 124.850 135.485 ;
        RECT 134.690 135.135 136.850 135.485 ;
        RECT 122.040 134.655 122.210 134.895 ;
        RECT 137.330 134.655 137.500 135.965 ;
        RECT 122.040 134.485 137.500 134.655 ;
        RECT 122.040 133.945 137.500 134.115 ;
        RECT 122.040 133.685 122.210 133.945 ;
        RECT 121.980 132.865 122.270 133.685 ;
        RECT 122.690 133.115 124.850 133.465 ;
        RECT 134.690 133.115 136.850 133.465 ;
        RECT 122.040 132.635 122.210 132.865 ;
        RECT 137.330 132.635 137.500 133.945 ;
        RECT 122.040 132.465 137.500 132.635 ;
        RECT 122.040 131.975 137.500 132.145 ;
        RECT 122.040 131.725 122.210 131.975 ;
        RECT 121.980 130.915 122.270 131.725 ;
        RECT 122.690 131.145 124.850 131.495 ;
        RECT 134.690 131.145 136.850 131.495 ;
        RECT 122.040 130.665 122.210 130.915 ;
        RECT 137.330 130.665 137.500 131.975 ;
        RECT 122.040 130.495 137.500 130.665 ;
        RECT 144.270 128.475 147.100 128.645 ;
        RECT 125.480 127.215 136.580 127.385 ;
        RECT 125.480 124.255 125.650 127.215 ;
        RECT 126.330 126.645 127.370 126.815 ;
        RECT 128.420 126.645 129.460 126.815 ;
        RECT 130.510 126.645 131.550 126.815 ;
        RECT 132.600 126.645 133.640 126.815 ;
        RECT 134.690 126.645 135.730 126.815 ;
        RECT 125.990 126.270 126.160 126.600 ;
        RECT 127.540 126.270 127.710 126.600 ;
        RECT 128.080 126.270 128.250 126.600 ;
        RECT 129.630 126.270 129.800 126.600 ;
        RECT 130.170 126.270 130.340 126.600 ;
        RECT 131.720 126.270 131.890 126.600 ;
        RECT 132.260 126.270 132.430 126.600 ;
        RECT 133.810 126.270 133.980 126.600 ;
        RECT 134.350 126.270 134.520 126.600 ;
        RECT 135.900 126.270 136.070 126.600 ;
        RECT 126.330 126.055 127.370 126.225 ;
        RECT 128.420 126.055 129.460 126.225 ;
        RECT 130.510 126.055 131.550 126.225 ;
        RECT 132.600 126.055 133.640 126.225 ;
        RECT 134.690 126.055 135.730 126.225 ;
        RECT 125.990 125.680 126.160 126.010 ;
        RECT 127.540 125.680 127.710 126.010 ;
        RECT 128.080 125.680 128.250 126.010 ;
        RECT 129.630 125.680 129.800 126.010 ;
        RECT 130.170 125.680 130.340 126.010 ;
        RECT 131.720 125.680 131.890 126.010 ;
        RECT 132.260 125.680 132.430 126.010 ;
        RECT 133.810 125.680 133.980 126.010 ;
        RECT 134.350 125.680 134.520 126.010 ;
        RECT 135.900 125.680 136.070 126.010 ;
        RECT 126.330 125.465 127.370 125.635 ;
        RECT 128.420 125.465 129.460 125.635 ;
        RECT 130.510 125.465 131.550 125.635 ;
        RECT 132.600 125.465 133.640 125.635 ;
        RECT 134.690 125.465 135.730 125.635 ;
        RECT 125.990 125.090 126.160 125.420 ;
        RECT 127.540 125.090 127.710 125.420 ;
        RECT 128.080 125.090 128.250 125.420 ;
        RECT 129.630 125.090 129.800 125.420 ;
        RECT 130.170 125.090 130.340 125.420 ;
        RECT 131.720 125.090 131.890 125.420 ;
        RECT 132.260 125.090 132.430 125.420 ;
        RECT 133.810 125.090 133.980 125.420 ;
        RECT 134.350 125.090 134.520 125.420 ;
        RECT 135.900 125.090 136.070 125.420 ;
        RECT 126.330 124.875 127.370 125.045 ;
        RECT 128.420 124.875 129.460 125.045 ;
        RECT 130.510 124.875 131.550 125.045 ;
        RECT 132.600 124.875 133.640 125.045 ;
        RECT 134.690 124.875 135.730 125.045 ;
        RECT 125.990 124.500 126.160 124.830 ;
        RECT 127.540 124.500 127.710 124.830 ;
        RECT 128.080 124.500 128.250 124.830 ;
        RECT 129.630 124.500 129.800 124.830 ;
        RECT 130.170 124.500 130.340 124.830 ;
        RECT 131.720 124.500 131.890 124.830 ;
        RECT 132.260 124.500 132.430 124.830 ;
        RECT 133.810 124.500 133.980 124.830 ;
        RECT 134.350 124.500 134.520 124.830 ;
        RECT 135.900 124.500 136.070 124.830 ;
        RECT 126.330 124.285 127.370 124.455 ;
        RECT 128.420 124.285 129.460 124.455 ;
        RECT 130.510 124.285 131.550 124.455 ;
        RECT 132.600 124.285 133.640 124.455 ;
        RECT 134.690 124.285 135.730 124.455 ;
        RECT 125.400 123.065 125.690 124.255 ;
        RECT 125.990 123.910 126.160 124.240 ;
        RECT 127.540 123.910 127.710 124.240 ;
        RECT 128.080 123.910 128.250 124.240 ;
        RECT 129.630 123.910 129.800 124.240 ;
        RECT 130.170 123.910 130.340 124.240 ;
        RECT 131.720 123.910 131.890 124.240 ;
        RECT 132.260 123.910 132.430 124.240 ;
        RECT 133.810 123.910 133.980 124.240 ;
        RECT 134.350 123.910 134.520 124.240 ;
        RECT 135.900 123.910 136.070 124.240 ;
        RECT 126.330 123.695 127.370 123.865 ;
        RECT 128.420 123.695 129.460 123.865 ;
        RECT 130.510 123.695 131.550 123.865 ;
        RECT 132.600 123.695 133.640 123.865 ;
        RECT 134.690 123.695 135.730 123.865 ;
        RECT 125.990 123.320 126.160 123.650 ;
        RECT 127.540 123.320 127.710 123.650 ;
        RECT 128.080 123.320 128.250 123.650 ;
        RECT 129.630 123.320 129.800 123.650 ;
        RECT 130.170 123.320 130.340 123.650 ;
        RECT 131.720 123.320 131.890 123.650 ;
        RECT 132.260 123.320 132.430 123.650 ;
        RECT 133.810 123.320 133.980 123.650 ;
        RECT 134.350 123.320 134.520 123.650 ;
        RECT 135.900 123.320 136.070 123.650 ;
        RECT 126.330 123.105 127.370 123.275 ;
        RECT 128.420 123.105 129.460 123.275 ;
        RECT 130.510 123.105 131.550 123.275 ;
        RECT 132.600 123.105 133.640 123.275 ;
        RECT 134.690 123.105 135.730 123.275 ;
        RECT 125.480 120.345 125.650 123.065 ;
        RECT 125.990 122.730 126.160 123.060 ;
        RECT 127.540 122.730 127.710 123.060 ;
        RECT 128.080 122.730 128.250 123.060 ;
        RECT 129.630 122.730 129.800 123.060 ;
        RECT 130.170 122.730 130.340 123.060 ;
        RECT 131.720 122.730 131.890 123.060 ;
        RECT 132.260 122.730 132.430 123.060 ;
        RECT 133.810 122.730 133.980 123.060 ;
        RECT 134.350 122.730 134.520 123.060 ;
        RECT 135.900 122.730 136.070 123.060 ;
        RECT 126.330 122.515 127.370 122.685 ;
        RECT 128.420 122.515 129.460 122.685 ;
        RECT 130.510 122.515 131.550 122.685 ;
        RECT 132.600 122.515 133.640 122.685 ;
        RECT 134.690 122.515 135.730 122.685 ;
        RECT 125.990 122.140 126.160 122.470 ;
        RECT 127.540 122.140 127.710 122.470 ;
        RECT 128.080 122.140 128.250 122.470 ;
        RECT 129.630 122.140 129.800 122.470 ;
        RECT 130.170 122.140 130.340 122.470 ;
        RECT 131.720 122.140 131.890 122.470 ;
        RECT 132.260 122.140 132.430 122.470 ;
        RECT 133.810 122.140 133.980 122.470 ;
        RECT 134.350 122.140 134.520 122.470 ;
        RECT 135.900 122.140 136.070 122.470 ;
        RECT 126.330 121.925 127.370 122.095 ;
        RECT 128.420 121.925 129.460 122.095 ;
        RECT 130.510 121.925 131.550 122.095 ;
        RECT 132.600 121.925 133.640 122.095 ;
        RECT 134.690 121.925 135.730 122.095 ;
        RECT 125.990 121.550 126.160 121.880 ;
        RECT 127.540 121.550 127.710 121.880 ;
        RECT 128.080 121.550 128.250 121.880 ;
        RECT 129.630 121.550 129.800 121.880 ;
        RECT 130.170 121.550 130.340 121.880 ;
        RECT 131.720 121.550 131.890 121.880 ;
        RECT 132.260 121.550 132.430 121.880 ;
        RECT 133.810 121.550 133.980 121.880 ;
        RECT 134.350 121.550 134.520 121.880 ;
        RECT 135.900 121.550 136.070 121.880 ;
        RECT 126.330 121.335 127.370 121.505 ;
        RECT 128.420 121.335 129.460 121.505 ;
        RECT 130.510 121.335 131.550 121.505 ;
        RECT 132.600 121.335 133.640 121.505 ;
        RECT 134.690 121.335 135.730 121.505 ;
        RECT 125.990 120.960 126.160 121.290 ;
        RECT 127.540 120.960 127.710 121.290 ;
        RECT 128.080 120.960 128.250 121.290 ;
        RECT 129.630 120.960 129.800 121.290 ;
        RECT 130.170 120.960 130.340 121.290 ;
        RECT 131.720 120.960 131.890 121.290 ;
        RECT 132.260 120.960 132.430 121.290 ;
        RECT 133.810 120.960 133.980 121.290 ;
        RECT 134.350 120.960 134.520 121.290 ;
        RECT 135.900 120.960 136.070 121.290 ;
        RECT 126.330 120.745 127.370 120.915 ;
        RECT 128.420 120.745 129.460 120.915 ;
        RECT 130.510 120.745 131.550 120.915 ;
        RECT 132.600 120.745 133.640 120.915 ;
        RECT 134.690 120.745 135.730 120.915 ;
        RECT 136.410 120.345 136.580 127.215 ;
        RECT 144.270 121.055 144.440 128.475 ;
        RECT 145.165 127.905 146.205 128.075 ;
        RECT 144.780 126.845 144.950 127.845 ;
        RECT 146.420 126.845 146.590 127.845 ;
        RECT 145.165 126.615 146.205 126.785 ;
        RECT 144.780 125.555 144.950 126.555 ;
        RECT 146.420 125.555 146.590 126.555 ;
        RECT 145.165 125.325 146.205 125.495 ;
        RECT 146.930 125.275 147.100 128.475 ;
        RECT 144.780 124.265 144.950 125.265 ;
        RECT 146.420 124.265 146.590 125.265 ;
        RECT 146.860 124.225 147.210 125.275 ;
        RECT 145.165 124.035 146.205 124.205 ;
        RECT 144.780 122.975 144.950 123.975 ;
        RECT 146.420 122.975 146.590 123.975 ;
        RECT 145.165 122.745 146.205 122.915 ;
        RECT 144.780 121.685 144.950 122.685 ;
        RECT 146.420 121.685 146.590 122.685 ;
        RECT 145.165 121.455 146.205 121.625 ;
        RECT 146.930 121.055 147.100 124.225 ;
        RECT 144.270 120.885 147.100 121.055 ;
        RECT 125.480 120.175 136.580 120.345 ;
        RECT 113.000 117.345 115.740 117.515 ;
        RECT 125.480 119.675 136.580 119.845 ;
        RECT 125.480 116.865 125.650 119.675 ;
        RECT 126.330 119.105 127.370 119.275 ;
        RECT 128.420 119.105 129.460 119.275 ;
        RECT 130.510 119.105 131.550 119.275 ;
        RECT 132.600 119.105 133.640 119.275 ;
        RECT 134.690 119.105 135.730 119.275 ;
        RECT 125.990 118.730 126.160 119.060 ;
        RECT 127.540 118.730 127.710 119.060 ;
        RECT 128.080 118.730 128.250 119.060 ;
        RECT 129.630 118.730 129.800 119.060 ;
        RECT 130.170 118.730 130.340 119.060 ;
        RECT 131.720 118.730 131.890 119.060 ;
        RECT 132.260 118.730 132.430 119.060 ;
        RECT 133.810 118.730 133.980 119.060 ;
        RECT 134.350 118.730 134.520 119.060 ;
        RECT 135.900 118.730 136.070 119.060 ;
        RECT 126.330 118.515 127.370 118.685 ;
        RECT 128.420 118.515 129.460 118.685 ;
        RECT 130.510 118.515 131.550 118.685 ;
        RECT 132.600 118.515 133.640 118.685 ;
        RECT 134.690 118.515 135.730 118.685 ;
        RECT 125.990 118.140 126.160 118.470 ;
        RECT 127.540 118.140 127.710 118.470 ;
        RECT 128.080 118.140 128.250 118.470 ;
        RECT 129.630 118.140 129.800 118.470 ;
        RECT 130.170 118.140 130.340 118.470 ;
        RECT 131.720 118.140 131.890 118.470 ;
        RECT 132.260 118.140 132.430 118.470 ;
        RECT 133.810 118.140 133.980 118.470 ;
        RECT 134.350 118.140 134.520 118.470 ;
        RECT 135.900 118.140 136.070 118.470 ;
        RECT 126.330 117.925 127.370 118.095 ;
        RECT 128.420 117.925 129.460 118.095 ;
        RECT 130.510 117.925 131.550 118.095 ;
        RECT 132.600 117.925 133.640 118.095 ;
        RECT 134.690 117.925 135.730 118.095 ;
        RECT 125.990 117.550 126.160 117.880 ;
        RECT 127.540 117.550 127.710 117.880 ;
        RECT 128.080 117.550 128.250 117.880 ;
        RECT 129.630 117.550 129.800 117.880 ;
        RECT 130.170 117.550 130.340 117.880 ;
        RECT 131.720 117.550 131.890 117.880 ;
        RECT 132.260 117.550 132.430 117.880 ;
        RECT 133.810 117.550 133.980 117.880 ;
        RECT 134.350 117.550 134.520 117.880 ;
        RECT 135.900 117.550 136.070 117.880 ;
        RECT 126.330 117.335 127.370 117.505 ;
        RECT 128.420 117.335 129.460 117.505 ;
        RECT 130.510 117.335 131.550 117.505 ;
        RECT 132.600 117.335 133.640 117.505 ;
        RECT 134.690 117.335 135.730 117.505 ;
        RECT 125.990 116.960 126.160 117.290 ;
        RECT 127.540 116.960 127.710 117.290 ;
        RECT 128.080 116.960 128.250 117.290 ;
        RECT 129.630 116.960 129.800 117.290 ;
        RECT 130.170 116.960 130.340 117.290 ;
        RECT 131.720 116.960 131.890 117.290 ;
        RECT 132.260 116.960 132.430 117.290 ;
        RECT 133.810 116.960 133.980 117.290 ;
        RECT 134.350 116.960 134.520 117.290 ;
        RECT 135.900 116.960 136.070 117.290 ;
        RECT 125.390 115.655 125.700 116.865 ;
        RECT 126.330 116.745 127.370 116.915 ;
        RECT 128.420 116.745 129.460 116.915 ;
        RECT 130.510 116.745 131.550 116.915 ;
        RECT 132.600 116.745 133.640 116.915 ;
        RECT 134.690 116.745 135.730 116.915 ;
        RECT 125.990 116.370 126.160 116.700 ;
        RECT 127.540 116.370 127.710 116.700 ;
        RECT 128.080 116.370 128.250 116.700 ;
        RECT 129.630 116.370 129.800 116.700 ;
        RECT 130.170 116.370 130.340 116.700 ;
        RECT 131.720 116.370 131.890 116.700 ;
        RECT 132.260 116.370 132.430 116.700 ;
        RECT 133.810 116.370 133.980 116.700 ;
        RECT 134.350 116.370 134.520 116.700 ;
        RECT 135.900 116.370 136.070 116.700 ;
        RECT 126.330 116.155 127.370 116.325 ;
        RECT 128.420 116.155 129.460 116.325 ;
        RECT 130.510 116.155 131.550 116.325 ;
        RECT 132.600 116.155 133.640 116.325 ;
        RECT 134.690 116.155 135.730 116.325 ;
        RECT 125.990 115.780 126.160 116.110 ;
        RECT 127.540 115.780 127.710 116.110 ;
        RECT 128.080 115.780 128.250 116.110 ;
        RECT 129.630 115.780 129.800 116.110 ;
        RECT 130.170 115.780 130.340 116.110 ;
        RECT 131.720 115.780 131.890 116.110 ;
        RECT 132.260 115.780 132.430 116.110 ;
        RECT 133.810 115.780 133.980 116.110 ;
        RECT 134.350 115.780 134.520 116.110 ;
        RECT 135.900 115.780 136.070 116.110 ;
        RECT 107.680 114.015 110.420 114.185 ;
        RECT 107.680 109.455 107.850 114.015 ;
        RECT 108.530 113.445 109.570 113.615 ;
        RECT 108.190 111.385 108.360 113.385 ;
        RECT 109.740 111.385 109.910 113.385 ;
        RECT 108.530 111.155 109.570 111.325 ;
        RECT 107.530 108.265 107.960 109.455 ;
        RECT 108.190 109.095 108.360 111.095 ;
        RECT 109.740 109.095 109.910 111.095 ;
        RECT 108.530 108.865 109.570 109.035 ;
        RECT 107.680 95.735 107.850 108.265 ;
        RECT 108.190 106.805 108.360 108.805 ;
        RECT 109.740 106.805 109.910 108.805 ;
        RECT 108.530 106.575 109.570 106.745 ;
        RECT 108.190 104.515 108.360 106.515 ;
        RECT 109.740 104.515 109.910 106.515 ;
        RECT 108.530 104.285 109.570 104.455 ;
        RECT 108.190 102.225 108.360 104.225 ;
        RECT 109.740 102.225 109.910 104.225 ;
        RECT 108.530 101.995 109.570 102.165 ;
        RECT 108.190 99.935 108.360 101.935 ;
        RECT 109.740 99.935 109.910 101.935 ;
        RECT 108.530 99.705 109.570 99.875 ;
        RECT 108.190 97.645 108.360 99.645 ;
        RECT 109.740 97.645 109.910 99.645 ;
        RECT 108.530 97.415 109.570 97.585 ;
        RECT 107.530 94.535 107.950 95.735 ;
        RECT 108.190 95.355 108.360 97.355 ;
        RECT 109.740 95.355 109.910 97.355 ;
        RECT 108.530 95.125 109.570 95.295 ;
        RECT 107.680 90.145 107.850 94.535 ;
        RECT 108.190 93.065 108.360 95.065 ;
        RECT 109.740 93.065 109.910 95.065 ;
        RECT 108.530 92.835 109.570 93.005 ;
        RECT 108.190 90.775 108.360 92.775 ;
        RECT 109.740 90.775 109.910 92.775 ;
        RECT 108.530 90.545 109.570 90.715 ;
        RECT 110.250 90.145 110.420 114.015 ;
        RECT 125.480 112.805 125.650 115.655 ;
        RECT 126.330 115.565 127.370 115.735 ;
        RECT 128.420 115.565 129.460 115.735 ;
        RECT 130.510 115.565 131.550 115.735 ;
        RECT 132.600 115.565 133.640 115.735 ;
        RECT 134.690 115.565 135.730 115.735 ;
        RECT 125.990 115.190 126.160 115.520 ;
        RECT 127.540 115.190 127.710 115.520 ;
        RECT 128.080 115.190 128.250 115.520 ;
        RECT 129.630 115.190 129.800 115.520 ;
        RECT 130.170 115.190 130.340 115.520 ;
        RECT 131.720 115.190 131.890 115.520 ;
        RECT 132.260 115.190 132.430 115.520 ;
        RECT 133.810 115.190 133.980 115.520 ;
        RECT 134.350 115.190 134.520 115.520 ;
        RECT 135.900 115.190 136.070 115.520 ;
        RECT 126.330 114.975 127.370 115.145 ;
        RECT 128.420 114.975 129.460 115.145 ;
        RECT 130.510 114.975 131.550 115.145 ;
        RECT 132.600 114.975 133.640 115.145 ;
        RECT 134.690 114.975 135.730 115.145 ;
        RECT 125.990 114.600 126.160 114.930 ;
        RECT 127.540 114.600 127.710 114.930 ;
        RECT 128.080 114.600 128.250 114.930 ;
        RECT 129.630 114.600 129.800 114.930 ;
        RECT 130.170 114.600 130.340 114.930 ;
        RECT 131.720 114.600 131.890 114.930 ;
        RECT 132.260 114.600 132.430 114.930 ;
        RECT 133.810 114.600 133.980 114.930 ;
        RECT 134.350 114.600 134.520 114.930 ;
        RECT 135.900 114.600 136.070 114.930 ;
        RECT 126.330 114.385 127.370 114.555 ;
        RECT 128.420 114.385 129.460 114.555 ;
        RECT 130.510 114.385 131.550 114.555 ;
        RECT 132.600 114.385 133.640 114.555 ;
        RECT 134.690 114.385 135.730 114.555 ;
        RECT 125.990 114.010 126.160 114.340 ;
        RECT 127.540 114.010 127.710 114.340 ;
        RECT 128.080 114.010 128.250 114.340 ;
        RECT 129.630 114.010 129.800 114.340 ;
        RECT 130.170 114.010 130.340 114.340 ;
        RECT 131.720 114.010 131.890 114.340 ;
        RECT 132.260 114.010 132.430 114.340 ;
        RECT 133.810 114.010 133.980 114.340 ;
        RECT 134.350 114.010 134.520 114.340 ;
        RECT 135.900 114.010 136.070 114.340 ;
        RECT 126.330 113.795 127.370 113.965 ;
        RECT 128.420 113.795 129.460 113.965 ;
        RECT 130.510 113.795 131.550 113.965 ;
        RECT 132.600 113.795 133.640 113.965 ;
        RECT 134.690 113.795 135.730 113.965 ;
        RECT 125.990 113.420 126.160 113.750 ;
        RECT 127.540 113.420 127.710 113.750 ;
        RECT 128.080 113.420 128.250 113.750 ;
        RECT 129.630 113.420 129.800 113.750 ;
        RECT 130.170 113.420 130.340 113.750 ;
        RECT 131.720 113.420 131.890 113.750 ;
        RECT 132.260 113.420 132.430 113.750 ;
        RECT 133.810 113.420 133.980 113.750 ;
        RECT 134.350 113.420 134.520 113.750 ;
        RECT 135.900 113.420 136.070 113.750 ;
        RECT 126.330 113.205 127.370 113.375 ;
        RECT 128.420 113.205 129.460 113.375 ;
        RECT 130.510 113.205 131.550 113.375 ;
        RECT 132.600 113.205 133.640 113.375 ;
        RECT 134.690 113.205 135.730 113.375 ;
        RECT 136.410 112.805 136.580 119.675 ;
        RECT 125.480 112.635 136.580 112.805 ;
        RECT 144.240 118.695 147.070 118.865 ;
        RECT 144.240 111.275 144.410 118.695 ;
        RECT 145.135 118.125 146.175 118.295 ;
        RECT 144.750 117.065 144.920 118.065 ;
        RECT 146.390 117.065 146.560 118.065 ;
        RECT 145.135 116.835 146.175 117.005 ;
        RECT 144.750 115.775 144.920 116.775 ;
        RECT 146.390 115.775 146.560 116.775 ;
        RECT 145.135 115.545 146.175 115.715 ;
        RECT 144.750 114.485 144.920 115.485 ;
        RECT 146.390 114.485 146.560 115.485 ;
        RECT 146.900 115.385 147.070 118.695 ;
        RECT 146.850 114.425 147.190 115.385 ;
        RECT 145.135 114.255 146.175 114.425 ;
        RECT 144.750 113.195 144.920 114.195 ;
        RECT 146.390 113.195 146.560 114.195 ;
        RECT 145.135 112.965 146.175 113.135 ;
        RECT 144.750 111.905 144.920 112.905 ;
        RECT 146.390 111.905 146.560 112.905 ;
        RECT 145.135 111.675 146.175 111.845 ;
        RECT 146.900 111.275 147.070 114.425 ;
        RECT 144.240 111.105 147.070 111.275 ;
        RECT 120.780 108.125 147.190 108.295 ;
        RECT 113.410 107.735 117.150 107.905 ;
        RECT 113.410 103.615 113.580 107.735 ;
        RECT 114.260 107.165 116.300 107.335 ;
        RECT 113.920 106.790 114.090 107.120 ;
        RECT 116.470 106.790 116.640 107.120 ;
        RECT 114.260 106.575 116.300 106.745 ;
        RECT 113.920 106.200 114.090 106.530 ;
        RECT 116.470 106.200 116.640 106.530 ;
        RECT 114.260 105.985 116.300 106.155 ;
        RECT 113.920 105.610 114.090 105.940 ;
        RECT 116.470 105.610 116.640 105.940 ;
        RECT 114.260 105.395 116.300 105.565 ;
        RECT 113.920 105.020 114.090 105.350 ;
        RECT 116.470 105.020 116.640 105.350 ;
        RECT 114.260 104.805 116.300 104.975 ;
        RECT 113.920 104.430 114.090 104.760 ;
        RECT 116.470 104.430 116.640 104.760 ;
        RECT 114.260 104.215 116.300 104.385 ;
        RECT 113.920 103.840 114.090 104.170 ;
        RECT 116.470 103.840 116.640 104.170 ;
        RECT 114.260 103.625 116.300 103.795 ;
        RECT 113.280 99.905 113.600 103.615 ;
        RECT 113.920 103.250 114.090 103.580 ;
        RECT 116.470 103.250 116.640 103.580 ;
        RECT 114.260 103.035 116.300 103.205 ;
        RECT 113.920 102.660 114.090 102.990 ;
        RECT 116.470 102.660 116.640 102.990 ;
        RECT 114.260 102.445 116.300 102.615 ;
        RECT 113.920 102.070 114.090 102.400 ;
        RECT 116.470 102.070 116.640 102.400 ;
        RECT 114.260 101.855 116.300 102.025 ;
        RECT 113.920 101.480 114.090 101.810 ;
        RECT 116.470 101.480 116.640 101.810 ;
        RECT 114.260 101.265 116.300 101.435 ;
        RECT 113.920 100.890 114.090 101.220 ;
        RECT 116.470 100.890 116.640 101.220 ;
        RECT 114.260 100.675 116.300 100.845 ;
        RECT 113.920 100.300 114.090 100.630 ;
        RECT 116.470 100.300 116.640 100.630 ;
        RECT 114.260 100.085 116.300 100.255 ;
        RECT 113.410 94.965 113.580 99.905 ;
        RECT 113.920 99.710 114.090 100.040 ;
        RECT 116.470 99.710 116.640 100.040 ;
        RECT 114.260 99.495 116.300 99.665 ;
        RECT 113.920 99.120 114.090 99.450 ;
        RECT 116.470 99.120 116.640 99.450 ;
        RECT 114.260 98.905 116.300 99.075 ;
        RECT 113.920 98.530 114.090 98.860 ;
        RECT 116.470 98.530 116.640 98.860 ;
        RECT 114.260 98.315 116.300 98.485 ;
        RECT 113.920 97.940 114.090 98.270 ;
        RECT 116.470 97.940 116.640 98.270 ;
        RECT 114.260 97.725 116.300 97.895 ;
        RECT 113.920 97.350 114.090 97.680 ;
        RECT 116.470 97.350 116.640 97.680 ;
        RECT 114.260 97.135 116.300 97.305 ;
        RECT 113.920 96.760 114.090 97.090 ;
        RECT 116.470 96.760 116.640 97.090 ;
        RECT 114.260 96.545 116.300 96.715 ;
        RECT 113.920 96.170 114.090 96.500 ;
        RECT 116.470 96.170 116.640 96.500 ;
        RECT 114.260 95.955 116.300 96.125 ;
        RECT 113.920 95.580 114.090 95.910 ;
        RECT 116.470 95.580 116.640 95.910 ;
        RECT 114.260 95.365 116.300 95.535 ;
        RECT 116.980 94.965 117.150 107.735 ;
        RECT 113.410 94.795 117.150 94.965 ;
        RECT 107.680 89.975 110.420 90.145 ;
        RECT 107.690 87.695 110.430 87.865 ;
        RECT 107.690 83.245 107.860 87.695 ;
        RECT 108.540 87.125 109.580 87.295 ;
        RECT 108.200 85.065 108.370 87.065 ;
        RECT 109.750 85.065 109.920 87.065 ;
        RECT 108.540 84.835 109.580 85.005 ;
        RECT 107.530 82.105 107.960 83.245 ;
        RECT 108.200 82.775 108.370 84.775 ;
        RECT 109.750 82.775 109.920 84.775 ;
        RECT 108.540 82.545 109.580 82.715 ;
        RECT 107.690 69.295 107.860 82.105 ;
        RECT 108.200 80.485 108.370 82.485 ;
        RECT 109.750 80.485 109.920 82.485 ;
        RECT 108.540 80.255 109.580 80.425 ;
        RECT 108.200 78.195 108.370 80.195 ;
        RECT 109.750 78.195 109.920 80.195 ;
        RECT 108.540 77.965 109.580 78.135 ;
        RECT 108.200 75.905 108.370 77.905 ;
        RECT 109.750 75.905 109.920 77.905 ;
        RECT 108.540 75.675 109.580 75.845 ;
        RECT 108.200 73.615 108.370 75.615 ;
        RECT 109.750 73.615 109.920 75.615 ;
        RECT 108.540 73.385 109.580 73.555 ;
        RECT 108.200 71.325 108.370 73.325 ;
        RECT 109.750 71.325 109.920 73.325 ;
        RECT 108.540 71.095 109.580 71.265 ;
        RECT 107.540 68.155 107.950 69.295 ;
        RECT 108.200 69.035 108.370 71.035 ;
        RECT 109.750 69.035 109.920 71.035 ;
        RECT 108.540 68.805 109.580 68.975 ;
        RECT 107.690 63.825 107.860 68.155 ;
        RECT 108.200 66.745 108.370 68.745 ;
        RECT 109.750 66.745 109.920 68.745 ;
        RECT 108.540 66.515 109.580 66.685 ;
        RECT 108.200 64.455 108.370 66.455 ;
        RECT 109.750 64.455 109.920 66.455 ;
        RECT 108.540 64.225 109.580 64.395 ;
        RECT 110.260 63.825 110.430 87.695 ;
        RECT 120.780 81.355 120.950 108.125 ;
        RECT 121.675 107.555 124.215 107.725 ;
        RECT 125.355 107.555 127.895 107.725 ;
        RECT 129.035 107.555 131.575 107.725 ;
        RECT 132.715 107.555 135.255 107.725 ;
        RECT 136.395 107.555 138.935 107.725 ;
        RECT 140.075 107.555 142.615 107.725 ;
        RECT 143.755 107.555 146.295 107.725 ;
        RECT 121.290 106.495 121.460 107.495 ;
        RECT 124.430 106.495 124.600 107.495 ;
        RECT 124.970 106.495 125.140 107.495 ;
        RECT 128.110 106.495 128.280 107.495 ;
        RECT 128.650 106.495 128.820 107.495 ;
        RECT 131.790 106.495 131.960 107.495 ;
        RECT 132.330 106.495 132.500 107.495 ;
        RECT 135.470 106.495 135.640 107.495 ;
        RECT 136.010 106.495 136.180 107.495 ;
        RECT 139.150 106.495 139.320 107.495 ;
        RECT 139.690 106.495 139.860 107.495 ;
        RECT 142.830 106.495 143.000 107.495 ;
        RECT 143.370 106.495 143.540 107.495 ;
        RECT 146.510 106.495 146.680 107.495 ;
        RECT 121.675 106.265 124.215 106.435 ;
        RECT 125.355 106.265 127.895 106.435 ;
        RECT 129.035 106.265 131.575 106.435 ;
        RECT 132.715 106.265 135.255 106.435 ;
        RECT 136.395 106.265 138.935 106.435 ;
        RECT 140.075 106.265 142.615 106.435 ;
        RECT 143.755 106.265 146.295 106.435 ;
        RECT 147.020 106.215 147.190 108.125 ;
        RECT 121.290 105.205 121.460 106.205 ;
        RECT 124.430 105.205 124.600 106.205 ;
        RECT 124.970 105.205 125.140 106.205 ;
        RECT 128.110 105.205 128.280 106.205 ;
        RECT 128.650 105.205 128.820 106.205 ;
        RECT 131.790 105.205 131.960 106.205 ;
        RECT 132.330 105.205 132.500 106.205 ;
        RECT 135.470 105.205 135.640 106.205 ;
        RECT 136.010 105.205 136.180 106.205 ;
        RECT 139.150 105.205 139.320 106.205 ;
        RECT 139.690 105.205 139.860 106.205 ;
        RECT 142.830 105.205 143.000 106.205 ;
        RECT 143.370 105.205 143.540 106.205 ;
        RECT 146.510 105.205 146.680 106.205 ;
        RECT 121.675 104.975 124.215 105.145 ;
        RECT 125.355 104.975 127.895 105.145 ;
        RECT 129.035 104.975 131.575 105.145 ;
        RECT 132.715 104.975 135.255 105.145 ;
        RECT 136.395 104.975 138.935 105.145 ;
        RECT 140.075 104.975 142.615 105.145 ;
        RECT 143.755 104.975 146.295 105.145 ;
        RECT 121.290 103.915 121.460 104.915 ;
        RECT 124.430 103.915 124.600 104.915 ;
        RECT 124.970 103.915 125.140 104.915 ;
        RECT 128.110 103.915 128.280 104.915 ;
        RECT 128.650 103.915 128.820 104.915 ;
        RECT 131.790 103.915 131.960 104.915 ;
        RECT 132.330 103.915 132.500 104.915 ;
        RECT 135.470 103.915 135.640 104.915 ;
        RECT 136.010 103.915 136.180 104.915 ;
        RECT 139.150 103.915 139.320 104.915 ;
        RECT 139.690 103.915 139.860 104.915 ;
        RECT 142.830 103.915 143.000 104.915 ;
        RECT 143.370 103.915 143.540 104.915 ;
        RECT 146.510 103.915 146.680 104.915 ;
        RECT 146.950 104.875 147.300 106.215 ;
        RECT 121.675 103.685 124.215 103.855 ;
        RECT 125.355 103.685 127.895 103.855 ;
        RECT 129.035 103.685 131.575 103.855 ;
        RECT 132.715 103.685 135.255 103.855 ;
        RECT 136.395 103.685 138.935 103.855 ;
        RECT 140.075 103.685 142.615 103.855 ;
        RECT 143.755 103.685 146.295 103.855 ;
        RECT 121.290 102.625 121.460 103.625 ;
        RECT 124.430 102.625 124.600 103.625 ;
        RECT 124.970 102.625 125.140 103.625 ;
        RECT 128.110 102.625 128.280 103.625 ;
        RECT 128.650 102.625 128.820 103.625 ;
        RECT 131.790 102.625 131.960 103.625 ;
        RECT 132.330 102.625 132.500 103.625 ;
        RECT 135.470 102.625 135.640 103.625 ;
        RECT 136.010 102.625 136.180 103.625 ;
        RECT 139.150 102.625 139.320 103.625 ;
        RECT 139.690 102.625 139.860 103.625 ;
        RECT 142.830 102.625 143.000 103.625 ;
        RECT 143.370 102.625 143.540 103.625 ;
        RECT 146.510 102.625 146.680 103.625 ;
        RECT 121.675 102.395 124.215 102.565 ;
        RECT 125.355 102.395 127.895 102.565 ;
        RECT 129.035 102.395 131.575 102.565 ;
        RECT 132.715 102.395 135.255 102.565 ;
        RECT 136.395 102.395 138.935 102.565 ;
        RECT 140.075 102.395 142.615 102.565 ;
        RECT 143.755 102.395 146.295 102.565 ;
        RECT 121.290 101.335 121.460 102.335 ;
        RECT 124.430 101.335 124.600 102.335 ;
        RECT 124.970 101.335 125.140 102.335 ;
        RECT 128.110 101.335 128.280 102.335 ;
        RECT 128.650 101.335 128.820 102.335 ;
        RECT 131.790 101.335 131.960 102.335 ;
        RECT 132.330 101.335 132.500 102.335 ;
        RECT 135.470 101.335 135.640 102.335 ;
        RECT 136.010 101.335 136.180 102.335 ;
        RECT 139.150 101.335 139.320 102.335 ;
        RECT 139.690 101.335 139.860 102.335 ;
        RECT 142.830 101.335 143.000 102.335 ;
        RECT 143.370 101.335 143.540 102.335 ;
        RECT 146.510 101.335 146.680 102.335 ;
        RECT 121.675 101.105 124.215 101.275 ;
        RECT 125.355 101.105 127.895 101.275 ;
        RECT 129.035 101.105 131.575 101.275 ;
        RECT 132.715 101.105 135.255 101.275 ;
        RECT 136.395 101.105 138.935 101.275 ;
        RECT 140.075 101.105 142.615 101.275 ;
        RECT 143.755 101.105 146.295 101.275 ;
        RECT 121.290 100.045 121.460 101.045 ;
        RECT 124.430 100.045 124.600 101.045 ;
        RECT 124.970 100.045 125.140 101.045 ;
        RECT 128.110 100.045 128.280 101.045 ;
        RECT 128.650 100.045 128.820 101.045 ;
        RECT 131.790 100.045 131.960 101.045 ;
        RECT 132.330 100.045 132.500 101.045 ;
        RECT 135.470 100.045 135.640 101.045 ;
        RECT 136.010 100.045 136.180 101.045 ;
        RECT 139.150 100.045 139.320 101.045 ;
        RECT 139.690 100.045 139.860 101.045 ;
        RECT 142.830 100.045 143.000 101.045 ;
        RECT 143.370 100.045 143.540 101.045 ;
        RECT 146.510 100.045 146.680 101.045 ;
        RECT 121.675 99.815 124.215 99.985 ;
        RECT 125.355 99.815 127.895 99.985 ;
        RECT 129.035 99.815 131.575 99.985 ;
        RECT 132.715 99.815 135.255 99.985 ;
        RECT 136.395 99.815 138.935 99.985 ;
        RECT 140.075 99.815 142.615 99.985 ;
        RECT 143.755 99.815 146.295 99.985 ;
        RECT 121.290 98.755 121.460 99.755 ;
        RECT 124.430 98.755 124.600 99.755 ;
        RECT 124.970 98.755 125.140 99.755 ;
        RECT 128.110 98.755 128.280 99.755 ;
        RECT 128.650 98.755 128.820 99.755 ;
        RECT 131.790 98.755 131.960 99.755 ;
        RECT 132.330 98.755 132.500 99.755 ;
        RECT 135.470 98.755 135.640 99.755 ;
        RECT 136.010 98.755 136.180 99.755 ;
        RECT 139.150 98.755 139.320 99.755 ;
        RECT 139.690 98.755 139.860 99.755 ;
        RECT 142.830 98.755 143.000 99.755 ;
        RECT 143.370 98.755 143.540 99.755 ;
        RECT 146.510 98.755 146.680 99.755 ;
        RECT 121.675 98.525 124.215 98.695 ;
        RECT 125.355 98.525 127.895 98.695 ;
        RECT 129.035 98.525 131.575 98.695 ;
        RECT 132.715 98.525 135.255 98.695 ;
        RECT 136.395 98.525 138.935 98.695 ;
        RECT 140.075 98.525 142.615 98.695 ;
        RECT 143.755 98.525 146.295 98.695 ;
        RECT 121.290 97.465 121.460 98.465 ;
        RECT 124.430 97.465 124.600 98.465 ;
        RECT 124.970 97.465 125.140 98.465 ;
        RECT 128.110 97.465 128.280 98.465 ;
        RECT 128.650 97.465 128.820 98.465 ;
        RECT 131.790 97.465 131.960 98.465 ;
        RECT 132.330 97.465 132.500 98.465 ;
        RECT 135.470 97.465 135.640 98.465 ;
        RECT 136.010 97.465 136.180 98.465 ;
        RECT 139.150 97.465 139.320 98.465 ;
        RECT 139.690 97.465 139.860 98.465 ;
        RECT 142.830 97.465 143.000 98.465 ;
        RECT 143.370 97.465 143.540 98.465 ;
        RECT 146.510 97.465 146.680 98.465 ;
        RECT 121.675 97.235 124.215 97.405 ;
        RECT 125.355 97.235 127.895 97.405 ;
        RECT 129.035 97.235 131.575 97.405 ;
        RECT 132.715 97.235 135.255 97.405 ;
        RECT 136.395 97.235 138.935 97.405 ;
        RECT 140.075 97.235 142.615 97.405 ;
        RECT 143.755 97.235 146.295 97.405 ;
        RECT 121.290 96.175 121.460 97.175 ;
        RECT 124.430 96.175 124.600 97.175 ;
        RECT 124.970 96.175 125.140 97.175 ;
        RECT 128.110 96.175 128.280 97.175 ;
        RECT 128.650 96.175 128.820 97.175 ;
        RECT 131.790 96.175 131.960 97.175 ;
        RECT 132.330 96.175 132.500 97.175 ;
        RECT 135.470 96.175 135.640 97.175 ;
        RECT 136.010 96.175 136.180 97.175 ;
        RECT 139.150 96.175 139.320 97.175 ;
        RECT 139.690 96.175 139.860 97.175 ;
        RECT 142.830 96.175 143.000 97.175 ;
        RECT 143.370 96.175 143.540 97.175 ;
        RECT 146.510 96.175 146.680 97.175 ;
        RECT 121.675 95.945 124.215 96.115 ;
        RECT 125.355 95.945 127.895 96.115 ;
        RECT 129.035 95.945 131.575 96.115 ;
        RECT 132.715 95.945 135.255 96.115 ;
        RECT 136.395 95.945 138.935 96.115 ;
        RECT 140.075 95.945 142.615 96.115 ;
        RECT 143.755 95.945 146.295 96.115 ;
        RECT 121.290 94.885 121.460 95.885 ;
        RECT 124.430 94.885 124.600 95.885 ;
        RECT 124.970 94.885 125.140 95.885 ;
        RECT 128.110 94.885 128.280 95.885 ;
        RECT 128.650 94.885 128.820 95.885 ;
        RECT 131.790 94.885 131.960 95.885 ;
        RECT 132.330 94.885 132.500 95.885 ;
        RECT 135.470 94.885 135.640 95.885 ;
        RECT 136.010 94.885 136.180 95.885 ;
        RECT 139.150 94.885 139.320 95.885 ;
        RECT 139.690 94.885 139.860 95.885 ;
        RECT 142.830 94.885 143.000 95.885 ;
        RECT 143.370 94.885 143.540 95.885 ;
        RECT 146.510 94.885 146.680 95.885 ;
        RECT 121.675 94.655 124.215 94.825 ;
        RECT 125.355 94.655 127.895 94.825 ;
        RECT 129.035 94.655 131.575 94.825 ;
        RECT 132.715 94.655 135.255 94.825 ;
        RECT 136.395 94.655 138.935 94.825 ;
        RECT 140.075 94.655 142.615 94.825 ;
        RECT 143.755 94.655 146.295 94.825 ;
        RECT 121.290 93.595 121.460 94.595 ;
        RECT 124.430 93.595 124.600 94.595 ;
        RECT 124.970 93.595 125.140 94.595 ;
        RECT 128.110 93.595 128.280 94.595 ;
        RECT 128.650 93.595 128.820 94.595 ;
        RECT 131.790 93.595 131.960 94.595 ;
        RECT 132.330 93.595 132.500 94.595 ;
        RECT 135.470 93.595 135.640 94.595 ;
        RECT 136.010 93.595 136.180 94.595 ;
        RECT 139.150 93.595 139.320 94.595 ;
        RECT 139.690 93.595 139.860 94.595 ;
        RECT 142.830 93.595 143.000 94.595 ;
        RECT 143.370 93.595 143.540 94.595 ;
        RECT 146.510 93.595 146.680 94.595 ;
        RECT 121.675 93.365 124.215 93.535 ;
        RECT 125.355 93.365 127.895 93.535 ;
        RECT 129.035 93.365 131.575 93.535 ;
        RECT 132.715 93.365 135.255 93.535 ;
        RECT 136.395 93.365 138.935 93.535 ;
        RECT 140.075 93.365 142.615 93.535 ;
        RECT 143.755 93.365 146.295 93.535 ;
        RECT 121.290 92.305 121.460 93.305 ;
        RECT 124.430 92.305 124.600 93.305 ;
        RECT 124.970 92.305 125.140 93.305 ;
        RECT 128.110 92.305 128.280 93.305 ;
        RECT 128.650 92.305 128.820 93.305 ;
        RECT 131.790 92.305 131.960 93.305 ;
        RECT 132.330 92.305 132.500 93.305 ;
        RECT 135.470 92.305 135.640 93.305 ;
        RECT 136.010 92.305 136.180 93.305 ;
        RECT 139.150 92.305 139.320 93.305 ;
        RECT 139.690 92.305 139.860 93.305 ;
        RECT 142.830 92.305 143.000 93.305 ;
        RECT 143.370 92.305 143.540 93.305 ;
        RECT 146.510 92.305 146.680 93.305 ;
        RECT 121.675 92.075 124.215 92.245 ;
        RECT 125.355 92.075 127.895 92.245 ;
        RECT 129.035 92.075 131.575 92.245 ;
        RECT 132.715 92.075 135.255 92.245 ;
        RECT 136.395 92.075 138.935 92.245 ;
        RECT 140.075 92.075 142.615 92.245 ;
        RECT 143.755 92.075 146.295 92.245 ;
        RECT 121.290 91.015 121.460 92.015 ;
        RECT 124.430 91.015 124.600 92.015 ;
        RECT 124.970 91.015 125.140 92.015 ;
        RECT 128.110 91.015 128.280 92.015 ;
        RECT 128.650 91.015 128.820 92.015 ;
        RECT 131.790 91.015 131.960 92.015 ;
        RECT 132.330 91.015 132.500 92.015 ;
        RECT 135.470 91.015 135.640 92.015 ;
        RECT 136.010 91.015 136.180 92.015 ;
        RECT 139.150 91.015 139.320 92.015 ;
        RECT 139.690 91.015 139.860 92.015 ;
        RECT 142.830 91.015 143.000 92.015 ;
        RECT 143.370 91.015 143.540 92.015 ;
        RECT 146.510 91.015 146.680 92.015 ;
        RECT 121.675 90.785 124.215 90.955 ;
        RECT 125.355 90.785 127.895 90.955 ;
        RECT 129.035 90.785 131.575 90.955 ;
        RECT 132.715 90.785 135.255 90.955 ;
        RECT 136.395 90.785 138.935 90.955 ;
        RECT 140.075 90.785 142.615 90.955 ;
        RECT 143.755 90.785 146.295 90.955 ;
        RECT 121.290 89.725 121.460 90.725 ;
        RECT 124.430 89.725 124.600 90.725 ;
        RECT 124.970 89.725 125.140 90.725 ;
        RECT 128.110 89.725 128.280 90.725 ;
        RECT 128.650 89.725 128.820 90.725 ;
        RECT 131.790 89.725 131.960 90.725 ;
        RECT 132.330 89.725 132.500 90.725 ;
        RECT 135.470 89.725 135.640 90.725 ;
        RECT 136.010 89.725 136.180 90.725 ;
        RECT 139.150 89.725 139.320 90.725 ;
        RECT 139.690 89.725 139.860 90.725 ;
        RECT 142.830 89.725 143.000 90.725 ;
        RECT 143.370 89.725 143.540 90.725 ;
        RECT 146.510 89.725 146.680 90.725 ;
        RECT 121.675 89.495 124.215 89.665 ;
        RECT 125.355 89.495 127.895 89.665 ;
        RECT 129.035 89.495 131.575 89.665 ;
        RECT 132.715 89.495 135.255 89.665 ;
        RECT 136.395 89.495 138.935 89.665 ;
        RECT 140.075 89.495 142.615 89.665 ;
        RECT 143.755 89.495 146.295 89.665 ;
        RECT 121.290 88.435 121.460 89.435 ;
        RECT 124.430 88.435 124.600 89.435 ;
        RECT 124.970 88.435 125.140 89.435 ;
        RECT 128.110 88.435 128.280 89.435 ;
        RECT 128.650 88.435 128.820 89.435 ;
        RECT 131.790 88.435 131.960 89.435 ;
        RECT 132.330 88.435 132.500 89.435 ;
        RECT 135.470 88.435 135.640 89.435 ;
        RECT 136.010 88.435 136.180 89.435 ;
        RECT 139.150 88.435 139.320 89.435 ;
        RECT 139.690 88.435 139.860 89.435 ;
        RECT 142.830 88.435 143.000 89.435 ;
        RECT 143.370 88.435 143.540 89.435 ;
        RECT 146.510 88.435 146.680 89.435 ;
        RECT 121.675 88.205 124.215 88.375 ;
        RECT 125.355 88.205 127.895 88.375 ;
        RECT 129.035 88.205 131.575 88.375 ;
        RECT 132.715 88.205 135.255 88.375 ;
        RECT 136.395 88.205 138.935 88.375 ;
        RECT 140.075 88.205 142.615 88.375 ;
        RECT 143.755 88.205 146.295 88.375 ;
        RECT 121.290 87.145 121.460 88.145 ;
        RECT 124.430 87.145 124.600 88.145 ;
        RECT 124.970 87.145 125.140 88.145 ;
        RECT 128.110 87.145 128.280 88.145 ;
        RECT 128.650 87.145 128.820 88.145 ;
        RECT 131.790 87.145 131.960 88.145 ;
        RECT 132.330 87.145 132.500 88.145 ;
        RECT 135.470 87.145 135.640 88.145 ;
        RECT 136.010 87.145 136.180 88.145 ;
        RECT 139.150 87.145 139.320 88.145 ;
        RECT 139.690 87.145 139.860 88.145 ;
        RECT 142.830 87.145 143.000 88.145 ;
        RECT 143.370 87.145 143.540 88.145 ;
        RECT 146.510 87.145 146.680 88.145 ;
        RECT 121.675 86.915 124.215 87.085 ;
        RECT 125.355 86.915 127.895 87.085 ;
        RECT 129.035 86.915 131.575 87.085 ;
        RECT 132.715 86.915 135.255 87.085 ;
        RECT 136.395 86.915 138.935 87.085 ;
        RECT 140.075 86.915 142.615 87.085 ;
        RECT 143.755 86.915 146.295 87.085 ;
        RECT 121.290 85.855 121.460 86.855 ;
        RECT 124.430 85.855 124.600 86.855 ;
        RECT 124.970 85.855 125.140 86.855 ;
        RECT 128.110 85.855 128.280 86.855 ;
        RECT 128.650 85.855 128.820 86.855 ;
        RECT 131.790 85.855 131.960 86.855 ;
        RECT 132.330 85.855 132.500 86.855 ;
        RECT 135.470 85.855 135.640 86.855 ;
        RECT 136.010 85.855 136.180 86.855 ;
        RECT 139.150 85.855 139.320 86.855 ;
        RECT 139.690 85.855 139.860 86.855 ;
        RECT 142.830 85.855 143.000 86.855 ;
        RECT 143.370 85.855 143.540 86.855 ;
        RECT 146.510 85.855 146.680 86.855 ;
        RECT 121.675 85.625 124.215 85.795 ;
        RECT 125.355 85.625 127.895 85.795 ;
        RECT 129.035 85.625 131.575 85.795 ;
        RECT 132.715 85.625 135.255 85.795 ;
        RECT 136.395 85.625 138.935 85.795 ;
        RECT 140.075 85.625 142.615 85.795 ;
        RECT 143.755 85.625 146.295 85.795 ;
        RECT 121.290 84.565 121.460 85.565 ;
        RECT 124.430 84.565 124.600 85.565 ;
        RECT 124.970 84.565 125.140 85.565 ;
        RECT 128.110 84.565 128.280 85.565 ;
        RECT 128.650 84.565 128.820 85.565 ;
        RECT 131.790 84.565 131.960 85.565 ;
        RECT 132.330 84.565 132.500 85.565 ;
        RECT 135.470 84.565 135.640 85.565 ;
        RECT 136.010 84.565 136.180 85.565 ;
        RECT 139.150 84.565 139.320 85.565 ;
        RECT 139.690 84.565 139.860 85.565 ;
        RECT 142.830 84.565 143.000 85.565 ;
        RECT 143.370 84.565 143.540 85.565 ;
        RECT 146.510 84.565 146.680 85.565 ;
        RECT 147.020 85.465 147.190 104.875 ;
        RECT 121.675 84.335 124.215 84.505 ;
        RECT 125.355 84.335 127.895 84.505 ;
        RECT 129.035 84.335 131.575 84.505 ;
        RECT 132.715 84.335 135.255 84.505 ;
        RECT 136.395 84.335 138.935 84.505 ;
        RECT 140.075 84.335 142.615 84.505 ;
        RECT 143.755 84.335 146.295 84.505 ;
        RECT 121.290 83.275 121.460 84.275 ;
        RECT 124.430 83.275 124.600 84.275 ;
        RECT 124.970 83.275 125.140 84.275 ;
        RECT 128.110 83.275 128.280 84.275 ;
        RECT 128.650 83.275 128.820 84.275 ;
        RECT 131.790 83.275 131.960 84.275 ;
        RECT 132.330 83.275 132.500 84.275 ;
        RECT 135.470 83.275 135.640 84.275 ;
        RECT 136.010 83.275 136.180 84.275 ;
        RECT 139.150 83.275 139.320 84.275 ;
        RECT 139.690 83.275 139.860 84.275 ;
        RECT 142.830 83.275 143.000 84.275 ;
        RECT 143.370 83.275 143.540 84.275 ;
        RECT 146.510 83.275 146.680 84.275 ;
        RECT 146.940 83.945 147.310 85.465 ;
        RECT 121.675 83.045 124.215 83.215 ;
        RECT 125.355 83.045 127.895 83.215 ;
        RECT 129.035 83.045 131.575 83.215 ;
        RECT 132.715 83.045 135.255 83.215 ;
        RECT 136.395 83.045 138.935 83.215 ;
        RECT 140.075 83.045 142.615 83.215 ;
        RECT 143.755 83.045 146.295 83.215 ;
        RECT 121.290 81.985 121.460 82.985 ;
        RECT 124.430 81.985 124.600 82.985 ;
        RECT 124.970 81.985 125.140 82.985 ;
        RECT 128.110 81.985 128.280 82.985 ;
        RECT 128.650 81.985 128.820 82.985 ;
        RECT 131.790 81.985 131.960 82.985 ;
        RECT 132.330 81.985 132.500 82.985 ;
        RECT 135.470 81.985 135.640 82.985 ;
        RECT 136.010 81.985 136.180 82.985 ;
        RECT 139.150 81.985 139.320 82.985 ;
        RECT 139.690 81.985 139.860 82.985 ;
        RECT 142.830 81.985 143.000 82.985 ;
        RECT 143.370 81.985 143.540 82.985 ;
        RECT 146.510 81.985 146.680 82.985 ;
        RECT 121.675 81.755 124.215 81.925 ;
        RECT 125.355 81.755 127.895 81.925 ;
        RECT 129.035 81.755 131.575 81.925 ;
        RECT 132.715 81.755 135.255 81.925 ;
        RECT 136.395 81.755 138.935 81.925 ;
        RECT 140.075 81.755 142.615 81.925 ;
        RECT 143.755 81.755 146.295 81.925 ;
        RECT 147.020 81.355 147.190 83.945 ;
        RECT 120.780 81.185 147.190 81.355 ;
        RECT 107.690 63.655 110.430 63.825 ;
        RECT 120.780 77.765 147.190 77.935 ;
        RECT 107.690 61.885 110.430 62.055 ;
        RECT 107.690 57.475 107.860 61.885 ;
        RECT 108.540 61.315 109.580 61.485 ;
        RECT 108.200 59.255 108.370 61.255 ;
        RECT 109.750 59.255 109.920 61.255 ;
        RECT 108.540 59.025 109.580 59.195 ;
        RECT 107.570 56.215 107.950 57.475 ;
        RECT 108.200 56.965 108.370 58.965 ;
        RECT 109.750 56.965 109.920 58.965 ;
        RECT 108.540 56.735 109.580 56.905 ;
        RECT 107.690 43.405 107.860 56.215 ;
        RECT 108.200 54.675 108.370 56.675 ;
        RECT 109.750 54.675 109.920 56.675 ;
        RECT 108.540 54.445 109.580 54.615 ;
        RECT 108.200 52.385 108.370 54.385 ;
        RECT 109.750 52.385 109.920 54.385 ;
        RECT 108.540 52.155 109.580 52.325 ;
        RECT 108.200 50.095 108.370 52.095 ;
        RECT 109.750 50.095 109.920 52.095 ;
        RECT 108.540 49.865 109.580 50.035 ;
        RECT 108.200 47.805 108.370 49.805 ;
        RECT 109.750 47.805 109.920 49.805 ;
        RECT 108.540 47.575 109.580 47.745 ;
        RECT 108.200 45.515 108.370 47.515 ;
        RECT 109.750 45.515 109.920 47.515 ;
        RECT 108.540 45.285 109.580 45.455 ;
        RECT 107.550 42.215 107.950 43.405 ;
        RECT 108.200 43.225 108.370 45.225 ;
        RECT 109.750 43.225 109.920 45.225 ;
        RECT 108.540 42.995 109.580 43.165 ;
        RECT 107.690 38.015 107.860 42.215 ;
        RECT 108.200 40.935 108.370 42.935 ;
        RECT 109.750 40.935 109.920 42.935 ;
        RECT 108.540 40.705 109.580 40.875 ;
        RECT 108.200 38.645 108.370 40.645 ;
        RECT 109.750 38.645 109.920 40.645 ;
        RECT 108.540 38.415 109.580 38.585 ;
        RECT 110.260 38.015 110.430 61.885 ;
        RECT 120.780 50.995 120.950 77.765 ;
        RECT 121.675 77.195 124.215 77.365 ;
        RECT 125.355 77.195 127.895 77.365 ;
        RECT 129.035 77.195 131.575 77.365 ;
        RECT 132.715 77.195 135.255 77.365 ;
        RECT 136.395 77.195 138.935 77.365 ;
        RECT 140.075 77.195 142.615 77.365 ;
        RECT 143.755 77.195 146.295 77.365 ;
        RECT 121.290 76.135 121.460 77.135 ;
        RECT 124.430 76.135 124.600 77.135 ;
        RECT 124.970 76.135 125.140 77.135 ;
        RECT 128.110 76.135 128.280 77.135 ;
        RECT 128.650 76.135 128.820 77.135 ;
        RECT 131.790 76.135 131.960 77.135 ;
        RECT 132.330 76.135 132.500 77.135 ;
        RECT 135.470 76.135 135.640 77.135 ;
        RECT 136.010 76.135 136.180 77.135 ;
        RECT 139.150 76.135 139.320 77.135 ;
        RECT 139.690 76.135 139.860 77.135 ;
        RECT 142.830 76.135 143.000 77.135 ;
        RECT 143.370 76.135 143.540 77.135 ;
        RECT 146.510 76.135 146.680 77.135 ;
        RECT 121.675 75.905 124.215 76.075 ;
        RECT 125.355 75.905 127.895 76.075 ;
        RECT 129.035 75.905 131.575 76.075 ;
        RECT 132.715 75.905 135.255 76.075 ;
        RECT 136.395 75.905 138.935 76.075 ;
        RECT 140.075 75.905 142.615 76.075 ;
        RECT 143.755 75.905 146.295 76.075 ;
        RECT 147.020 75.925 147.190 77.765 ;
        RECT 121.290 74.845 121.460 75.845 ;
        RECT 124.430 74.845 124.600 75.845 ;
        RECT 124.970 74.845 125.140 75.845 ;
        RECT 128.110 74.845 128.280 75.845 ;
        RECT 128.650 74.845 128.820 75.845 ;
        RECT 131.790 74.845 131.960 75.845 ;
        RECT 132.330 74.845 132.500 75.845 ;
        RECT 135.470 74.845 135.640 75.845 ;
        RECT 136.010 74.845 136.180 75.845 ;
        RECT 139.150 74.845 139.320 75.845 ;
        RECT 139.690 74.845 139.860 75.845 ;
        RECT 142.830 74.845 143.000 75.845 ;
        RECT 143.370 74.845 143.540 75.845 ;
        RECT 146.510 74.845 146.680 75.845 ;
        RECT 121.675 74.615 124.215 74.785 ;
        RECT 125.355 74.615 127.895 74.785 ;
        RECT 129.035 74.615 131.575 74.785 ;
        RECT 132.715 74.615 135.255 74.785 ;
        RECT 136.395 74.615 138.935 74.785 ;
        RECT 140.075 74.615 142.615 74.785 ;
        RECT 143.755 74.615 146.295 74.785 ;
        RECT 121.290 73.555 121.460 74.555 ;
        RECT 124.430 73.555 124.600 74.555 ;
        RECT 124.970 73.555 125.140 74.555 ;
        RECT 128.110 73.555 128.280 74.555 ;
        RECT 128.650 73.555 128.820 74.555 ;
        RECT 131.790 73.555 131.960 74.555 ;
        RECT 132.330 73.555 132.500 74.555 ;
        RECT 135.470 73.555 135.640 74.555 ;
        RECT 136.010 73.555 136.180 74.555 ;
        RECT 139.150 73.555 139.320 74.555 ;
        RECT 139.690 73.555 139.860 74.555 ;
        RECT 142.830 73.555 143.000 74.555 ;
        RECT 143.370 73.555 143.540 74.555 ;
        RECT 146.510 73.555 146.680 74.555 ;
        RECT 146.950 74.485 147.300 75.925 ;
        RECT 121.675 73.325 124.215 73.495 ;
        RECT 125.355 73.325 127.895 73.495 ;
        RECT 129.035 73.325 131.575 73.495 ;
        RECT 132.715 73.325 135.255 73.495 ;
        RECT 136.395 73.325 138.935 73.495 ;
        RECT 140.075 73.325 142.615 73.495 ;
        RECT 143.755 73.325 146.295 73.495 ;
        RECT 121.290 72.265 121.460 73.265 ;
        RECT 124.430 72.265 124.600 73.265 ;
        RECT 124.970 72.265 125.140 73.265 ;
        RECT 128.110 72.265 128.280 73.265 ;
        RECT 128.650 72.265 128.820 73.265 ;
        RECT 131.790 72.265 131.960 73.265 ;
        RECT 132.330 72.265 132.500 73.265 ;
        RECT 135.470 72.265 135.640 73.265 ;
        RECT 136.010 72.265 136.180 73.265 ;
        RECT 139.150 72.265 139.320 73.265 ;
        RECT 139.690 72.265 139.860 73.265 ;
        RECT 142.830 72.265 143.000 73.265 ;
        RECT 143.370 72.265 143.540 73.265 ;
        RECT 146.510 72.265 146.680 73.265 ;
        RECT 121.675 72.035 124.215 72.205 ;
        RECT 125.355 72.035 127.895 72.205 ;
        RECT 129.035 72.035 131.575 72.205 ;
        RECT 132.715 72.035 135.255 72.205 ;
        RECT 136.395 72.035 138.935 72.205 ;
        RECT 140.075 72.035 142.615 72.205 ;
        RECT 143.755 72.035 146.295 72.205 ;
        RECT 121.290 70.975 121.460 71.975 ;
        RECT 124.430 70.975 124.600 71.975 ;
        RECT 124.970 70.975 125.140 71.975 ;
        RECT 128.110 70.975 128.280 71.975 ;
        RECT 128.650 70.975 128.820 71.975 ;
        RECT 131.790 70.975 131.960 71.975 ;
        RECT 132.330 70.975 132.500 71.975 ;
        RECT 135.470 70.975 135.640 71.975 ;
        RECT 136.010 70.975 136.180 71.975 ;
        RECT 139.150 70.975 139.320 71.975 ;
        RECT 139.690 70.975 139.860 71.975 ;
        RECT 142.830 70.975 143.000 71.975 ;
        RECT 143.370 70.975 143.540 71.975 ;
        RECT 146.510 70.975 146.680 71.975 ;
        RECT 121.675 70.745 124.215 70.915 ;
        RECT 125.355 70.745 127.895 70.915 ;
        RECT 129.035 70.745 131.575 70.915 ;
        RECT 132.715 70.745 135.255 70.915 ;
        RECT 136.395 70.745 138.935 70.915 ;
        RECT 140.075 70.745 142.615 70.915 ;
        RECT 143.755 70.745 146.295 70.915 ;
        RECT 121.290 69.685 121.460 70.685 ;
        RECT 124.430 69.685 124.600 70.685 ;
        RECT 124.970 69.685 125.140 70.685 ;
        RECT 128.110 69.685 128.280 70.685 ;
        RECT 128.650 69.685 128.820 70.685 ;
        RECT 131.790 69.685 131.960 70.685 ;
        RECT 132.330 69.685 132.500 70.685 ;
        RECT 135.470 69.685 135.640 70.685 ;
        RECT 136.010 69.685 136.180 70.685 ;
        RECT 139.150 69.685 139.320 70.685 ;
        RECT 139.690 69.685 139.860 70.685 ;
        RECT 142.830 69.685 143.000 70.685 ;
        RECT 143.370 69.685 143.540 70.685 ;
        RECT 146.510 69.685 146.680 70.685 ;
        RECT 121.675 69.455 124.215 69.625 ;
        RECT 125.355 69.455 127.895 69.625 ;
        RECT 129.035 69.455 131.575 69.625 ;
        RECT 132.715 69.455 135.255 69.625 ;
        RECT 136.395 69.455 138.935 69.625 ;
        RECT 140.075 69.455 142.615 69.625 ;
        RECT 143.755 69.455 146.295 69.625 ;
        RECT 121.290 68.395 121.460 69.395 ;
        RECT 124.430 68.395 124.600 69.395 ;
        RECT 124.970 68.395 125.140 69.395 ;
        RECT 128.110 68.395 128.280 69.395 ;
        RECT 128.650 68.395 128.820 69.395 ;
        RECT 131.790 68.395 131.960 69.395 ;
        RECT 132.330 68.395 132.500 69.395 ;
        RECT 135.470 68.395 135.640 69.395 ;
        RECT 136.010 68.395 136.180 69.395 ;
        RECT 139.150 68.395 139.320 69.395 ;
        RECT 139.690 68.395 139.860 69.395 ;
        RECT 142.830 68.395 143.000 69.395 ;
        RECT 143.370 68.395 143.540 69.395 ;
        RECT 146.510 68.395 146.680 69.395 ;
        RECT 121.675 68.165 124.215 68.335 ;
        RECT 125.355 68.165 127.895 68.335 ;
        RECT 129.035 68.165 131.575 68.335 ;
        RECT 132.715 68.165 135.255 68.335 ;
        RECT 136.395 68.165 138.935 68.335 ;
        RECT 140.075 68.165 142.615 68.335 ;
        RECT 143.755 68.165 146.295 68.335 ;
        RECT 121.290 67.105 121.460 68.105 ;
        RECT 124.430 67.105 124.600 68.105 ;
        RECT 124.970 67.105 125.140 68.105 ;
        RECT 128.110 67.105 128.280 68.105 ;
        RECT 128.650 67.105 128.820 68.105 ;
        RECT 131.790 67.105 131.960 68.105 ;
        RECT 132.330 67.105 132.500 68.105 ;
        RECT 135.470 67.105 135.640 68.105 ;
        RECT 136.010 67.105 136.180 68.105 ;
        RECT 139.150 67.105 139.320 68.105 ;
        RECT 139.690 67.105 139.860 68.105 ;
        RECT 142.830 67.105 143.000 68.105 ;
        RECT 143.370 67.105 143.540 68.105 ;
        RECT 146.510 67.105 146.680 68.105 ;
        RECT 121.675 66.875 124.215 67.045 ;
        RECT 125.355 66.875 127.895 67.045 ;
        RECT 129.035 66.875 131.575 67.045 ;
        RECT 132.715 66.875 135.255 67.045 ;
        RECT 136.395 66.875 138.935 67.045 ;
        RECT 140.075 66.875 142.615 67.045 ;
        RECT 143.755 66.875 146.295 67.045 ;
        RECT 121.290 65.815 121.460 66.815 ;
        RECT 124.430 65.815 124.600 66.815 ;
        RECT 124.970 65.815 125.140 66.815 ;
        RECT 128.110 65.815 128.280 66.815 ;
        RECT 128.650 65.815 128.820 66.815 ;
        RECT 131.790 65.815 131.960 66.815 ;
        RECT 132.330 65.815 132.500 66.815 ;
        RECT 135.470 65.815 135.640 66.815 ;
        RECT 136.010 65.815 136.180 66.815 ;
        RECT 139.150 65.815 139.320 66.815 ;
        RECT 139.690 65.815 139.860 66.815 ;
        RECT 142.830 65.815 143.000 66.815 ;
        RECT 143.370 65.815 143.540 66.815 ;
        RECT 146.510 65.815 146.680 66.815 ;
        RECT 121.675 65.585 124.215 65.755 ;
        RECT 125.355 65.585 127.895 65.755 ;
        RECT 129.035 65.585 131.575 65.755 ;
        RECT 132.715 65.585 135.255 65.755 ;
        RECT 136.395 65.585 138.935 65.755 ;
        RECT 140.075 65.585 142.615 65.755 ;
        RECT 143.755 65.585 146.295 65.755 ;
        RECT 121.290 64.525 121.460 65.525 ;
        RECT 124.430 64.525 124.600 65.525 ;
        RECT 124.970 64.525 125.140 65.525 ;
        RECT 128.110 64.525 128.280 65.525 ;
        RECT 128.650 64.525 128.820 65.525 ;
        RECT 131.790 64.525 131.960 65.525 ;
        RECT 132.330 64.525 132.500 65.525 ;
        RECT 135.470 64.525 135.640 65.525 ;
        RECT 136.010 64.525 136.180 65.525 ;
        RECT 139.150 64.525 139.320 65.525 ;
        RECT 139.690 64.525 139.860 65.525 ;
        RECT 142.830 64.525 143.000 65.525 ;
        RECT 143.370 64.525 143.540 65.525 ;
        RECT 146.510 64.525 146.680 65.525 ;
        RECT 121.675 64.295 124.215 64.465 ;
        RECT 125.355 64.295 127.895 64.465 ;
        RECT 129.035 64.295 131.575 64.465 ;
        RECT 132.715 64.295 135.255 64.465 ;
        RECT 136.395 64.295 138.935 64.465 ;
        RECT 140.075 64.295 142.615 64.465 ;
        RECT 143.755 64.295 146.295 64.465 ;
        RECT 121.290 63.235 121.460 64.235 ;
        RECT 124.430 63.235 124.600 64.235 ;
        RECT 124.970 63.235 125.140 64.235 ;
        RECT 128.110 63.235 128.280 64.235 ;
        RECT 128.650 63.235 128.820 64.235 ;
        RECT 131.790 63.235 131.960 64.235 ;
        RECT 132.330 63.235 132.500 64.235 ;
        RECT 135.470 63.235 135.640 64.235 ;
        RECT 136.010 63.235 136.180 64.235 ;
        RECT 139.150 63.235 139.320 64.235 ;
        RECT 139.690 63.235 139.860 64.235 ;
        RECT 142.830 63.235 143.000 64.235 ;
        RECT 143.370 63.235 143.540 64.235 ;
        RECT 146.510 63.235 146.680 64.235 ;
        RECT 121.675 63.005 124.215 63.175 ;
        RECT 125.355 63.005 127.895 63.175 ;
        RECT 129.035 63.005 131.575 63.175 ;
        RECT 132.715 63.005 135.255 63.175 ;
        RECT 136.395 63.005 138.935 63.175 ;
        RECT 140.075 63.005 142.615 63.175 ;
        RECT 143.755 63.005 146.295 63.175 ;
        RECT 121.290 61.945 121.460 62.945 ;
        RECT 124.430 61.945 124.600 62.945 ;
        RECT 124.970 61.945 125.140 62.945 ;
        RECT 128.110 61.945 128.280 62.945 ;
        RECT 128.650 61.945 128.820 62.945 ;
        RECT 131.790 61.945 131.960 62.945 ;
        RECT 132.330 61.945 132.500 62.945 ;
        RECT 135.470 61.945 135.640 62.945 ;
        RECT 136.010 61.945 136.180 62.945 ;
        RECT 139.150 61.945 139.320 62.945 ;
        RECT 139.690 61.945 139.860 62.945 ;
        RECT 142.830 61.945 143.000 62.945 ;
        RECT 143.370 61.945 143.540 62.945 ;
        RECT 146.510 61.945 146.680 62.945 ;
        RECT 121.675 61.715 124.215 61.885 ;
        RECT 125.355 61.715 127.895 61.885 ;
        RECT 129.035 61.715 131.575 61.885 ;
        RECT 132.715 61.715 135.255 61.885 ;
        RECT 136.395 61.715 138.935 61.885 ;
        RECT 140.075 61.715 142.615 61.885 ;
        RECT 143.755 61.715 146.295 61.885 ;
        RECT 121.290 60.655 121.460 61.655 ;
        RECT 124.430 60.655 124.600 61.655 ;
        RECT 124.970 60.655 125.140 61.655 ;
        RECT 128.110 60.655 128.280 61.655 ;
        RECT 128.650 60.655 128.820 61.655 ;
        RECT 131.790 60.655 131.960 61.655 ;
        RECT 132.330 60.655 132.500 61.655 ;
        RECT 135.470 60.655 135.640 61.655 ;
        RECT 136.010 60.655 136.180 61.655 ;
        RECT 139.150 60.655 139.320 61.655 ;
        RECT 139.690 60.655 139.860 61.655 ;
        RECT 142.830 60.655 143.000 61.655 ;
        RECT 143.370 60.655 143.540 61.655 ;
        RECT 146.510 60.655 146.680 61.655 ;
        RECT 121.675 60.425 124.215 60.595 ;
        RECT 125.355 60.425 127.895 60.595 ;
        RECT 129.035 60.425 131.575 60.595 ;
        RECT 132.715 60.425 135.255 60.595 ;
        RECT 136.395 60.425 138.935 60.595 ;
        RECT 140.075 60.425 142.615 60.595 ;
        RECT 143.755 60.425 146.295 60.595 ;
        RECT 121.290 59.365 121.460 60.365 ;
        RECT 124.430 59.365 124.600 60.365 ;
        RECT 124.970 59.365 125.140 60.365 ;
        RECT 128.110 59.365 128.280 60.365 ;
        RECT 128.650 59.365 128.820 60.365 ;
        RECT 131.790 59.365 131.960 60.365 ;
        RECT 132.330 59.365 132.500 60.365 ;
        RECT 135.470 59.365 135.640 60.365 ;
        RECT 136.010 59.365 136.180 60.365 ;
        RECT 139.150 59.365 139.320 60.365 ;
        RECT 139.690 59.365 139.860 60.365 ;
        RECT 142.830 59.365 143.000 60.365 ;
        RECT 143.370 59.365 143.540 60.365 ;
        RECT 146.510 59.365 146.680 60.365 ;
        RECT 121.675 59.135 124.215 59.305 ;
        RECT 125.355 59.135 127.895 59.305 ;
        RECT 129.035 59.135 131.575 59.305 ;
        RECT 132.715 59.135 135.255 59.305 ;
        RECT 136.395 59.135 138.935 59.305 ;
        RECT 140.075 59.135 142.615 59.305 ;
        RECT 143.755 59.135 146.295 59.305 ;
        RECT 121.290 58.075 121.460 59.075 ;
        RECT 124.430 58.075 124.600 59.075 ;
        RECT 124.970 58.075 125.140 59.075 ;
        RECT 128.110 58.075 128.280 59.075 ;
        RECT 128.650 58.075 128.820 59.075 ;
        RECT 131.790 58.075 131.960 59.075 ;
        RECT 132.330 58.075 132.500 59.075 ;
        RECT 135.470 58.075 135.640 59.075 ;
        RECT 136.010 58.075 136.180 59.075 ;
        RECT 139.150 58.075 139.320 59.075 ;
        RECT 139.690 58.075 139.860 59.075 ;
        RECT 142.830 58.075 143.000 59.075 ;
        RECT 143.370 58.075 143.540 59.075 ;
        RECT 146.510 58.075 146.680 59.075 ;
        RECT 121.675 57.845 124.215 58.015 ;
        RECT 125.355 57.845 127.895 58.015 ;
        RECT 129.035 57.845 131.575 58.015 ;
        RECT 132.715 57.845 135.255 58.015 ;
        RECT 136.395 57.845 138.935 58.015 ;
        RECT 140.075 57.845 142.615 58.015 ;
        RECT 143.755 57.845 146.295 58.015 ;
        RECT 121.290 56.785 121.460 57.785 ;
        RECT 124.430 56.785 124.600 57.785 ;
        RECT 124.970 56.785 125.140 57.785 ;
        RECT 128.110 56.785 128.280 57.785 ;
        RECT 128.650 56.785 128.820 57.785 ;
        RECT 131.790 56.785 131.960 57.785 ;
        RECT 132.330 56.785 132.500 57.785 ;
        RECT 135.470 56.785 135.640 57.785 ;
        RECT 136.010 56.785 136.180 57.785 ;
        RECT 139.150 56.785 139.320 57.785 ;
        RECT 139.690 56.785 139.860 57.785 ;
        RECT 142.830 56.785 143.000 57.785 ;
        RECT 143.370 56.785 143.540 57.785 ;
        RECT 146.510 56.785 146.680 57.785 ;
        RECT 121.675 56.555 124.215 56.725 ;
        RECT 125.355 56.555 127.895 56.725 ;
        RECT 129.035 56.555 131.575 56.725 ;
        RECT 132.715 56.555 135.255 56.725 ;
        RECT 136.395 56.555 138.935 56.725 ;
        RECT 140.075 56.555 142.615 56.725 ;
        RECT 143.755 56.555 146.295 56.725 ;
        RECT 121.290 55.495 121.460 56.495 ;
        RECT 124.430 55.495 124.600 56.495 ;
        RECT 124.970 55.495 125.140 56.495 ;
        RECT 128.110 55.495 128.280 56.495 ;
        RECT 128.650 55.495 128.820 56.495 ;
        RECT 131.790 55.495 131.960 56.495 ;
        RECT 132.330 55.495 132.500 56.495 ;
        RECT 135.470 55.495 135.640 56.495 ;
        RECT 136.010 55.495 136.180 56.495 ;
        RECT 139.150 55.495 139.320 56.495 ;
        RECT 139.690 55.495 139.860 56.495 ;
        RECT 142.830 55.495 143.000 56.495 ;
        RECT 143.370 55.495 143.540 56.495 ;
        RECT 146.510 55.495 146.680 56.495 ;
        RECT 121.675 55.265 124.215 55.435 ;
        RECT 125.355 55.265 127.895 55.435 ;
        RECT 129.035 55.265 131.575 55.435 ;
        RECT 132.715 55.265 135.255 55.435 ;
        RECT 136.395 55.265 138.935 55.435 ;
        RECT 140.075 55.265 142.615 55.435 ;
        RECT 143.755 55.265 146.295 55.435 ;
        RECT 121.290 54.205 121.460 55.205 ;
        RECT 124.430 54.205 124.600 55.205 ;
        RECT 124.970 54.205 125.140 55.205 ;
        RECT 128.110 54.205 128.280 55.205 ;
        RECT 128.650 54.205 128.820 55.205 ;
        RECT 131.790 54.205 131.960 55.205 ;
        RECT 132.330 54.205 132.500 55.205 ;
        RECT 135.470 54.205 135.640 55.205 ;
        RECT 136.010 54.205 136.180 55.205 ;
        RECT 139.150 54.205 139.320 55.205 ;
        RECT 139.690 54.205 139.860 55.205 ;
        RECT 142.830 54.205 143.000 55.205 ;
        RECT 143.370 54.205 143.540 55.205 ;
        RECT 146.510 54.205 146.680 55.205 ;
        RECT 147.020 55.155 147.190 74.485 ;
        RECT 121.675 53.975 124.215 54.145 ;
        RECT 125.355 53.975 127.895 54.145 ;
        RECT 129.035 53.975 131.575 54.145 ;
        RECT 132.715 53.975 135.255 54.145 ;
        RECT 136.395 53.975 138.935 54.145 ;
        RECT 140.075 53.975 142.615 54.145 ;
        RECT 143.755 53.975 146.295 54.145 ;
        RECT 121.290 52.915 121.460 53.915 ;
        RECT 124.430 52.915 124.600 53.915 ;
        RECT 124.970 52.915 125.140 53.915 ;
        RECT 128.110 52.915 128.280 53.915 ;
        RECT 128.650 52.915 128.820 53.915 ;
        RECT 131.790 52.915 131.960 53.915 ;
        RECT 132.330 52.915 132.500 53.915 ;
        RECT 135.470 52.915 135.640 53.915 ;
        RECT 136.010 52.915 136.180 53.915 ;
        RECT 139.150 52.915 139.320 53.915 ;
        RECT 139.690 52.915 139.860 53.915 ;
        RECT 142.830 52.915 143.000 53.915 ;
        RECT 143.370 52.915 143.540 53.915 ;
        RECT 146.510 52.915 146.680 53.915 ;
        RECT 146.930 53.695 147.310 55.155 ;
        RECT 121.675 52.685 124.215 52.855 ;
        RECT 125.355 52.685 127.895 52.855 ;
        RECT 129.035 52.685 131.575 52.855 ;
        RECT 132.715 52.685 135.255 52.855 ;
        RECT 136.395 52.685 138.935 52.855 ;
        RECT 140.075 52.685 142.615 52.855 ;
        RECT 143.755 52.685 146.295 52.855 ;
        RECT 121.290 51.625 121.460 52.625 ;
        RECT 124.430 51.625 124.600 52.625 ;
        RECT 124.970 51.625 125.140 52.625 ;
        RECT 128.110 51.625 128.280 52.625 ;
        RECT 128.650 51.625 128.820 52.625 ;
        RECT 131.790 51.625 131.960 52.625 ;
        RECT 132.330 51.625 132.500 52.625 ;
        RECT 135.470 51.625 135.640 52.625 ;
        RECT 136.010 51.625 136.180 52.625 ;
        RECT 139.150 51.625 139.320 52.625 ;
        RECT 139.690 51.625 139.860 52.625 ;
        RECT 142.830 51.625 143.000 52.625 ;
        RECT 143.370 51.625 143.540 52.625 ;
        RECT 146.510 51.625 146.680 52.625 ;
        RECT 121.675 51.395 124.215 51.565 ;
        RECT 125.355 51.395 127.895 51.565 ;
        RECT 129.035 51.395 131.575 51.565 ;
        RECT 132.715 51.395 135.255 51.565 ;
        RECT 136.395 51.395 138.935 51.565 ;
        RECT 140.075 51.395 142.615 51.565 ;
        RECT 143.755 51.395 146.295 51.565 ;
        RECT 147.020 50.995 147.190 53.695 ;
        RECT 120.780 50.825 147.190 50.995 ;
        RECT 140.080 46.395 146.910 46.565 ;
        RECT 117.840 44.365 128.670 44.535 ;
        RECT 112.800 44.185 115.540 44.355 ;
        RECT 112.800 43.035 112.970 44.185 ;
        RECT 113.650 43.615 114.690 43.785 ;
        RECT 112.700 39.785 113.000 43.035 ;
        RECT 113.310 41.555 113.480 43.555 ;
        RECT 114.860 41.555 115.030 43.555 ;
        RECT 113.650 41.325 114.690 41.495 ;
        RECT 112.800 38.635 112.970 39.785 ;
        RECT 113.310 39.265 113.480 41.265 ;
        RECT 114.860 39.265 115.030 41.265 ;
        RECT 113.650 39.035 114.690 39.205 ;
        RECT 115.370 38.635 115.540 44.185 ;
        RECT 117.840 43.435 118.010 44.365 ;
        RECT 118.350 43.475 118.520 43.805 ;
        RECT 118.690 43.795 122.730 43.965 ;
        RECT 123.780 43.795 127.820 43.965 ;
        RECT 117.780 39.605 118.030 43.435 ;
        RECT 118.690 43.315 122.730 43.485 ;
        RECT 118.350 42.515 118.520 42.845 ;
        RECT 118.690 42.835 122.730 43.005 ;
        RECT 122.900 42.995 123.070 43.325 ;
        RECT 123.440 42.995 123.610 43.325 ;
        RECT 123.780 43.315 127.820 43.485 ;
        RECT 127.990 43.475 128.160 43.805 ;
        RECT 123.780 42.835 127.820 43.005 ;
        RECT 118.690 42.355 122.730 42.525 ;
        RECT 118.350 41.555 118.520 41.885 ;
        RECT 118.690 41.875 122.730 42.045 ;
        RECT 122.900 42.035 123.070 42.365 ;
        RECT 123.440 42.035 123.610 42.365 ;
        RECT 123.780 42.355 127.820 42.525 ;
        RECT 127.990 42.515 128.160 42.845 ;
        RECT 123.780 41.875 127.820 42.045 ;
        RECT 118.690 41.395 122.730 41.565 ;
        RECT 118.350 40.595 118.520 40.925 ;
        RECT 118.690 40.915 122.730 41.085 ;
        RECT 122.900 41.075 123.070 41.405 ;
        RECT 123.440 41.075 123.610 41.405 ;
        RECT 123.780 41.395 127.820 41.565 ;
        RECT 127.990 41.555 128.160 41.885 ;
        RECT 123.780 40.915 127.820 41.085 ;
        RECT 118.690 40.435 122.730 40.605 ;
        RECT 118.350 39.635 118.520 39.965 ;
        RECT 118.690 39.955 122.730 40.125 ;
        RECT 122.900 40.115 123.070 40.445 ;
        RECT 123.440 40.115 123.610 40.445 ;
        RECT 123.780 40.435 127.820 40.605 ;
        RECT 127.990 40.595 128.160 40.925 ;
        RECT 123.780 39.955 127.820 40.125 ;
        RECT 112.800 38.465 115.540 38.635 ;
        RECT 117.840 38.595 118.010 39.605 ;
        RECT 118.690 39.475 122.730 39.645 ;
        RECT 118.690 38.995 122.730 39.165 ;
        RECT 122.900 39.155 123.070 39.485 ;
        RECT 123.440 39.155 123.610 39.485 ;
        RECT 123.780 39.475 127.820 39.645 ;
        RECT 127.990 39.635 128.160 39.965 ;
        RECT 123.780 38.995 127.820 39.165 ;
        RECT 128.500 38.595 128.670 44.365 ;
        RECT 117.840 38.425 128.670 38.595 ;
        RECT 130.680 44.305 137.510 44.475 ;
        RECT 130.680 38.535 130.850 44.305 ;
        RECT 131.190 43.415 131.360 43.745 ;
        RECT 131.575 43.735 136.615 43.905 ;
        RECT 131.575 43.255 136.615 43.425 ;
        RECT 131.190 42.455 131.360 42.785 ;
        RECT 131.575 42.775 136.615 42.945 ;
        RECT 136.830 42.935 137.000 43.265 ;
        RECT 137.340 42.815 137.510 44.305 ;
        RECT 140.080 44.135 140.250 46.395 ;
        RECT 140.975 45.825 146.015 45.995 ;
        RECT 140.590 44.765 140.760 45.765 ;
        RECT 146.230 44.765 146.400 45.765 ;
        RECT 146.740 45.665 146.910 46.395 ;
        RECT 146.660 44.795 147.040 45.665 ;
        RECT 140.975 44.535 146.015 44.705 ;
        RECT 146.740 44.135 146.910 44.795 ;
        RECT 140.080 43.965 146.910 44.135 ;
        RECT 131.575 42.295 136.615 42.465 ;
        RECT 131.190 41.495 131.360 41.825 ;
        RECT 131.575 41.815 136.615 41.985 ;
        RECT 136.830 41.975 137.000 42.305 ;
        RECT 131.575 41.335 136.615 41.505 ;
        RECT 131.190 40.535 131.360 40.865 ;
        RECT 131.575 40.855 136.615 41.025 ;
        RECT 136.830 41.015 137.000 41.345 ;
        RECT 131.575 40.375 136.615 40.545 ;
        RECT 131.190 39.575 131.360 39.905 ;
        RECT 131.575 39.895 136.615 40.065 ;
        RECT 136.830 40.055 137.000 40.385 ;
        RECT 137.300 40.115 137.610 42.815 ;
        RECT 140.070 40.935 146.900 41.105 ;
        RECT 131.575 39.415 136.615 39.585 ;
        RECT 131.575 38.935 136.615 39.105 ;
        RECT 136.830 39.095 137.000 39.425 ;
        RECT 137.340 38.535 137.510 40.115 ;
        RECT 130.680 38.365 137.510 38.535 ;
        RECT 140.070 38.675 140.240 40.935 ;
        RECT 140.965 40.365 146.005 40.535 ;
        RECT 140.580 39.305 140.750 40.305 ;
        RECT 146.220 39.305 146.390 40.305 ;
        RECT 146.730 40.205 146.900 40.935 ;
        RECT 146.670 39.395 147.050 40.205 ;
        RECT 140.965 39.075 146.005 39.245 ;
        RECT 146.730 38.675 146.900 39.395 ;
        RECT 140.070 38.505 146.900 38.675 ;
        RECT 107.690 37.845 110.430 38.015 ;
      LAYER mcon ;
        RECT 108.620 140.815 109.500 140.985 ;
        RECT 108.200 138.835 108.370 140.675 ;
        RECT 109.750 138.835 109.920 140.675 ;
        RECT 108.620 138.525 109.500 138.695 ;
        RECT 107.480 135.805 107.940 136.845 ;
        RECT 108.200 136.545 108.370 138.385 ;
        RECT 109.750 136.545 109.920 138.385 ;
        RECT 108.620 136.235 109.500 136.405 ;
        RECT 108.200 134.255 108.370 136.095 ;
        RECT 109.750 134.255 109.920 136.095 ;
        RECT 108.620 133.945 109.500 134.115 ;
        RECT 108.200 131.965 108.370 133.805 ;
        RECT 109.750 131.965 109.920 133.805 ;
        RECT 108.620 131.655 109.500 131.825 ;
        RECT 108.200 129.675 108.370 131.515 ;
        RECT 109.750 129.675 109.920 131.515 ;
        RECT 108.620 129.365 109.500 129.535 ;
        RECT 108.200 127.385 108.370 129.225 ;
        RECT 109.750 127.385 109.920 129.225 ;
        RECT 108.620 127.075 109.500 127.245 ;
        RECT 108.200 125.095 108.370 126.935 ;
        RECT 109.750 125.095 109.920 126.935 ;
        RECT 108.620 124.785 109.500 124.955 ;
        RECT 107.500 121.805 107.940 122.965 ;
        RECT 108.200 122.805 108.370 124.645 ;
        RECT 109.750 122.805 109.920 124.645 ;
        RECT 108.620 122.495 109.500 122.665 ;
        RECT 108.200 120.515 108.370 122.355 ;
        RECT 109.750 120.515 109.920 122.355 ;
        RECT 108.620 120.205 109.500 120.375 ;
        RECT 108.200 118.225 108.370 120.065 ;
        RECT 109.750 118.225 109.920 120.065 ;
        RECT 108.620 117.915 109.500 118.085 ;
        RECT 113.930 140.815 114.810 140.985 ;
        RECT 113.510 138.835 113.680 140.675 ;
        RECT 115.060 138.835 115.230 140.675 ;
        RECT 113.930 138.525 114.810 138.695 ;
        RECT 113.510 136.545 113.680 138.385 ;
        RECT 115.060 136.545 115.230 138.385 ;
        RECT 113.930 136.235 114.810 136.405 ;
        RECT 113.510 134.255 113.680 136.095 ;
        RECT 115.060 134.255 115.230 136.095 ;
        RECT 113.930 133.945 114.810 134.115 ;
        RECT 113.510 131.965 113.680 133.805 ;
        RECT 115.060 131.965 115.230 133.805 ;
        RECT 113.930 131.655 114.810 131.825 ;
        RECT 113.510 129.675 113.680 131.515 ;
        RECT 115.060 129.675 115.230 131.515 ;
        RECT 113.930 129.365 114.810 129.535 ;
        RECT 113.510 127.385 113.680 129.225 ;
        RECT 115.060 127.385 115.230 129.225 ;
        RECT 113.930 127.075 114.810 127.245 ;
        RECT 113.510 125.095 113.680 126.935 ;
        RECT 115.060 125.095 115.230 126.935 ;
        RECT 113.930 124.785 114.810 124.955 ;
        RECT 113.510 122.805 113.680 124.645 ;
        RECT 115.060 122.805 115.230 124.645 ;
        RECT 113.930 122.495 114.810 122.665 ;
        RECT 113.510 120.515 113.680 122.355 ;
        RECT 115.060 120.515 115.230 122.355 ;
        RECT 113.930 120.205 114.810 120.375 ;
        RECT 113.510 118.225 113.680 120.065 ;
        RECT 115.060 118.225 115.230 120.065 ;
        RECT 113.930 117.915 114.810 118.085 ;
        RECT 122.780 141.135 124.765 141.325 ;
        RECT 132.775 141.135 134.760 141.325 ;
        RECT 122.780 139.175 124.765 139.365 ;
        RECT 132.775 139.175 134.760 139.365 ;
        RECT 122.780 137.205 124.765 137.395 ;
        RECT 132.775 137.205 134.760 137.395 ;
        RECT 122.780 135.215 124.765 135.405 ;
        RECT 134.775 135.215 136.760 135.405 ;
        RECT 122.780 133.195 124.765 133.385 ;
        RECT 134.775 133.195 136.760 133.385 ;
        RECT 122.780 131.225 124.765 131.415 ;
        RECT 134.775 131.225 136.760 131.415 ;
        RECT 126.410 126.645 127.290 126.815 ;
        RECT 128.500 126.645 129.380 126.815 ;
        RECT 130.590 126.645 131.470 126.815 ;
        RECT 132.680 126.645 133.560 126.815 ;
        RECT 134.770 126.645 135.650 126.815 ;
        RECT 125.990 126.350 126.160 126.520 ;
        RECT 127.540 126.350 127.710 126.520 ;
        RECT 128.080 126.350 128.250 126.520 ;
        RECT 129.630 126.350 129.800 126.520 ;
        RECT 130.170 126.350 130.340 126.520 ;
        RECT 131.720 126.350 131.890 126.520 ;
        RECT 132.260 126.350 132.430 126.520 ;
        RECT 133.810 126.350 133.980 126.520 ;
        RECT 134.350 126.350 134.520 126.520 ;
        RECT 135.900 126.350 136.070 126.520 ;
        RECT 126.410 126.055 127.290 126.225 ;
        RECT 128.500 126.055 129.380 126.225 ;
        RECT 130.590 126.055 131.470 126.225 ;
        RECT 132.680 126.055 133.560 126.225 ;
        RECT 134.770 126.055 135.650 126.225 ;
        RECT 125.990 125.760 126.160 125.930 ;
        RECT 127.540 125.760 127.710 125.930 ;
        RECT 128.080 125.760 128.250 125.930 ;
        RECT 129.630 125.760 129.800 125.930 ;
        RECT 130.170 125.760 130.340 125.930 ;
        RECT 131.720 125.760 131.890 125.930 ;
        RECT 132.260 125.760 132.430 125.930 ;
        RECT 133.810 125.760 133.980 125.930 ;
        RECT 134.350 125.760 134.520 125.930 ;
        RECT 135.900 125.760 136.070 125.930 ;
        RECT 126.410 125.465 127.290 125.635 ;
        RECT 128.500 125.465 129.380 125.635 ;
        RECT 130.590 125.465 131.470 125.635 ;
        RECT 132.680 125.465 133.560 125.635 ;
        RECT 134.770 125.465 135.650 125.635 ;
        RECT 125.990 125.170 126.160 125.340 ;
        RECT 127.540 125.170 127.710 125.340 ;
        RECT 128.080 125.170 128.250 125.340 ;
        RECT 129.630 125.170 129.800 125.340 ;
        RECT 130.170 125.170 130.340 125.340 ;
        RECT 131.720 125.170 131.890 125.340 ;
        RECT 132.260 125.170 132.430 125.340 ;
        RECT 133.810 125.170 133.980 125.340 ;
        RECT 134.350 125.170 134.520 125.340 ;
        RECT 135.900 125.170 136.070 125.340 ;
        RECT 126.410 124.875 127.290 125.045 ;
        RECT 128.500 124.875 129.380 125.045 ;
        RECT 130.590 124.875 131.470 125.045 ;
        RECT 132.680 124.875 133.560 125.045 ;
        RECT 134.770 124.875 135.650 125.045 ;
        RECT 125.990 124.580 126.160 124.750 ;
        RECT 127.540 124.580 127.710 124.750 ;
        RECT 128.080 124.580 128.250 124.750 ;
        RECT 129.630 124.580 129.800 124.750 ;
        RECT 130.170 124.580 130.340 124.750 ;
        RECT 131.720 124.580 131.890 124.750 ;
        RECT 132.260 124.580 132.430 124.750 ;
        RECT 133.810 124.580 133.980 124.750 ;
        RECT 134.350 124.580 134.520 124.750 ;
        RECT 135.900 124.580 136.070 124.750 ;
        RECT 126.410 124.285 127.290 124.455 ;
        RECT 128.500 124.285 129.380 124.455 ;
        RECT 130.590 124.285 131.470 124.455 ;
        RECT 132.680 124.285 133.560 124.455 ;
        RECT 134.770 124.285 135.650 124.455 ;
        RECT 125.400 123.065 125.690 124.255 ;
        RECT 125.990 123.990 126.160 124.160 ;
        RECT 127.540 123.990 127.710 124.160 ;
        RECT 128.080 123.990 128.250 124.160 ;
        RECT 129.630 123.990 129.800 124.160 ;
        RECT 130.170 123.990 130.340 124.160 ;
        RECT 131.720 123.990 131.890 124.160 ;
        RECT 132.260 123.990 132.430 124.160 ;
        RECT 133.810 123.990 133.980 124.160 ;
        RECT 134.350 123.990 134.520 124.160 ;
        RECT 135.900 123.990 136.070 124.160 ;
        RECT 126.410 123.695 127.290 123.865 ;
        RECT 128.500 123.695 129.380 123.865 ;
        RECT 130.590 123.695 131.470 123.865 ;
        RECT 132.680 123.695 133.560 123.865 ;
        RECT 134.770 123.695 135.650 123.865 ;
        RECT 125.990 123.400 126.160 123.570 ;
        RECT 127.540 123.400 127.710 123.570 ;
        RECT 128.080 123.400 128.250 123.570 ;
        RECT 129.630 123.400 129.800 123.570 ;
        RECT 130.170 123.400 130.340 123.570 ;
        RECT 131.720 123.400 131.890 123.570 ;
        RECT 132.260 123.400 132.430 123.570 ;
        RECT 133.810 123.400 133.980 123.570 ;
        RECT 134.350 123.400 134.520 123.570 ;
        RECT 135.900 123.400 136.070 123.570 ;
        RECT 126.410 123.105 127.290 123.275 ;
        RECT 128.500 123.105 129.380 123.275 ;
        RECT 130.590 123.105 131.470 123.275 ;
        RECT 132.680 123.105 133.560 123.275 ;
        RECT 134.770 123.105 135.650 123.275 ;
        RECT 125.990 122.810 126.160 122.980 ;
        RECT 127.540 122.810 127.710 122.980 ;
        RECT 128.080 122.810 128.250 122.980 ;
        RECT 129.630 122.810 129.800 122.980 ;
        RECT 130.170 122.810 130.340 122.980 ;
        RECT 131.720 122.810 131.890 122.980 ;
        RECT 132.260 122.810 132.430 122.980 ;
        RECT 133.810 122.810 133.980 122.980 ;
        RECT 134.350 122.810 134.520 122.980 ;
        RECT 135.900 122.810 136.070 122.980 ;
        RECT 126.410 122.515 127.290 122.685 ;
        RECT 128.500 122.515 129.380 122.685 ;
        RECT 130.590 122.515 131.470 122.685 ;
        RECT 132.680 122.515 133.560 122.685 ;
        RECT 134.770 122.515 135.650 122.685 ;
        RECT 125.990 122.220 126.160 122.390 ;
        RECT 127.540 122.220 127.710 122.390 ;
        RECT 128.080 122.220 128.250 122.390 ;
        RECT 129.630 122.220 129.800 122.390 ;
        RECT 130.170 122.220 130.340 122.390 ;
        RECT 131.720 122.220 131.890 122.390 ;
        RECT 132.260 122.220 132.430 122.390 ;
        RECT 133.810 122.220 133.980 122.390 ;
        RECT 134.350 122.220 134.520 122.390 ;
        RECT 135.900 122.220 136.070 122.390 ;
        RECT 126.410 121.925 127.290 122.095 ;
        RECT 128.500 121.925 129.380 122.095 ;
        RECT 130.590 121.925 131.470 122.095 ;
        RECT 132.680 121.925 133.560 122.095 ;
        RECT 134.770 121.925 135.650 122.095 ;
        RECT 125.990 121.630 126.160 121.800 ;
        RECT 127.540 121.630 127.710 121.800 ;
        RECT 128.080 121.630 128.250 121.800 ;
        RECT 129.630 121.630 129.800 121.800 ;
        RECT 130.170 121.630 130.340 121.800 ;
        RECT 131.720 121.630 131.890 121.800 ;
        RECT 132.260 121.630 132.430 121.800 ;
        RECT 133.810 121.630 133.980 121.800 ;
        RECT 134.350 121.630 134.520 121.800 ;
        RECT 135.900 121.630 136.070 121.800 ;
        RECT 126.410 121.335 127.290 121.505 ;
        RECT 128.500 121.335 129.380 121.505 ;
        RECT 130.590 121.335 131.470 121.505 ;
        RECT 132.680 121.335 133.560 121.505 ;
        RECT 134.770 121.335 135.650 121.505 ;
        RECT 125.990 121.040 126.160 121.210 ;
        RECT 127.540 121.040 127.710 121.210 ;
        RECT 128.080 121.040 128.250 121.210 ;
        RECT 129.630 121.040 129.800 121.210 ;
        RECT 130.170 121.040 130.340 121.210 ;
        RECT 131.720 121.040 131.890 121.210 ;
        RECT 132.260 121.040 132.430 121.210 ;
        RECT 133.810 121.040 133.980 121.210 ;
        RECT 134.350 121.040 134.520 121.210 ;
        RECT 135.900 121.040 136.070 121.210 ;
        RECT 126.410 120.745 127.290 120.915 ;
        RECT 128.500 120.745 129.380 120.915 ;
        RECT 130.590 120.745 131.470 120.915 ;
        RECT 132.680 120.745 133.560 120.915 ;
        RECT 134.770 120.745 135.650 120.915 ;
        RECT 145.245 127.905 146.125 128.075 ;
        RECT 144.780 126.925 144.950 127.765 ;
        RECT 146.420 126.925 146.590 127.765 ;
        RECT 145.245 126.615 146.125 126.785 ;
        RECT 144.780 125.635 144.950 126.475 ;
        RECT 146.420 125.635 146.590 126.475 ;
        RECT 145.245 125.325 146.125 125.495 ;
        RECT 144.780 124.345 144.950 125.185 ;
        RECT 146.420 124.345 146.590 125.185 ;
        RECT 146.860 124.225 147.210 125.275 ;
        RECT 145.245 124.035 146.125 124.205 ;
        RECT 144.780 123.055 144.950 123.895 ;
        RECT 146.420 123.055 146.590 123.895 ;
        RECT 145.245 122.745 146.125 122.915 ;
        RECT 144.780 121.765 144.950 122.605 ;
        RECT 146.420 121.765 146.590 122.605 ;
        RECT 145.245 121.455 146.125 121.625 ;
        RECT 126.410 119.105 127.290 119.275 ;
        RECT 128.500 119.105 129.380 119.275 ;
        RECT 130.590 119.105 131.470 119.275 ;
        RECT 132.680 119.105 133.560 119.275 ;
        RECT 134.770 119.105 135.650 119.275 ;
        RECT 125.990 118.810 126.160 118.980 ;
        RECT 127.540 118.810 127.710 118.980 ;
        RECT 128.080 118.810 128.250 118.980 ;
        RECT 129.630 118.810 129.800 118.980 ;
        RECT 130.170 118.810 130.340 118.980 ;
        RECT 131.720 118.810 131.890 118.980 ;
        RECT 132.260 118.810 132.430 118.980 ;
        RECT 133.810 118.810 133.980 118.980 ;
        RECT 134.350 118.810 134.520 118.980 ;
        RECT 135.900 118.810 136.070 118.980 ;
        RECT 126.410 118.515 127.290 118.685 ;
        RECT 128.500 118.515 129.380 118.685 ;
        RECT 130.590 118.515 131.470 118.685 ;
        RECT 132.680 118.515 133.560 118.685 ;
        RECT 134.770 118.515 135.650 118.685 ;
        RECT 125.990 118.220 126.160 118.390 ;
        RECT 127.540 118.220 127.710 118.390 ;
        RECT 128.080 118.220 128.250 118.390 ;
        RECT 129.630 118.220 129.800 118.390 ;
        RECT 130.170 118.220 130.340 118.390 ;
        RECT 131.720 118.220 131.890 118.390 ;
        RECT 132.260 118.220 132.430 118.390 ;
        RECT 133.810 118.220 133.980 118.390 ;
        RECT 134.350 118.220 134.520 118.390 ;
        RECT 135.900 118.220 136.070 118.390 ;
        RECT 126.410 117.925 127.290 118.095 ;
        RECT 128.500 117.925 129.380 118.095 ;
        RECT 130.590 117.925 131.470 118.095 ;
        RECT 132.680 117.925 133.560 118.095 ;
        RECT 134.770 117.925 135.650 118.095 ;
        RECT 125.990 117.630 126.160 117.800 ;
        RECT 127.540 117.630 127.710 117.800 ;
        RECT 128.080 117.630 128.250 117.800 ;
        RECT 129.630 117.630 129.800 117.800 ;
        RECT 130.170 117.630 130.340 117.800 ;
        RECT 131.720 117.630 131.890 117.800 ;
        RECT 132.260 117.630 132.430 117.800 ;
        RECT 133.810 117.630 133.980 117.800 ;
        RECT 134.350 117.630 134.520 117.800 ;
        RECT 135.900 117.630 136.070 117.800 ;
        RECT 126.410 117.335 127.290 117.505 ;
        RECT 128.500 117.335 129.380 117.505 ;
        RECT 130.590 117.335 131.470 117.505 ;
        RECT 132.680 117.335 133.560 117.505 ;
        RECT 134.770 117.335 135.650 117.505 ;
        RECT 125.990 117.040 126.160 117.210 ;
        RECT 127.540 117.040 127.710 117.210 ;
        RECT 128.080 117.040 128.250 117.210 ;
        RECT 129.630 117.040 129.800 117.210 ;
        RECT 130.170 117.040 130.340 117.210 ;
        RECT 131.720 117.040 131.890 117.210 ;
        RECT 132.260 117.040 132.430 117.210 ;
        RECT 133.810 117.040 133.980 117.210 ;
        RECT 134.350 117.040 134.520 117.210 ;
        RECT 135.900 117.040 136.070 117.210 ;
        RECT 125.390 115.655 125.700 116.865 ;
        RECT 126.410 116.745 127.290 116.915 ;
        RECT 128.500 116.745 129.380 116.915 ;
        RECT 130.590 116.745 131.470 116.915 ;
        RECT 132.680 116.745 133.560 116.915 ;
        RECT 134.770 116.745 135.650 116.915 ;
        RECT 125.990 116.450 126.160 116.620 ;
        RECT 127.540 116.450 127.710 116.620 ;
        RECT 128.080 116.450 128.250 116.620 ;
        RECT 129.630 116.450 129.800 116.620 ;
        RECT 130.170 116.450 130.340 116.620 ;
        RECT 131.720 116.450 131.890 116.620 ;
        RECT 132.260 116.450 132.430 116.620 ;
        RECT 133.810 116.450 133.980 116.620 ;
        RECT 134.350 116.450 134.520 116.620 ;
        RECT 135.900 116.450 136.070 116.620 ;
        RECT 126.410 116.155 127.290 116.325 ;
        RECT 128.500 116.155 129.380 116.325 ;
        RECT 130.590 116.155 131.470 116.325 ;
        RECT 132.680 116.155 133.560 116.325 ;
        RECT 134.770 116.155 135.650 116.325 ;
        RECT 125.990 115.860 126.160 116.030 ;
        RECT 127.540 115.860 127.710 116.030 ;
        RECT 128.080 115.860 128.250 116.030 ;
        RECT 129.630 115.860 129.800 116.030 ;
        RECT 130.170 115.860 130.340 116.030 ;
        RECT 131.720 115.860 131.890 116.030 ;
        RECT 132.260 115.860 132.430 116.030 ;
        RECT 133.810 115.860 133.980 116.030 ;
        RECT 134.350 115.860 134.520 116.030 ;
        RECT 135.900 115.860 136.070 116.030 ;
        RECT 108.610 113.445 109.490 113.615 ;
        RECT 108.190 111.465 108.360 113.305 ;
        RECT 109.740 111.465 109.910 113.305 ;
        RECT 108.610 111.155 109.490 111.325 ;
        RECT 107.530 108.265 107.960 109.455 ;
        RECT 108.190 109.175 108.360 111.015 ;
        RECT 109.740 109.175 109.910 111.015 ;
        RECT 108.610 108.865 109.490 109.035 ;
        RECT 108.190 106.885 108.360 108.725 ;
        RECT 109.740 106.885 109.910 108.725 ;
        RECT 108.610 106.575 109.490 106.745 ;
        RECT 108.190 104.595 108.360 106.435 ;
        RECT 109.740 104.595 109.910 106.435 ;
        RECT 108.610 104.285 109.490 104.455 ;
        RECT 108.190 102.305 108.360 104.145 ;
        RECT 109.740 102.305 109.910 104.145 ;
        RECT 108.610 101.995 109.490 102.165 ;
        RECT 108.190 100.015 108.360 101.855 ;
        RECT 109.740 100.015 109.910 101.855 ;
        RECT 108.610 99.705 109.490 99.875 ;
        RECT 108.190 97.725 108.360 99.565 ;
        RECT 109.740 97.725 109.910 99.565 ;
        RECT 108.610 97.415 109.490 97.585 ;
        RECT 107.530 94.535 107.950 95.735 ;
        RECT 108.190 95.435 108.360 97.275 ;
        RECT 109.740 95.435 109.910 97.275 ;
        RECT 108.610 95.125 109.490 95.295 ;
        RECT 108.190 93.145 108.360 94.985 ;
        RECT 109.740 93.145 109.910 94.985 ;
        RECT 108.610 92.835 109.490 93.005 ;
        RECT 108.190 90.855 108.360 92.695 ;
        RECT 109.740 90.855 109.910 92.695 ;
        RECT 108.610 90.545 109.490 90.715 ;
        RECT 126.410 115.565 127.290 115.735 ;
        RECT 128.500 115.565 129.380 115.735 ;
        RECT 130.590 115.565 131.470 115.735 ;
        RECT 132.680 115.565 133.560 115.735 ;
        RECT 134.770 115.565 135.650 115.735 ;
        RECT 125.990 115.270 126.160 115.440 ;
        RECT 127.540 115.270 127.710 115.440 ;
        RECT 128.080 115.270 128.250 115.440 ;
        RECT 129.630 115.270 129.800 115.440 ;
        RECT 130.170 115.270 130.340 115.440 ;
        RECT 131.720 115.270 131.890 115.440 ;
        RECT 132.260 115.270 132.430 115.440 ;
        RECT 133.810 115.270 133.980 115.440 ;
        RECT 134.350 115.270 134.520 115.440 ;
        RECT 135.900 115.270 136.070 115.440 ;
        RECT 126.410 114.975 127.290 115.145 ;
        RECT 128.500 114.975 129.380 115.145 ;
        RECT 130.590 114.975 131.470 115.145 ;
        RECT 132.680 114.975 133.560 115.145 ;
        RECT 134.770 114.975 135.650 115.145 ;
        RECT 125.990 114.680 126.160 114.850 ;
        RECT 127.540 114.680 127.710 114.850 ;
        RECT 128.080 114.680 128.250 114.850 ;
        RECT 129.630 114.680 129.800 114.850 ;
        RECT 130.170 114.680 130.340 114.850 ;
        RECT 131.720 114.680 131.890 114.850 ;
        RECT 132.260 114.680 132.430 114.850 ;
        RECT 133.810 114.680 133.980 114.850 ;
        RECT 134.350 114.680 134.520 114.850 ;
        RECT 135.900 114.680 136.070 114.850 ;
        RECT 126.410 114.385 127.290 114.555 ;
        RECT 128.500 114.385 129.380 114.555 ;
        RECT 130.590 114.385 131.470 114.555 ;
        RECT 132.680 114.385 133.560 114.555 ;
        RECT 134.770 114.385 135.650 114.555 ;
        RECT 125.990 114.090 126.160 114.260 ;
        RECT 127.540 114.090 127.710 114.260 ;
        RECT 128.080 114.090 128.250 114.260 ;
        RECT 129.630 114.090 129.800 114.260 ;
        RECT 130.170 114.090 130.340 114.260 ;
        RECT 131.720 114.090 131.890 114.260 ;
        RECT 132.260 114.090 132.430 114.260 ;
        RECT 133.810 114.090 133.980 114.260 ;
        RECT 134.350 114.090 134.520 114.260 ;
        RECT 135.900 114.090 136.070 114.260 ;
        RECT 126.410 113.795 127.290 113.965 ;
        RECT 128.500 113.795 129.380 113.965 ;
        RECT 130.590 113.795 131.470 113.965 ;
        RECT 132.680 113.795 133.560 113.965 ;
        RECT 134.770 113.795 135.650 113.965 ;
        RECT 125.990 113.500 126.160 113.670 ;
        RECT 127.540 113.500 127.710 113.670 ;
        RECT 128.080 113.500 128.250 113.670 ;
        RECT 129.630 113.500 129.800 113.670 ;
        RECT 130.170 113.500 130.340 113.670 ;
        RECT 131.720 113.500 131.890 113.670 ;
        RECT 132.260 113.500 132.430 113.670 ;
        RECT 133.810 113.500 133.980 113.670 ;
        RECT 134.350 113.500 134.520 113.670 ;
        RECT 135.900 113.500 136.070 113.670 ;
        RECT 126.410 113.205 127.290 113.375 ;
        RECT 128.500 113.205 129.380 113.375 ;
        RECT 130.590 113.205 131.470 113.375 ;
        RECT 132.680 113.205 133.560 113.375 ;
        RECT 134.770 113.205 135.650 113.375 ;
        RECT 145.215 118.125 146.095 118.295 ;
        RECT 144.750 117.145 144.920 117.985 ;
        RECT 146.390 117.145 146.560 117.985 ;
        RECT 145.215 116.835 146.095 117.005 ;
        RECT 144.750 115.855 144.920 116.695 ;
        RECT 146.390 115.855 146.560 116.695 ;
        RECT 145.215 115.545 146.095 115.715 ;
        RECT 144.750 114.565 144.920 115.405 ;
        RECT 146.390 114.565 146.560 115.405 ;
        RECT 146.850 114.425 147.190 115.385 ;
        RECT 145.215 114.255 146.095 114.425 ;
        RECT 144.750 113.275 144.920 114.115 ;
        RECT 146.390 113.275 146.560 114.115 ;
        RECT 145.215 112.965 146.095 113.135 ;
        RECT 144.750 111.985 144.920 112.825 ;
        RECT 146.390 111.985 146.560 112.825 ;
        RECT 145.215 111.675 146.095 111.845 ;
        RECT 114.340 107.165 116.220 107.335 ;
        RECT 113.920 106.870 114.090 107.040 ;
        RECT 116.470 106.870 116.640 107.040 ;
        RECT 114.340 106.575 116.220 106.745 ;
        RECT 113.920 106.280 114.090 106.450 ;
        RECT 116.470 106.280 116.640 106.450 ;
        RECT 114.340 105.985 116.220 106.155 ;
        RECT 113.920 105.690 114.090 105.860 ;
        RECT 116.470 105.690 116.640 105.860 ;
        RECT 114.340 105.395 116.220 105.565 ;
        RECT 113.920 105.100 114.090 105.270 ;
        RECT 116.470 105.100 116.640 105.270 ;
        RECT 114.340 104.805 116.220 104.975 ;
        RECT 113.920 104.510 114.090 104.680 ;
        RECT 116.470 104.510 116.640 104.680 ;
        RECT 114.340 104.215 116.220 104.385 ;
        RECT 113.920 103.920 114.090 104.090 ;
        RECT 116.470 103.920 116.640 104.090 ;
        RECT 114.340 103.625 116.220 103.795 ;
        RECT 113.280 99.905 113.600 103.615 ;
        RECT 113.920 103.330 114.090 103.500 ;
        RECT 116.470 103.330 116.640 103.500 ;
        RECT 114.340 103.035 116.220 103.205 ;
        RECT 113.920 102.740 114.090 102.910 ;
        RECT 116.470 102.740 116.640 102.910 ;
        RECT 114.340 102.445 116.220 102.615 ;
        RECT 113.920 102.150 114.090 102.320 ;
        RECT 116.470 102.150 116.640 102.320 ;
        RECT 114.340 101.855 116.220 102.025 ;
        RECT 113.920 101.560 114.090 101.730 ;
        RECT 116.470 101.560 116.640 101.730 ;
        RECT 114.340 101.265 116.220 101.435 ;
        RECT 113.920 100.970 114.090 101.140 ;
        RECT 116.470 100.970 116.640 101.140 ;
        RECT 114.340 100.675 116.220 100.845 ;
        RECT 113.920 100.380 114.090 100.550 ;
        RECT 116.470 100.380 116.640 100.550 ;
        RECT 114.340 100.085 116.220 100.255 ;
        RECT 113.920 99.790 114.090 99.960 ;
        RECT 116.470 99.790 116.640 99.960 ;
        RECT 114.340 99.495 116.220 99.665 ;
        RECT 113.920 99.200 114.090 99.370 ;
        RECT 116.470 99.200 116.640 99.370 ;
        RECT 114.340 98.905 116.220 99.075 ;
        RECT 113.920 98.610 114.090 98.780 ;
        RECT 116.470 98.610 116.640 98.780 ;
        RECT 114.340 98.315 116.220 98.485 ;
        RECT 113.920 98.020 114.090 98.190 ;
        RECT 116.470 98.020 116.640 98.190 ;
        RECT 114.340 97.725 116.220 97.895 ;
        RECT 113.920 97.430 114.090 97.600 ;
        RECT 116.470 97.430 116.640 97.600 ;
        RECT 114.340 97.135 116.220 97.305 ;
        RECT 113.920 96.840 114.090 97.010 ;
        RECT 116.470 96.840 116.640 97.010 ;
        RECT 114.340 96.545 116.220 96.715 ;
        RECT 113.920 96.250 114.090 96.420 ;
        RECT 116.470 96.250 116.640 96.420 ;
        RECT 114.340 95.955 116.220 96.125 ;
        RECT 113.920 95.660 114.090 95.830 ;
        RECT 116.470 95.660 116.640 95.830 ;
        RECT 114.340 95.365 116.220 95.535 ;
        RECT 108.620 87.125 109.500 87.295 ;
        RECT 108.200 85.145 108.370 86.985 ;
        RECT 109.750 85.145 109.920 86.985 ;
        RECT 108.620 84.835 109.500 85.005 ;
        RECT 107.530 82.105 107.960 83.245 ;
        RECT 108.200 82.855 108.370 84.695 ;
        RECT 109.750 82.855 109.920 84.695 ;
        RECT 108.620 82.545 109.500 82.715 ;
        RECT 108.200 80.565 108.370 82.405 ;
        RECT 109.750 80.565 109.920 82.405 ;
        RECT 108.620 80.255 109.500 80.425 ;
        RECT 108.200 78.275 108.370 80.115 ;
        RECT 109.750 78.275 109.920 80.115 ;
        RECT 108.620 77.965 109.500 78.135 ;
        RECT 108.200 75.985 108.370 77.825 ;
        RECT 109.750 75.985 109.920 77.825 ;
        RECT 108.620 75.675 109.500 75.845 ;
        RECT 108.200 73.695 108.370 75.535 ;
        RECT 109.750 73.695 109.920 75.535 ;
        RECT 108.620 73.385 109.500 73.555 ;
        RECT 108.200 71.405 108.370 73.245 ;
        RECT 109.750 71.405 109.920 73.245 ;
        RECT 108.620 71.095 109.500 71.265 ;
        RECT 107.540 68.155 107.950 69.295 ;
        RECT 108.200 69.115 108.370 70.955 ;
        RECT 109.750 69.115 109.920 70.955 ;
        RECT 108.620 68.805 109.500 68.975 ;
        RECT 108.200 66.825 108.370 68.665 ;
        RECT 109.750 66.825 109.920 68.665 ;
        RECT 108.620 66.515 109.500 66.685 ;
        RECT 108.200 64.535 108.370 66.375 ;
        RECT 109.750 64.535 109.920 66.375 ;
        RECT 108.620 64.225 109.500 64.395 ;
        RECT 121.755 107.555 124.135 107.725 ;
        RECT 125.435 107.555 127.815 107.725 ;
        RECT 129.115 107.555 131.495 107.725 ;
        RECT 132.795 107.555 135.175 107.725 ;
        RECT 136.475 107.555 138.855 107.725 ;
        RECT 140.155 107.555 142.535 107.725 ;
        RECT 143.835 107.555 146.215 107.725 ;
        RECT 121.290 106.575 121.460 107.415 ;
        RECT 124.430 106.575 124.600 107.415 ;
        RECT 124.970 106.575 125.140 107.415 ;
        RECT 128.110 106.575 128.280 107.415 ;
        RECT 128.650 106.575 128.820 107.415 ;
        RECT 131.790 106.575 131.960 107.415 ;
        RECT 132.330 106.575 132.500 107.415 ;
        RECT 135.470 106.575 135.640 107.415 ;
        RECT 136.010 106.575 136.180 107.415 ;
        RECT 139.150 106.575 139.320 107.415 ;
        RECT 139.690 106.575 139.860 107.415 ;
        RECT 142.830 106.575 143.000 107.415 ;
        RECT 143.370 106.575 143.540 107.415 ;
        RECT 146.510 106.575 146.680 107.415 ;
        RECT 121.755 106.265 124.135 106.435 ;
        RECT 125.435 106.265 127.815 106.435 ;
        RECT 129.115 106.265 131.495 106.435 ;
        RECT 132.795 106.265 135.175 106.435 ;
        RECT 136.475 106.265 138.855 106.435 ;
        RECT 140.155 106.265 142.535 106.435 ;
        RECT 143.835 106.265 146.215 106.435 ;
        RECT 121.290 105.285 121.460 106.125 ;
        RECT 124.430 105.285 124.600 106.125 ;
        RECT 124.970 105.285 125.140 106.125 ;
        RECT 128.110 105.285 128.280 106.125 ;
        RECT 128.650 105.285 128.820 106.125 ;
        RECT 131.790 105.285 131.960 106.125 ;
        RECT 132.330 105.285 132.500 106.125 ;
        RECT 135.470 105.285 135.640 106.125 ;
        RECT 136.010 105.285 136.180 106.125 ;
        RECT 139.150 105.285 139.320 106.125 ;
        RECT 139.690 105.285 139.860 106.125 ;
        RECT 142.830 105.285 143.000 106.125 ;
        RECT 143.370 105.285 143.540 106.125 ;
        RECT 146.510 105.285 146.680 106.125 ;
        RECT 121.755 104.975 124.135 105.145 ;
        RECT 125.435 104.975 127.815 105.145 ;
        RECT 129.115 104.975 131.495 105.145 ;
        RECT 132.795 104.975 135.175 105.145 ;
        RECT 136.475 104.975 138.855 105.145 ;
        RECT 140.155 104.975 142.535 105.145 ;
        RECT 143.835 104.975 146.215 105.145 ;
        RECT 121.290 103.995 121.460 104.835 ;
        RECT 124.430 103.995 124.600 104.835 ;
        RECT 124.970 103.995 125.140 104.835 ;
        RECT 128.110 103.995 128.280 104.835 ;
        RECT 128.650 103.995 128.820 104.835 ;
        RECT 131.790 103.995 131.960 104.835 ;
        RECT 132.330 103.995 132.500 104.835 ;
        RECT 135.470 103.995 135.640 104.835 ;
        RECT 136.010 103.995 136.180 104.835 ;
        RECT 139.150 103.995 139.320 104.835 ;
        RECT 139.690 103.995 139.860 104.835 ;
        RECT 142.830 103.995 143.000 104.835 ;
        RECT 143.370 103.995 143.540 104.835 ;
        RECT 146.950 104.875 147.300 106.215 ;
        RECT 146.510 103.995 146.680 104.835 ;
        RECT 121.755 103.685 124.135 103.855 ;
        RECT 125.435 103.685 127.815 103.855 ;
        RECT 129.115 103.685 131.495 103.855 ;
        RECT 132.795 103.685 135.175 103.855 ;
        RECT 136.475 103.685 138.855 103.855 ;
        RECT 140.155 103.685 142.535 103.855 ;
        RECT 143.835 103.685 146.215 103.855 ;
        RECT 121.290 102.705 121.460 103.545 ;
        RECT 124.430 102.705 124.600 103.545 ;
        RECT 124.970 102.705 125.140 103.545 ;
        RECT 128.110 102.705 128.280 103.545 ;
        RECT 128.650 102.705 128.820 103.545 ;
        RECT 131.790 102.705 131.960 103.545 ;
        RECT 132.330 102.705 132.500 103.545 ;
        RECT 135.470 102.705 135.640 103.545 ;
        RECT 136.010 102.705 136.180 103.545 ;
        RECT 139.150 102.705 139.320 103.545 ;
        RECT 139.690 102.705 139.860 103.545 ;
        RECT 142.830 102.705 143.000 103.545 ;
        RECT 143.370 102.705 143.540 103.545 ;
        RECT 146.510 102.705 146.680 103.545 ;
        RECT 121.755 102.395 124.135 102.565 ;
        RECT 125.435 102.395 127.815 102.565 ;
        RECT 129.115 102.395 131.495 102.565 ;
        RECT 132.795 102.395 135.175 102.565 ;
        RECT 136.475 102.395 138.855 102.565 ;
        RECT 140.155 102.395 142.535 102.565 ;
        RECT 143.835 102.395 146.215 102.565 ;
        RECT 121.290 101.415 121.460 102.255 ;
        RECT 124.430 101.415 124.600 102.255 ;
        RECT 124.970 101.415 125.140 102.255 ;
        RECT 128.110 101.415 128.280 102.255 ;
        RECT 128.650 101.415 128.820 102.255 ;
        RECT 131.790 101.415 131.960 102.255 ;
        RECT 132.330 101.415 132.500 102.255 ;
        RECT 135.470 101.415 135.640 102.255 ;
        RECT 136.010 101.415 136.180 102.255 ;
        RECT 139.150 101.415 139.320 102.255 ;
        RECT 139.690 101.415 139.860 102.255 ;
        RECT 142.830 101.415 143.000 102.255 ;
        RECT 143.370 101.415 143.540 102.255 ;
        RECT 146.510 101.415 146.680 102.255 ;
        RECT 121.755 101.105 124.135 101.275 ;
        RECT 125.435 101.105 127.815 101.275 ;
        RECT 129.115 101.105 131.495 101.275 ;
        RECT 132.795 101.105 135.175 101.275 ;
        RECT 136.475 101.105 138.855 101.275 ;
        RECT 140.155 101.105 142.535 101.275 ;
        RECT 143.835 101.105 146.215 101.275 ;
        RECT 121.290 100.125 121.460 100.965 ;
        RECT 124.430 100.125 124.600 100.965 ;
        RECT 124.970 100.125 125.140 100.965 ;
        RECT 128.110 100.125 128.280 100.965 ;
        RECT 128.650 100.125 128.820 100.965 ;
        RECT 131.790 100.125 131.960 100.965 ;
        RECT 132.330 100.125 132.500 100.965 ;
        RECT 135.470 100.125 135.640 100.965 ;
        RECT 136.010 100.125 136.180 100.965 ;
        RECT 139.150 100.125 139.320 100.965 ;
        RECT 139.690 100.125 139.860 100.965 ;
        RECT 142.830 100.125 143.000 100.965 ;
        RECT 143.370 100.125 143.540 100.965 ;
        RECT 146.510 100.125 146.680 100.965 ;
        RECT 121.755 99.815 124.135 99.985 ;
        RECT 125.435 99.815 127.815 99.985 ;
        RECT 129.115 99.815 131.495 99.985 ;
        RECT 132.795 99.815 135.175 99.985 ;
        RECT 136.475 99.815 138.855 99.985 ;
        RECT 140.155 99.815 142.535 99.985 ;
        RECT 143.835 99.815 146.215 99.985 ;
        RECT 121.290 98.835 121.460 99.675 ;
        RECT 124.430 98.835 124.600 99.675 ;
        RECT 124.970 98.835 125.140 99.675 ;
        RECT 128.110 98.835 128.280 99.675 ;
        RECT 128.650 98.835 128.820 99.675 ;
        RECT 131.790 98.835 131.960 99.675 ;
        RECT 132.330 98.835 132.500 99.675 ;
        RECT 135.470 98.835 135.640 99.675 ;
        RECT 136.010 98.835 136.180 99.675 ;
        RECT 139.150 98.835 139.320 99.675 ;
        RECT 139.690 98.835 139.860 99.675 ;
        RECT 142.830 98.835 143.000 99.675 ;
        RECT 143.370 98.835 143.540 99.675 ;
        RECT 146.510 98.835 146.680 99.675 ;
        RECT 121.755 98.525 124.135 98.695 ;
        RECT 125.435 98.525 127.815 98.695 ;
        RECT 129.115 98.525 131.495 98.695 ;
        RECT 132.795 98.525 135.175 98.695 ;
        RECT 136.475 98.525 138.855 98.695 ;
        RECT 140.155 98.525 142.535 98.695 ;
        RECT 143.835 98.525 146.215 98.695 ;
        RECT 121.290 97.545 121.460 98.385 ;
        RECT 124.430 97.545 124.600 98.385 ;
        RECT 124.970 97.545 125.140 98.385 ;
        RECT 128.110 97.545 128.280 98.385 ;
        RECT 128.650 97.545 128.820 98.385 ;
        RECT 131.790 97.545 131.960 98.385 ;
        RECT 132.330 97.545 132.500 98.385 ;
        RECT 135.470 97.545 135.640 98.385 ;
        RECT 136.010 97.545 136.180 98.385 ;
        RECT 139.150 97.545 139.320 98.385 ;
        RECT 139.690 97.545 139.860 98.385 ;
        RECT 142.830 97.545 143.000 98.385 ;
        RECT 143.370 97.545 143.540 98.385 ;
        RECT 146.510 97.545 146.680 98.385 ;
        RECT 121.755 97.235 124.135 97.405 ;
        RECT 125.435 97.235 127.815 97.405 ;
        RECT 129.115 97.235 131.495 97.405 ;
        RECT 132.795 97.235 135.175 97.405 ;
        RECT 136.475 97.235 138.855 97.405 ;
        RECT 140.155 97.235 142.535 97.405 ;
        RECT 143.835 97.235 146.215 97.405 ;
        RECT 121.290 96.255 121.460 97.095 ;
        RECT 124.430 96.255 124.600 97.095 ;
        RECT 124.970 96.255 125.140 97.095 ;
        RECT 128.110 96.255 128.280 97.095 ;
        RECT 128.650 96.255 128.820 97.095 ;
        RECT 131.790 96.255 131.960 97.095 ;
        RECT 132.330 96.255 132.500 97.095 ;
        RECT 135.470 96.255 135.640 97.095 ;
        RECT 136.010 96.255 136.180 97.095 ;
        RECT 139.150 96.255 139.320 97.095 ;
        RECT 139.690 96.255 139.860 97.095 ;
        RECT 142.830 96.255 143.000 97.095 ;
        RECT 143.370 96.255 143.540 97.095 ;
        RECT 146.510 96.255 146.680 97.095 ;
        RECT 121.755 95.945 124.135 96.115 ;
        RECT 125.435 95.945 127.815 96.115 ;
        RECT 129.115 95.945 131.495 96.115 ;
        RECT 132.795 95.945 135.175 96.115 ;
        RECT 136.475 95.945 138.855 96.115 ;
        RECT 140.155 95.945 142.535 96.115 ;
        RECT 143.835 95.945 146.215 96.115 ;
        RECT 121.290 94.965 121.460 95.805 ;
        RECT 124.430 94.965 124.600 95.805 ;
        RECT 124.970 94.965 125.140 95.805 ;
        RECT 128.110 94.965 128.280 95.805 ;
        RECT 128.650 94.965 128.820 95.805 ;
        RECT 131.790 94.965 131.960 95.805 ;
        RECT 132.330 94.965 132.500 95.805 ;
        RECT 135.470 94.965 135.640 95.805 ;
        RECT 136.010 94.965 136.180 95.805 ;
        RECT 139.150 94.965 139.320 95.805 ;
        RECT 139.690 94.965 139.860 95.805 ;
        RECT 142.830 94.965 143.000 95.805 ;
        RECT 143.370 94.965 143.540 95.805 ;
        RECT 146.510 94.965 146.680 95.805 ;
        RECT 121.755 94.655 124.135 94.825 ;
        RECT 125.435 94.655 127.815 94.825 ;
        RECT 129.115 94.655 131.495 94.825 ;
        RECT 132.795 94.655 135.175 94.825 ;
        RECT 136.475 94.655 138.855 94.825 ;
        RECT 140.155 94.655 142.535 94.825 ;
        RECT 143.835 94.655 146.215 94.825 ;
        RECT 121.290 93.675 121.460 94.515 ;
        RECT 124.430 93.675 124.600 94.515 ;
        RECT 124.970 93.675 125.140 94.515 ;
        RECT 128.110 93.675 128.280 94.515 ;
        RECT 128.650 93.675 128.820 94.515 ;
        RECT 131.790 93.675 131.960 94.515 ;
        RECT 132.330 93.675 132.500 94.515 ;
        RECT 135.470 93.675 135.640 94.515 ;
        RECT 136.010 93.675 136.180 94.515 ;
        RECT 139.150 93.675 139.320 94.515 ;
        RECT 139.690 93.675 139.860 94.515 ;
        RECT 142.830 93.675 143.000 94.515 ;
        RECT 143.370 93.675 143.540 94.515 ;
        RECT 146.510 93.675 146.680 94.515 ;
        RECT 121.755 93.365 124.135 93.535 ;
        RECT 125.435 93.365 127.815 93.535 ;
        RECT 129.115 93.365 131.495 93.535 ;
        RECT 132.795 93.365 135.175 93.535 ;
        RECT 136.475 93.365 138.855 93.535 ;
        RECT 140.155 93.365 142.535 93.535 ;
        RECT 143.835 93.365 146.215 93.535 ;
        RECT 121.290 92.385 121.460 93.225 ;
        RECT 124.430 92.385 124.600 93.225 ;
        RECT 124.970 92.385 125.140 93.225 ;
        RECT 128.110 92.385 128.280 93.225 ;
        RECT 128.650 92.385 128.820 93.225 ;
        RECT 131.790 92.385 131.960 93.225 ;
        RECT 132.330 92.385 132.500 93.225 ;
        RECT 135.470 92.385 135.640 93.225 ;
        RECT 136.010 92.385 136.180 93.225 ;
        RECT 139.150 92.385 139.320 93.225 ;
        RECT 139.690 92.385 139.860 93.225 ;
        RECT 142.830 92.385 143.000 93.225 ;
        RECT 143.370 92.385 143.540 93.225 ;
        RECT 146.510 92.385 146.680 93.225 ;
        RECT 121.755 92.075 124.135 92.245 ;
        RECT 125.435 92.075 127.815 92.245 ;
        RECT 129.115 92.075 131.495 92.245 ;
        RECT 132.795 92.075 135.175 92.245 ;
        RECT 136.475 92.075 138.855 92.245 ;
        RECT 140.155 92.075 142.535 92.245 ;
        RECT 143.835 92.075 146.215 92.245 ;
        RECT 121.290 91.095 121.460 91.935 ;
        RECT 124.430 91.095 124.600 91.935 ;
        RECT 124.970 91.095 125.140 91.935 ;
        RECT 128.110 91.095 128.280 91.935 ;
        RECT 128.650 91.095 128.820 91.935 ;
        RECT 131.790 91.095 131.960 91.935 ;
        RECT 132.330 91.095 132.500 91.935 ;
        RECT 135.470 91.095 135.640 91.935 ;
        RECT 136.010 91.095 136.180 91.935 ;
        RECT 139.150 91.095 139.320 91.935 ;
        RECT 139.690 91.095 139.860 91.935 ;
        RECT 142.830 91.095 143.000 91.935 ;
        RECT 143.370 91.095 143.540 91.935 ;
        RECT 146.510 91.095 146.680 91.935 ;
        RECT 121.755 90.785 124.135 90.955 ;
        RECT 125.435 90.785 127.815 90.955 ;
        RECT 129.115 90.785 131.495 90.955 ;
        RECT 132.795 90.785 135.175 90.955 ;
        RECT 136.475 90.785 138.855 90.955 ;
        RECT 140.155 90.785 142.535 90.955 ;
        RECT 143.835 90.785 146.215 90.955 ;
        RECT 121.290 89.805 121.460 90.645 ;
        RECT 124.430 89.805 124.600 90.645 ;
        RECT 124.970 89.805 125.140 90.645 ;
        RECT 128.110 89.805 128.280 90.645 ;
        RECT 128.650 89.805 128.820 90.645 ;
        RECT 131.790 89.805 131.960 90.645 ;
        RECT 132.330 89.805 132.500 90.645 ;
        RECT 135.470 89.805 135.640 90.645 ;
        RECT 136.010 89.805 136.180 90.645 ;
        RECT 139.150 89.805 139.320 90.645 ;
        RECT 139.690 89.805 139.860 90.645 ;
        RECT 142.830 89.805 143.000 90.645 ;
        RECT 143.370 89.805 143.540 90.645 ;
        RECT 146.510 89.805 146.680 90.645 ;
        RECT 121.755 89.495 124.135 89.665 ;
        RECT 125.435 89.495 127.815 89.665 ;
        RECT 129.115 89.495 131.495 89.665 ;
        RECT 132.795 89.495 135.175 89.665 ;
        RECT 136.475 89.495 138.855 89.665 ;
        RECT 140.155 89.495 142.535 89.665 ;
        RECT 143.835 89.495 146.215 89.665 ;
        RECT 121.290 88.515 121.460 89.355 ;
        RECT 124.430 88.515 124.600 89.355 ;
        RECT 124.970 88.515 125.140 89.355 ;
        RECT 128.110 88.515 128.280 89.355 ;
        RECT 128.650 88.515 128.820 89.355 ;
        RECT 131.790 88.515 131.960 89.355 ;
        RECT 132.330 88.515 132.500 89.355 ;
        RECT 135.470 88.515 135.640 89.355 ;
        RECT 136.010 88.515 136.180 89.355 ;
        RECT 139.150 88.515 139.320 89.355 ;
        RECT 139.690 88.515 139.860 89.355 ;
        RECT 142.830 88.515 143.000 89.355 ;
        RECT 143.370 88.515 143.540 89.355 ;
        RECT 146.510 88.515 146.680 89.355 ;
        RECT 121.755 88.205 124.135 88.375 ;
        RECT 125.435 88.205 127.815 88.375 ;
        RECT 129.115 88.205 131.495 88.375 ;
        RECT 132.795 88.205 135.175 88.375 ;
        RECT 136.475 88.205 138.855 88.375 ;
        RECT 140.155 88.205 142.535 88.375 ;
        RECT 143.835 88.205 146.215 88.375 ;
        RECT 121.290 87.225 121.460 88.065 ;
        RECT 124.430 87.225 124.600 88.065 ;
        RECT 124.970 87.225 125.140 88.065 ;
        RECT 128.110 87.225 128.280 88.065 ;
        RECT 128.650 87.225 128.820 88.065 ;
        RECT 131.790 87.225 131.960 88.065 ;
        RECT 132.330 87.225 132.500 88.065 ;
        RECT 135.470 87.225 135.640 88.065 ;
        RECT 136.010 87.225 136.180 88.065 ;
        RECT 139.150 87.225 139.320 88.065 ;
        RECT 139.690 87.225 139.860 88.065 ;
        RECT 142.830 87.225 143.000 88.065 ;
        RECT 143.370 87.225 143.540 88.065 ;
        RECT 146.510 87.225 146.680 88.065 ;
        RECT 121.755 86.915 124.135 87.085 ;
        RECT 125.435 86.915 127.815 87.085 ;
        RECT 129.115 86.915 131.495 87.085 ;
        RECT 132.795 86.915 135.175 87.085 ;
        RECT 136.475 86.915 138.855 87.085 ;
        RECT 140.155 86.915 142.535 87.085 ;
        RECT 143.835 86.915 146.215 87.085 ;
        RECT 121.290 85.935 121.460 86.775 ;
        RECT 124.430 85.935 124.600 86.775 ;
        RECT 124.970 85.935 125.140 86.775 ;
        RECT 128.110 85.935 128.280 86.775 ;
        RECT 128.650 85.935 128.820 86.775 ;
        RECT 131.790 85.935 131.960 86.775 ;
        RECT 132.330 85.935 132.500 86.775 ;
        RECT 135.470 85.935 135.640 86.775 ;
        RECT 136.010 85.935 136.180 86.775 ;
        RECT 139.150 85.935 139.320 86.775 ;
        RECT 139.690 85.935 139.860 86.775 ;
        RECT 142.830 85.935 143.000 86.775 ;
        RECT 143.370 85.935 143.540 86.775 ;
        RECT 146.510 85.935 146.680 86.775 ;
        RECT 121.755 85.625 124.135 85.795 ;
        RECT 125.435 85.625 127.815 85.795 ;
        RECT 129.115 85.625 131.495 85.795 ;
        RECT 132.795 85.625 135.175 85.795 ;
        RECT 136.475 85.625 138.855 85.795 ;
        RECT 140.155 85.625 142.535 85.795 ;
        RECT 143.835 85.625 146.215 85.795 ;
        RECT 121.290 84.645 121.460 85.485 ;
        RECT 124.430 84.645 124.600 85.485 ;
        RECT 124.970 84.645 125.140 85.485 ;
        RECT 128.110 84.645 128.280 85.485 ;
        RECT 128.650 84.645 128.820 85.485 ;
        RECT 131.790 84.645 131.960 85.485 ;
        RECT 132.330 84.645 132.500 85.485 ;
        RECT 135.470 84.645 135.640 85.485 ;
        RECT 136.010 84.645 136.180 85.485 ;
        RECT 139.150 84.645 139.320 85.485 ;
        RECT 139.690 84.645 139.860 85.485 ;
        RECT 142.830 84.645 143.000 85.485 ;
        RECT 143.370 84.645 143.540 85.485 ;
        RECT 146.510 84.645 146.680 85.485 ;
        RECT 121.755 84.335 124.135 84.505 ;
        RECT 125.435 84.335 127.815 84.505 ;
        RECT 129.115 84.335 131.495 84.505 ;
        RECT 132.795 84.335 135.175 84.505 ;
        RECT 136.475 84.335 138.855 84.505 ;
        RECT 140.155 84.335 142.535 84.505 ;
        RECT 143.835 84.335 146.215 84.505 ;
        RECT 121.290 83.355 121.460 84.195 ;
        RECT 124.430 83.355 124.600 84.195 ;
        RECT 124.970 83.355 125.140 84.195 ;
        RECT 128.110 83.355 128.280 84.195 ;
        RECT 128.650 83.355 128.820 84.195 ;
        RECT 131.790 83.355 131.960 84.195 ;
        RECT 132.330 83.355 132.500 84.195 ;
        RECT 135.470 83.355 135.640 84.195 ;
        RECT 136.010 83.355 136.180 84.195 ;
        RECT 139.150 83.355 139.320 84.195 ;
        RECT 139.690 83.355 139.860 84.195 ;
        RECT 142.830 83.355 143.000 84.195 ;
        RECT 143.370 83.355 143.540 84.195 ;
        RECT 146.510 83.355 146.680 84.195 ;
        RECT 146.940 83.945 147.310 85.465 ;
        RECT 121.755 83.045 124.135 83.215 ;
        RECT 125.435 83.045 127.815 83.215 ;
        RECT 129.115 83.045 131.495 83.215 ;
        RECT 132.795 83.045 135.175 83.215 ;
        RECT 136.475 83.045 138.855 83.215 ;
        RECT 140.155 83.045 142.535 83.215 ;
        RECT 143.835 83.045 146.215 83.215 ;
        RECT 121.290 82.065 121.460 82.905 ;
        RECT 124.430 82.065 124.600 82.905 ;
        RECT 124.970 82.065 125.140 82.905 ;
        RECT 128.110 82.065 128.280 82.905 ;
        RECT 128.650 82.065 128.820 82.905 ;
        RECT 131.790 82.065 131.960 82.905 ;
        RECT 132.330 82.065 132.500 82.905 ;
        RECT 135.470 82.065 135.640 82.905 ;
        RECT 136.010 82.065 136.180 82.905 ;
        RECT 139.150 82.065 139.320 82.905 ;
        RECT 139.690 82.065 139.860 82.905 ;
        RECT 142.830 82.065 143.000 82.905 ;
        RECT 143.370 82.065 143.540 82.905 ;
        RECT 146.510 82.065 146.680 82.905 ;
        RECT 121.755 81.755 124.135 81.925 ;
        RECT 125.435 81.755 127.815 81.925 ;
        RECT 129.115 81.755 131.495 81.925 ;
        RECT 132.795 81.755 135.175 81.925 ;
        RECT 136.475 81.755 138.855 81.925 ;
        RECT 140.155 81.755 142.535 81.925 ;
        RECT 143.835 81.755 146.215 81.925 ;
        RECT 108.620 61.315 109.500 61.485 ;
        RECT 108.200 59.335 108.370 61.175 ;
        RECT 109.750 59.335 109.920 61.175 ;
        RECT 108.620 59.025 109.500 59.195 ;
        RECT 107.570 56.215 107.950 57.475 ;
        RECT 108.200 57.045 108.370 58.885 ;
        RECT 109.750 57.045 109.920 58.885 ;
        RECT 108.620 56.735 109.500 56.905 ;
        RECT 108.200 54.755 108.370 56.595 ;
        RECT 109.750 54.755 109.920 56.595 ;
        RECT 108.620 54.445 109.500 54.615 ;
        RECT 108.200 52.465 108.370 54.305 ;
        RECT 109.750 52.465 109.920 54.305 ;
        RECT 108.620 52.155 109.500 52.325 ;
        RECT 108.200 50.175 108.370 52.015 ;
        RECT 109.750 50.175 109.920 52.015 ;
        RECT 108.620 49.865 109.500 50.035 ;
        RECT 108.200 47.885 108.370 49.725 ;
        RECT 109.750 47.885 109.920 49.725 ;
        RECT 108.620 47.575 109.500 47.745 ;
        RECT 108.200 45.595 108.370 47.435 ;
        RECT 109.750 45.595 109.920 47.435 ;
        RECT 108.620 45.285 109.500 45.455 ;
        RECT 107.550 42.215 107.950 43.405 ;
        RECT 108.200 43.305 108.370 45.145 ;
        RECT 109.750 43.305 109.920 45.145 ;
        RECT 108.620 42.995 109.500 43.165 ;
        RECT 108.200 41.015 108.370 42.855 ;
        RECT 109.750 41.015 109.920 42.855 ;
        RECT 108.620 40.705 109.500 40.875 ;
        RECT 108.200 38.725 108.370 40.565 ;
        RECT 109.750 38.725 109.920 40.565 ;
        RECT 108.620 38.415 109.500 38.585 ;
        RECT 121.755 77.195 124.135 77.365 ;
        RECT 125.435 77.195 127.815 77.365 ;
        RECT 129.115 77.195 131.495 77.365 ;
        RECT 132.795 77.195 135.175 77.365 ;
        RECT 136.475 77.195 138.855 77.365 ;
        RECT 140.155 77.195 142.535 77.365 ;
        RECT 143.835 77.195 146.215 77.365 ;
        RECT 121.290 76.215 121.460 77.055 ;
        RECT 124.430 76.215 124.600 77.055 ;
        RECT 124.970 76.215 125.140 77.055 ;
        RECT 128.110 76.215 128.280 77.055 ;
        RECT 128.650 76.215 128.820 77.055 ;
        RECT 131.790 76.215 131.960 77.055 ;
        RECT 132.330 76.215 132.500 77.055 ;
        RECT 135.470 76.215 135.640 77.055 ;
        RECT 136.010 76.215 136.180 77.055 ;
        RECT 139.150 76.215 139.320 77.055 ;
        RECT 139.690 76.215 139.860 77.055 ;
        RECT 142.830 76.215 143.000 77.055 ;
        RECT 143.370 76.215 143.540 77.055 ;
        RECT 146.510 76.215 146.680 77.055 ;
        RECT 121.755 75.905 124.135 76.075 ;
        RECT 125.435 75.905 127.815 76.075 ;
        RECT 129.115 75.905 131.495 76.075 ;
        RECT 132.795 75.905 135.175 76.075 ;
        RECT 136.475 75.905 138.855 76.075 ;
        RECT 140.155 75.905 142.535 76.075 ;
        RECT 143.835 75.905 146.215 76.075 ;
        RECT 121.290 74.925 121.460 75.765 ;
        RECT 124.430 74.925 124.600 75.765 ;
        RECT 124.970 74.925 125.140 75.765 ;
        RECT 128.110 74.925 128.280 75.765 ;
        RECT 128.650 74.925 128.820 75.765 ;
        RECT 131.790 74.925 131.960 75.765 ;
        RECT 132.330 74.925 132.500 75.765 ;
        RECT 135.470 74.925 135.640 75.765 ;
        RECT 136.010 74.925 136.180 75.765 ;
        RECT 139.150 74.925 139.320 75.765 ;
        RECT 139.690 74.925 139.860 75.765 ;
        RECT 142.830 74.925 143.000 75.765 ;
        RECT 143.370 74.925 143.540 75.765 ;
        RECT 146.510 74.925 146.680 75.765 ;
        RECT 121.755 74.615 124.135 74.785 ;
        RECT 125.435 74.615 127.815 74.785 ;
        RECT 129.115 74.615 131.495 74.785 ;
        RECT 132.795 74.615 135.175 74.785 ;
        RECT 136.475 74.615 138.855 74.785 ;
        RECT 140.155 74.615 142.535 74.785 ;
        RECT 143.835 74.615 146.215 74.785 ;
        RECT 121.290 73.635 121.460 74.475 ;
        RECT 124.430 73.635 124.600 74.475 ;
        RECT 124.970 73.635 125.140 74.475 ;
        RECT 128.110 73.635 128.280 74.475 ;
        RECT 128.650 73.635 128.820 74.475 ;
        RECT 131.790 73.635 131.960 74.475 ;
        RECT 132.330 73.635 132.500 74.475 ;
        RECT 135.470 73.635 135.640 74.475 ;
        RECT 136.010 73.635 136.180 74.475 ;
        RECT 139.150 73.635 139.320 74.475 ;
        RECT 139.690 73.635 139.860 74.475 ;
        RECT 142.830 73.635 143.000 74.475 ;
        RECT 143.370 73.635 143.540 74.475 ;
        RECT 146.950 74.485 147.300 75.925 ;
        RECT 146.510 73.635 146.680 74.475 ;
        RECT 121.755 73.325 124.135 73.495 ;
        RECT 125.435 73.325 127.815 73.495 ;
        RECT 129.115 73.325 131.495 73.495 ;
        RECT 132.795 73.325 135.175 73.495 ;
        RECT 136.475 73.325 138.855 73.495 ;
        RECT 140.155 73.325 142.535 73.495 ;
        RECT 143.835 73.325 146.215 73.495 ;
        RECT 121.290 72.345 121.460 73.185 ;
        RECT 124.430 72.345 124.600 73.185 ;
        RECT 124.970 72.345 125.140 73.185 ;
        RECT 128.110 72.345 128.280 73.185 ;
        RECT 128.650 72.345 128.820 73.185 ;
        RECT 131.790 72.345 131.960 73.185 ;
        RECT 132.330 72.345 132.500 73.185 ;
        RECT 135.470 72.345 135.640 73.185 ;
        RECT 136.010 72.345 136.180 73.185 ;
        RECT 139.150 72.345 139.320 73.185 ;
        RECT 139.690 72.345 139.860 73.185 ;
        RECT 142.830 72.345 143.000 73.185 ;
        RECT 143.370 72.345 143.540 73.185 ;
        RECT 146.510 72.345 146.680 73.185 ;
        RECT 121.755 72.035 124.135 72.205 ;
        RECT 125.435 72.035 127.815 72.205 ;
        RECT 129.115 72.035 131.495 72.205 ;
        RECT 132.795 72.035 135.175 72.205 ;
        RECT 136.475 72.035 138.855 72.205 ;
        RECT 140.155 72.035 142.535 72.205 ;
        RECT 143.835 72.035 146.215 72.205 ;
        RECT 121.290 71.055 121.460 71.895 ;
        RECT 124.430 71.055 124.600 71.895 ;
        RECT 124.970 71.055 125.140 71.895 ;
        RECT 128.110 71.055 128.280 71.895 ;
        RECT 128.650 71.055 128.820 71.895 ;
        RECT 131.790 71.055 131.960 71.895 ;
        RECT 132.330 71.055 132.500 71.895 ;
        RECT 135.470 71.055 135.640 71.895 ;
        RECT 136.010 71.055 136.180 71.895 ;
        RECT 139.150 71.055 139.320 71.895 ;
        RECT 139.690 71.055 139.860 71.895 ;
        RECT 142.830 71.055 143.000 71.895 ;
        RECT 143.370 71.055 143.540 71.895 ;
        RECT 146.510 71.055 146.680 71.895 ;
        RECT 121.755 70.745 124.135 70.915 ;
        RECT 125.435 70.745 127.815 70.915 ;
        RECT 129.115 70.745 131.495 70.915 ;
        RECT 132.795 70.745 135.175 70.915 ;
        RECT 136.475 70.745 138.855 70.915 ;
        RECT 140.155 70.745 142.535 70.915 ;
        RECT 143.835 70.745 146.215 70.915 ;
        RECT 121.290 69.765 121.460 70.605 ;
        RECT 124.430 69.765 124.600 70.605 ;
        RECT 124.970 69.765 125.140 70.605 ;
        RECT 128.110 69.765 128.280 70.605 ;
        RECT 128.650 69.765 128.820 70.605 ;
        RECT 131.790 69.765 131.960 70.605 ;
        RECT 132.330 69.765 132.500 70.605 ;
        RECT 135.470 69.765 135.640 70.605 ;
        RECT 136.010 69.765 136.180 70.605 ;
        RECT 139.150 69.765 139.320 70.605 ;
        RECT 139.690 69.765 139.860 70.605 ;
        RECT 142.830 69.765 143.000 70.605 ;
        RECT 143.370 69.765 143.540 70.605 ;
        RECT 146.510 69.765 146.680 70.605 ;
        RECT 121.755 69.455 124.135 69.625 ;
        RECT 125.435 69.455 127.815 69.625 ;
        RECT 129.115 69.455 131.495 69.625 ;
        RECT 132.795 69.455 135.175 69.625 ;
        RECT 136.475 69.455 138.855 69.625 ;
        RECT 140.155 69.455 142.535 69.625 ;
        RECT 143.835 69.455 146.215 69.625 ;
        RECT 121.290 68.475 121.460 69.315 ;
        RECT 124.430 68.475 124.600 69.315 ;
        RECT 124.970 68.475 125.140 69.315 ;
        RECT 128.110 68.475 128.280 69.315 ;
        RECT 128.650 68.475 128.820 69.315 ;
        RECT 131.790 68.475 131.960 69.315 ;
        RECT 132.330 68.475 132.500 69.315 ;
        RECT 135.470 68.475 135.640 69.315 ;
        RECT 136.010 68.475 136.180 69.315 ;
        RECT 139.150 68.475 139.320 69.315 ;
        RECT 139.690 68.475 139.860 69.315 ;
        RECT 142.830 68.475 143.000 69.315 ;
        RECT 143.370 68.475 143.540 69.315 ;
        RECT 146.510 68.475 146.680 69.315 ;
        RECT 121.755 68.165 124.135 68.335 ;
        RECT 125.435 68.165 127.815 68.335 ;
        RECT 129.115 68.165 131.495 68.335 ;
        RECT 132.795 68.165 135.175 68.335 ;
        RECT 136.475 68.165 138.855 68.335 ;
        RECT 140.155 68.165 142.535 68.335 ;
        RECT 143.835 68.165 146.215 68.335 ;
        RECT 121.290 67.185 121.460 68.025 ;
        RECT 124.430 67.185 124.600 68.025 ;
        RECT 124.970 67.185 125.140 68.025 ;
        RECT 128.110 67.185 128.280 68.025 ;
        RECT 128.650 67.185 128.820 68.025 ;
        RECT 131.790 67.185 131.960 68.025 ;
        RECT 132.330 67.185 132.500 68.025 ;
        RECT 135.470 67.185 135.640 68.025 ;
        RECT 136.010 67.185 136.180 68.025 ;
        RECT 139.150 67.185 139.320 68.025 ;
        RECT 139.690 67.185 139.860 68.025 ;
        RECT 142.830 67.185 143.000 68.025 ;
        RECT 143.370 67.185 143.540 68.025 ;
        RECT 146.510 67.185 146.680 68.025 ;
        RECT 121.755 66.875 124.135 67.045 ;
        RECT 125.435 66.875 127.815 67.045 ;
        RECT 129.115 66.875 131.495 67.045 ;
        RECT 132.795 66.875 135.175 67.045 ;
        RECT 136.475 66.875 138.855 67.045 ;
        RECT 140.155 66.875 142.535 67.045 ;
        RECT 143.835 66.875 146.215 67.045 ;
        RECT 121.290 65.895 121.460 66.735 ;
        RECT 124.430 65.895 124.600 66.735 ;
        RECT 124.970 65.895 125.140 66.735 ;
        RECT 128.110 65.895 128.280 66.735 ;
        RECT 128.650 65.895 128.820 66.735 ;
        RECT 131.790 65.895 131.960 66.735 ;
        RECT 132.330 65.895 132.500 66.735 ;
        RECT 135.470 65.895 135.640 66.735 ;
        RECT 136.010 65.895 136.180 66.735 ;
        RECT 139.150 65.895 139.320 66.735 ;
        RECT 139.690 65.895 139.860 66.735 ;
        RECT 142.830 65.895 143.000 66.735 ;
        RECT 143.370 65.895 143.540 66.735 ;
        RECT 146.510 65.895 146.680 66.735 ;
        RECT 121.755 65.585 124.135 65.755 ;
        RECT 125.435 65.585 127.815 65.755 ;
        RECT 129.115 65.585 131.495 65.755 ;
        RECT 132.795 65.585 135.175 65.755 ;
        RECT 136.475 65.585 138.855 65.755 ;
        RECT 140.155 65.585 142.535 65.755 ;
        RECT 143.835 65.585 146.215 65.755 ;
        RECT 121.290 64.605 121.460 65.445 ;
        RECT 124.430 64.605 124.600 65.445 ;
        RECT 124.970 64.605 125.140 65.445 ;
        RECT 128.110 64.605 128.280 65.445 ;
        RECT 128.650 64.605 128.820 65.445 ;
        RECT 131.790 64.605 131.960 65.445 ;
        RECT 132.330 64.605 132.500 65.445 ;
        RECT 135.470 64.605 135.640 65.445 ;
        RECT 136.010 64.605 136.180 65.445 ;
        RECT 139.150 64.605 139.320 65.445 ;
        RECT 139.690 64.605 139.860 65.445 ;
        RECT 142.830 64.605 143.000 65.445 ;
        RECT 143.370 64.605 143.540 65.445 ;
        RECT 146.510 64.605 146.680 65.445 ;
        RECT 121.755 64.295 124.135 64.465 ;
        RECT 125.435 64.295 127.815 64.465 ;
        RECT 129.115 64.295 131.495 64.465 ;
        RECT 132.795 64.295 135.175 64.465 ;
        RECT 136.475 64.295 138.855 64.465 ;
        RECT 140.155 64.295 142.535 64.465 ;
        RECT 143.835 64.295 146.215 64.465 ;
        RECT 121.290 63.315 121.460 64.155 ;
        RECT 124.430 63.315 124.600 64.155 ;
        RECT 124.970 63.315 125.140 64.155 ;
        RECT 128.110 63.315 128.280 64.155 ;
        RECT 128.650 63.315 128.820 64.155 ;
        RECT 131.790 63.315 131.960 64.155 ;
        RECT 132.330 63.315 132.500 64.155 ;
        RECT 135.470 63.315 135.640 64.155 ;
        RECT 136.010 63.315 136.180 64.155 ;
        RECT 139.150 63.315 139.320 64.155 ;
        RECT 139.690 63.315 139.860 64.155 ;
        RECT 142.830 63.315 143.000 64.155 ;
        RECT 143.370 63.315 143.540 64.155 ;
        RECT 146.510 63.315 146.680 64.155 ;
        RECT 121.755 63.005 124.135 63.175 ;
        RECT 125.435 63.005 127.815 63.175 ;
        RECT 129.115 63.005 131.495 63.175 ;
        RECT 132.795 63.005 135.175 63.175 ;
        RECT 136.475 63.005 138.855 63.175 ;
        RECT 140.155 63.005 142.535 63.175 ;
        RECT 143.835 63.005 146.215 63.175 ;
        RECT 121.290 62.025 121.460 62.865 ;
        RECT 124.430 62.025 124.600 62.865 ;
        RECT 124.970 62.025 125.140 62.865 ;
        RECT 128.110 62.025 128.280 62.865 ;
        RECT 128.650 62.025 128.820 62.865 ;
        RECT 131.790 62.025 131.960 62.865 ;
        RECT 132.330 62.025 132.500 62.865 ;
        RECT 135.470 62.025 135.640 62.865 ;
        RECT 136.010 62.025 136.180 62.865 ;
        RECT 139.150 62.025 139.320 62.865 ;
        RECT 139.690 62.025 139.860 62.865 ;
        RECT 142.830 62.025 143.000 62.865 ;
        RECT 143.370 62.025 143.540 62.865 ;
        RECT 146.510 62.025 146.680 62.865 ;
        RECT 121.755 61.715 124.135 61.885 ;
        RECT 125.435 61.715 127.815 61.885 ;
        RECT 129.115 61.715 131.495 61.885 ;
        RECT 132.795 61.715 135.175 61.885 ;
        RECT 136.475 61.715 138.855 61.885 ;
        RECT 140.155 61.715 142.535 61.885 ;
        RECT 143.835 61.715 146.215 61.885 ;
        RECT 121.290 60.735 121.460 61.575 ;
        RECT 124.430 60.735 124.600 61.575 ;
        RECT 124.970 60.735 125.140 61.575 ;
        RECT 128.110 60.735 128.280 61.575 ;
        RECT 128.650 60.735 128.820 61.575 ;
        RECT 131.790 60.735 131.960 61.575 ;
        RECT 132.330 60.735 132.500 61.575 ;
        RECT 135.470 60.735 135.640 61.575 ;
        RECT 136.010 60.735 136.180 61.575 ;
        RECT 139.150 60.735 139.320 61.575 ;
        RECT 139.690 60.735 139.860 61.575 ;
        RECT 142.830 60.735 143.000 61.575 ;
        RECT 143.370 60.735 143.540 61.575 ;
        RECT 146.510 60.735 146.680 61.575 ;
        RECT 121.755 60.425 124.135 60.595 ;
        RECT 125.435 60.425 127.815 60.595 ;
        RECT 129.115 60.425 131.495 60.595 ;
        RECT 132.795 60.425 135.175 60.595 ;
        RECT 136.475 60.425 138.855 60.595 ;
        RECT 140.155 60.425 142.535 60.595 ;
        RECT 143.835 60.425 146.215 60.595 ;
        RECT 121.290 59.445 121.460 60.285 ;
        RECT 124.430 59.445 124.600 60.285 ;
        RECT 124.970 59.445 125.140 60.285 ;
        RECT 128.110 59.445 128.280 60.285 ;
        RECT 128.650 59.445 128.820 60.285 ;
        RECT 131.790 59.445 131.960 60.285 ;
        RECT 132.330 59.445 132.500 60.285 ;
        RECT 135.470 59.445 135.640 60.285 ;
        RECT 136.010 59.445 136.180 60.285 ;
        RECT 139.150 59.445 139.320 60.285 ;
        RECT 139.690 59.445 139.860 60.285 ;
        RECT 142.830 59.445 143.000 60.285 ;
        RECT 143.370 59.445 143.540 60.285 ;
        RECT 146.510 59.445 146.680 60.285 ;
        RECT 121.755 59.135 124.135 59.305 ;
        RECT 125.435 59.135 127.815 59.305 ;
        RECT 129.115 59.135 131.495 59.305 ;
        RECT 132.795 59.135 135.175 59.305 ;
        RECT 136.475 59.135 138.855 59.305 ;
        RECT 140.155 59.135 142.535 59.305 ;
        RECT 143.835 59.135 146.215 59.305 ;
        RECT 121.290 58.155 121.460 58.995 ;
        RECT 124.430 58.155 124.600 58.995 ;
        RECT 124.970 58.155 125.140 58.995 ;
        RECT 128.110 58.155 128.280 58.995 ;
        RECT 128.650 58.155 128.820 58.995 ;
        RECT 131.790 58.155 131.960 58.995 ;
        RECT 132.330 58.155 132.500 58.995 ;
        RECT 135.470 58.155 135.640 58.995 ;
        RECT 136.010 58.155 136.180 58.995 ;
        RECT 139.150 58.155 139.320 58.995 ;
        RECT 139.690 58.155 139.860 58.995 ;
        RECT 142.830 58.155 143.000 58.995 ;
        RECT 143.370 58.155 143.540 58.995 ;
        RECT 146.510 58.155 146.680 58.995 ;
        RECT 121.755 57.845 124.135 58.015 ;
        RECT 125.435 57.845 127.815 58.015 ;
        RECT 129.115 57.845 131.495 58.015 ;
        RECT 132.795 57.845 135.175 58.015 ;
        RECT 136.475 57.845 138.855 58.015 ;
        RECT 140.155 57.845 142.535 58.015 ;
        RECT 143.835 57.845 146.215 58.015 ;
        RECT 121.290 56.865 121.460 57.705 ;
        RECT 124.430 56.865 124.600 57.705 ;
        RECT 124.970 56.865 125.140 57.705 ;
        RECT 128.110 56.865 128.280 57.705 ;
        RECT 128.650 56.865 128.820 57.705 ;
        RECT 131.790 56.865 131.960 57.705 ;
        RECT 132.330 56.865 132.500 57.705 ;
        RECT 135.470 56.865 135.640 57.705 ;
        RECT 136.010 56.865 136.180 57.705 ;
        RECT 139.150 56.865 139.320 57.705 ;
        RECT 139.690 56.865 139.860 57.705 ;
        RECT 142.830 56.865 143.000 57.705 ;
        RECT 143.370 56.865 143.540 57.705 ;
        RECT 146.510 56.865 146.680 57.705 ;
        RECT 121.755 56.555 124.135 56.725 ;
        RECT 125.435 56.555 127.815 56.725 ;
        RECT 129.115 56.555 131.495 56.725 ;
        RECT 132.795 56.555 135.175 56.725 ;
        RECT 136.475 56.555 138.855 56.725 ;
        RECT 140.155 56.555 142.535 56.725 ;
        RECT 143.835 56.555 146.215 56.725 ;
        RECT 121.290 55.575 121.460 56.415 ;
        RECT 124.430 55.575 124.600 56.415 ;
        RECT 124.970 55.575 125.140 56.415 ;
        RECT 128.110 55.575 128.280 56.415 ;
        RECT 128.650 55.575 128.820 56.415 ;
        RECT 131.790 55.575 131.960 56.415 ;
        RECT 132.330 55.575 132.500 56.415 ;
        RECT 135.470 55.575 135.640 56.415 ;
        RECT 136.010 55.575 136.180 56.415 ;
        RECT 139.150 55.575 139.320 56.415 ;
        RECT 139.690 55.575 139.860 56.415 ;
        RECT 142.830 55.575 143.000 56.415 ;
        RECT 143.370 55.575 143.540 56.415 ;
        RECT 146.510 55.575 146.680 56.415 ;
        RECT 121.755 55.265 124.135 55.435 ;
        RECT 125.435 55.265 127.815 55.435 ;
        RECT 129.115 55.265 131.495 55.435 ;
        RECT 132.795 55.265 135.175 55.435 ;
        RECT 136.475 55.265 138.855 55.435 ;
        RECT 140.155 55.265 142.535 55.435 ;
        RECT 143.835 55.265 146.215 55.435 ;
        RECT 121.290 54.285 121.460 55.125 ;
        RECT 124.430 54.285 124.600 55.125 ;
        RECT 124.970 54.285 125.140 55.125 ;
        RECT 128.110 54.285 128.280 55.125 ;
        RECT 128.650 54.285 128.820 55.125 ;
        RECT 131.790 54.285 131.960 55.125 ;
        RECT 132.330 54.285 132.500 55.125 ;
        RECT 135.470 54.285 135.640 55.125 ;
        RECT 136.010 54.285 136.180 55.125 ;
        RECT 139.150 54.285 139.320 55.125 ;
        RECT 139.690 54.285 139.860 55.125 ;
        RECT 142.830 54.285 143.000 55.125 ;
        RECT 143.370 54.285 143.540 55.125 ;
        RECT 146.510 54.285 146.680 55.125 ;
        RECT 121.755 53.975 124.135 54.145 ;
        RECT 125.435 53.975 127.815 54.145 ;
        RECT 129.115 53.975 131.495 54.145 ;
        RECT 132.795 53.975 135.175 54.145 ;
        RECT 136.475 53.975 138.855 54.145 ;
        RECT 140.155 53.975 142.535 54.145 ;
        RECT 143.835 53.975 146.215 54.145 ;
        RECT 121.290 52.995 121.460 53.835 ;
        RECT 124.430 52.995 124.600 53.835 ;
        RECT 124.970 52.995 125.140 53.835 ;
        RECT 128.110 52.995 128.280 53.835 ;
        RECT 128.650 52.995 128.820 53.835 ;
        RECT 131.790 52.995 131.960 53.835 ;
        RECT 132.330 52.995 132.500 53.835 ;
        RECT 135.470 52.995 135.640 53.835 ;
        RECT 136.010 52.995 136.180 53.835 ;
        RECT 139.150 52.995 139.320 53.835 ;
        RECT 139.690 52.995 139.860 53.835 ;
        RECT 142.830 52.995 143.000 53.835 ;
        RECT 143.370 52.995 143.540 53.835 ;
        RECT 146.510 52.995 146.680 53.835 ;
        RECT 146.930 53.695 147.310 55.155 ;
        RECT 121.755 52.685 124.135 52.855 ;
        RECT 125.435 52.685 127.815 52.855 ;
        RECT 129.115 52.685 131.495 52.855 ;
        RECT 132.795 52.685 135.175 52.855 ;
        RECT 136.475 52.685 138.855 52.855 ;
        RECT 140.155 52.685 142.535 52.855 ;
        RECT 143.835 52.685 146.215 52.855 ;
        RECT 121.290 51.705 121.460 52.545 ;
        RECT 124.430 51.705 124.600 52.545 ;
        RECT 124.970 51.705 125.140 52.545 ;
        RECT 128.110 51.705 128.280 52.545 ;
        RECT 128.650 51.705 128.820 52.545 ;
        RECT 131.790 51.705 131.960 52.545 ;
        RECT 132.330 51.705 132.500 52.545 ;
        RECT 135.470 51.705 135.640 52.545 ;
        RECT 136.010 51.705 136.180 52.545 ;
        RECT 139.150 51.705 139.320 52.545 ;
        RECT 139.690 51.705 139.860 52.545 ;
        RECT 142.830 51.705 143.000 52.545 ;
        RECT 143.370 51.705 143.540 52.545 ;
        RECT 146.510 51.705 146.680 52.545 ;
        RECT 121.755 51.395 124.135 51.565 ;
        RECT 125.435 51.395 127.815 51.565 ;
        RECT 129.115 51.395 131.495 51.565 ;
        RECT 132.795 51.395 135.175 51.565 ;
        RECT 136.475 51.395 138.855 51.565 ;
        RECT 140.155 51.395 142.535 51.565 ;
        RECT 143.835 51.395 146.215 51.565 ;
        RECT 113.730 43.615 114.610 43.785 ;
        RECT 112.700 39.785 113.000 43.035 ;
        RECT 113.310 41.635 113.480 43.475 ;
        RECT 114.860 41.635 115.030 43.475 ;
        RECT 113.730 41.325 114.610 41.495 ;
        RECT 113.310 39.345 113.480 41.185 ;
        RECT 114.860 39.345 115.030 41.185 ;
        RECT 113.730 39.035 114.610 39.205 ;
        RECT 118.770 43.795 122.650 43.965 ;
        RECT 123.860 43.795 127.740 43.965 ;
        RECT 118.350 43.555 118.520 43.725 ;
        RECT 127.990 43.555 128.160 43.725 ;
        RECT 117.780 39.605 118.030 43.435 ;
        RECT 118.770 43.315 122.650 43.485 ;
        RECT 122.900 43.075 123.070 43.245 ;
        RECT 118.770 42.835 122.650 43.005 ;
        RECT 123.860 43.315 127.740 43.485 ;
        RECT 123.440 43.075 123.610 43.245 ;
        RECT 123.860 42.835 127.740 43.005 ;
        RECT 118.350 42.595 118.520 42.765 ;
        RECT 127.990 42.595 128.160 42.765 ;
        RECT 118.770 42.355 122.650 42.525 ;
        RECT 122.900 42.115 123.070 42.285 ;
        RECT 118.770 41.875 122.650 42.045 ;
        RECT 123.860 42.355 127.740 42.525 ;
        RECT 123.440 42.115 123.610 42.285 ;
        RECT 123.860 41.875 127.740 42.045 ;
        RECT 118.350 41.635 118.520 41.805 ;
        RECT 127.990 41.635 128.160 41.805 ;
        RECT 118.770 41.395 122.650 41.565 ;
        RECT 122.900 41.155 123.070 41.325 ;
        RECT 118.770 40.915 122.650 41.085 ;
        RECT 123.860 41.395 127.740 41.565 ;
        RECT 123.440 41.155 123.610 41.325 ;
        RECT 123.860 40.915 127.740 41.085 ;
        RECT 118.350 40.675 118.520 40.845 ;
        RECT 127.990 40.675 128.160 40.845 ;
        RECT 118.770 40.435 122.650 40.605 ;
        RECT 122.900 40.195 123.070 40.365 ;
        RECT 118.770 39.955 122.650 40.125 ;
        RECT 123.860 40.435 127.740 40.605 ;
        RECT 123.440 40.195 123.610 40.365 ;
        RECT 123.860 39.955 127.740 40.125 ;
        RECT 118.350 39.715 118.520 39.885 ;
        RECT 127.990 39.715 128.160 39.885 ;
        RECT 118.770 39.475 122.650 39.645 ;
        RECT 122.900 39.235 123.070 39.405 ;
        RECT 118.770 38.995 122.650 39.165 ;
        RECT 123.860 39.475 127.740 39.645 ;
        RECT 123.440 39.235 123.610 39.405 ;
        RECT 123.860 38.995 127.740 39.165 ;
        RECT 131.655 43.735 136.535 43.905 ;
        RECT 131.190 43.495 131.360 43.665 ;
        RECT 131.655 43.255 136.535 43.425 ;
        RECT 136.830 43.015 137.000 43.185 ;
        RECT 131.655 42.775 136.535 42.945 ;
        RECT 141.055 45.825 145.935 45.995 ;
        RECT 140.590 44.845 140.760 45.685 ;
        RECT 146.230 44.845 146.400 45.685 ;
        RECT 146.660 44.795 147.040 45.665 ;
        RECT 141.055 44.535 145.935 44.705 ;
        RECT 131.190 42.535 131.360 42.705 ;
        RECT 131.655 42.295 136.535 42.465 ;
        RECT 136.830 42.055 137.000 42.225 ;
        RECT 131.655 41.815 136.535 41.985 ;
        RECT 131.190 41.575 131.360 41.745 ;
        RECT 131.655 41.335 136.535 41.505 ;
        RECT 136.830 41.095 137.000 41.265 ;
        RECT 131.655 40.855 136.535 41.025 ;
        RECT 131.190 40.615 131.360 40.785 ;
        RECT 131.655 40.375 136.535 40.545 ;
        RECT 136.830 40.135 137.000 40.305 ;
        RECT 131.655 39.895 136.535 40.065 ;
        RECT 137.300 40.115 137.610 42.815 ;
        RECT 131.190 39.655 131.360 39.825 ;
        RECT 131.655 39.415 136.535 39.585 ;
        RECT 136.830 39.175 137.000 39.345 ;
        RECT 131.655 38.935 136.535 39.105 ;
        RECT 141.045 40.365 145.925 40.535 ;
        RECT 140.580 39.385 140.750 40.225 ;
        RECT 146.220 39.385 146.390 40.225 ;
        RECT 146.670 39.395 147.050 40.205 ;
        RECT 141.045 39.075 145.925 39.245 ;
      LAYER met1 ;
        RECT 102.730 146.985 105.075 162.755 ;
        RECT 118.135 147.805 119.085 148.695 ;
        RECT 138.725 148.600 139.590 148.605 ;
        RECT 102.680 146.790 105.075 146.985 ;
        RECT 102.680 145.240 115.180 146.790 ;
        RECT 118.165 146.545 119.055 147.805 ;
        RECT 138.700 147.745 139.615 148.600 ;
        RECT 118.165 145.555 119.200 146.545 ;
        RECT 138.725 146.525 139.590 147.745 ;
        RECT 149.000 146.885 151.200 162.960 ;
        RECT 118.200 145.545 119.200 145.555 ;
        RECT 102.680 144.160 104.910 145.240 ;
        RECT 113.630 144.160 115.180 145.240 ;
        RECT 118.265 144.660 119.060 145.545 ;
        RECT 102.680 142.885 104.920 144.160 ;
        RECT 108.170 143.135 109.995 143.145 ;
        RECT 110.590 143.135 111.915 143.305 ;
        RECT 113.620 143.195 115.180 144.160 ;
        RECT 118.205 143.810 119.115 144.660 ;
        RECT 131.955 144.305 132.985 144.335 ;
        RECT 108.170 142.895 111.915 143.135 ;
        RECT 102.680 137.175 104.910 142.885 ;
        RECT 102.680 135.485 108.010 137.175 ;
        RECT 102.680 123.225 104.910 135.485 ;
        RECT 102.680 121.545 108.010 123.225 ;
        RECT 102.680 116.350 104.910 121.545 ;
        RECT 108.170 118.045 108.420 142.895 ;
        RECT 109.710 142.845 111.915 142.895 ;
        RECT 108.580 141.015 108.860 141.135 ;
        RECT 108.560 140.785 109.560 141.015 ;
        RECT 108.580 140.685 108.860 140.785 ;
        RECT 109.710 138.775 110.000 142.845 ;
        RECT 110.590 142.670 111.915 142.845 ;
        RECT 113.630 142.965 115.180 143.195 ;
        RECT 122.930 143.275 132.985 144.305 ;
        RECT 113.630 142.545 122.340 142.965 ;
        RECT 113.630 141.295 115.180 142.545 ;
        RECT 114.570 141.015 114.880 141.085 ;
        RECT 109.130 138.725 110.000 138.775 ;
        RECT 108.560 138.495 110.000 138.725 ;
        RECT 109.130 138.435 110.000 138.495 ;
        RECT 108.590 136.435 108.870 136.545 ;
        RECT 108.560 136.205 109.560 136.435 ;
        RECT 108.590 136.095 108.870 136.205 ;
        RECT 109.710 134.215 110.000 138.435 ;
        RECT 109.130 134.145 110.000 134.215 ;
        RECT 108.560 133.915 110.000 134.145 ;
        RECT 109.130 133.875 110.000 133.915 ;
        RECT 108.590 131.855 108.870 131.975 ;
        RECT 108.560 131.625 109.560 131.855 ;
        RECT 108.590 131.525 108.870 131.625 ;
        RECT 109.710 129.615 110.000 133.875 ;
        RECT 109.130 129.565 110.000 129.615 ;
        RECT 108.560 129.335 110.000 129.565 ;
        RECT 109.130 129.275 110.000 129.335 ;
        RECT 108.590 127.275 108.870 127.385 ;
        RECT 108.560 127.045 109.560 127.275 ;
        RECT 108.590 126.935 108.870 127.045 ;
        RECT 109.710 125.045 110.000 129.275 ;
        RECT 109.130 124.985 110.000 125.045 ;
        RECT 108.560 124.755 110.000 124.985 ;
        RECT 109.130 124.705 110.000 124.755 ;
        RECT 108.590 122.695 108.870 122.815 ;
        RECT 108.560 122.465 109.560 122.695 ;
        RECT 108.590 122.365 108.870 122.465 ;
        RECT 109.710 120.465 110.000 124.705 ;
        RECT 109.130 120.405 110.000 120.465 ;
        RECT 108.560 120.175 110.000 120.405 ;
        RECT 109.130 120.125 110.000 120.175 ;
        RECT 108.590 118.115 108.870 118.215 ;
        RECT 108.560 117.885 109.560 118.115 ;
        RECT 109.710 118.035 110.000 120.125 ;
        RECT 113.310 140.735 113.680 140.925 ;
        RECT 113.870 140.785 114.880 141.015 ;
        RECT 113.310 138.775 113.710 140.735 ;
        RECT 114.570 140.705 114.880 140.785 ;
        RECT 115.050 140.735 115.420 140.945 ;
        RECT 113.310 138.445 113.680 138.775 ;
        RECT 113.860 138.725 114.140 138.825 ;
        RECT 115.030 138.775 115.420 140.735 ;
        RECT 113.860 138.495 114.870 138.725 ;
        RECT 113.310 136.485 113.710 138.445 ;
        RECT 113.860 138.375 114.140 138.495 ;
        RECT 115.050 138.445 115.420 138.775 ;
        RECT 116.505 138.625 117.310 139.370 ;
        RECT 113.310 136.155 113.680 136.485 ;
        RECT 114.570 136.435 114.880 136.505 ;
        RECT 115.030 136.485 115.420 138.445 ;
        RECT 113.870 136.205 114.880 136.435 ;
        RECT 113.310 134.195 113.710 136.155 ;
        RECT 114.570 136.125 114.880 136.205 ;
        RECT 115.050 136.155 115.420 136.485 ;
        RECT 113.310 133.865 113.680 134.195 ;
        RECT 113.860 134.145 114.140 134.245 ;
        RECT 115.030 134.195 115.420 136.155 ;
        RECT 113.860 133.915 114.870 134.145 ;
        RECT 113.310 131.905 113.710 133.865 ;
        RECT 113.860 133.795 114.140 133.915 ;
        RECT 115.050 133.865 115.420 134.195 ;
        RECT 113.310 131.575 113.680 131.905 ;
        RECT 114.570 131.855 114.880 131.925 ;
        RECT 115.030 131.905 115.420 133.865 ;
        RECT 113.870 131.625 114.880 131.855 ;
        RECT 113.310 129.615 113.710 131.575 ;
        RECT 114.570 131.545 114.880 131.625 ;
        RECT 115.050 131.575 115.420 131.905 ;
        RECT 113.310 129.285 113.680 129.615 ;
        RECT 113.870 129.565 114.150 129.675 ;
        RECT 115.030 129.615 115.420 131.575 ;
        RECT 113.870 129.335 114.870 129.565 ;
        RECT 113.310 127.325 113.710 129.285 ;
        RECT 113.870 129.225 114.150 129.335 ;
        RECT 115.050 129.285 115.420 129.615 ;
        RECT 113.310 126.995 113.680 127.325 ;
        RECT 114.570 127.275 114.880 127.345 ;
        RECT 115.030 127.325 115.420 129.285 ;
        RECT 116.535 129.895 117.280 138.625 ;
        RECT 121.920 130.825 122.340 142.545 ;
        RECT 122.930 141.485 123.960 143.275 ;
        RECT 131.955 143.245 132.985 143.275 ;
        RECT 122.930 141.355 124.960 141.485 ;
        RECT 122.720 141.105 124.960 141.355 ;
        RECT 122.930 140.945 124.960 141.105 ;
        RECT 132.640 140.925 134.950 141.395 ;
        RECT 122.610 139.005 124.910 139.525 ;
        RECT 134.450 139.485 134.950 140.925 ;
        RECT 122.610 137.645 123.130 139.005 ;
        RECT 132.670 138.985 134.950 139.485 ;
        RECT 122.610 137.125 124.890 137.645 ;
        RECT 132.620 137.125 134.980 137.675 ;
        RECT 122.590 135.015 124.910 135.585 ;
        RECT 134.430 135.570 134.980 137.125 ;
        RECT 134.430 135.020 136.975 135.570 ;
        RECT 122.590 133.590 123.160 135.015 ;
        RECT 122.590 133.020 125.015 133.590 ;
        RECT 134.630 133.035 136.990 133.615 ;
        RECT 122.660 131.595 123.140 131.615 ;
        RECT 136.410 131.605 136.990 133.035 ;
        RECT 122.645 131.095 124.950 131.595 ;
        RECT 122.660 129.895 123.140 131.095 ;
        RECT 134.520 131.025 136.990 131.605 ;
        RECT 116.535 129.435 123.140 129.895 ;
        RECT 116.535 128.855 123.110 129.435 ;
        RECT 138.690 128.885 139.690 146.525 ;
        RECT 149.000 144.560 151.240 146.885 ;
        RECT 149.010 144.305 151.240 144.560 ;
        RECT 146.890 143.275 151.240 144.305 ;
        RECT 147.700 129.495 148.160 129.525 ;
        RECT 149.010 129.495 151.240 143.275 ;
        RECT 147.700 129.035 151.240 129.495 ;
        RECT 147.700 129.005 148.160 129.035 ;
        RECT 116.535 128.645 117.630 128.855 ;
        RECT 137.750 128.745 139.690 128.885 ;
        RECT 113.870 127.045 114.880 127.275 ;
        RECT 113.310 125.035 113.710 126.995 ;
        RECT 114.570 126.965 114.880 127.045 ;
        RECT 115.050 126.995 115.420 127.325 ;
        RECT 113.310 124.705 113.680 125.035 ;
        RECT 113.860 124.985 114.140 125.085 ;
        RECT 115.030 125.035 115.420 126.995 ;
        RECT 113.860 124.755 114.870 124.985 ;
        RECT 113.310 122.745 113.710 124.705 ;
        RECT 113.860 124.635 114.140 124.755 ;
        RECT 115.050 124.705 115.420 125.035 ;
        RECT 113.310 122.415 113.680 122.745 ;
        RECT 114.550 122.695 114.860 122.775 ;
        RECT 115.030 122.745 115.420 124.705 ;
        RECT 113.870 122.465 114.870 122.695 ;
        RECT 113.310 120.455 113.710 122.415 ;
        RECT 114.550 122.395 114.860 122.465 ;
        RECT 115.050 122.415 115.420 122.745 ;
        RECT 113.310 120.125 113.680 120.455 ;
        RECT 113.860 120.405 114.140 120.505 ;
        RECT 115.030 120.455 115.420 122.415 ;
        RECT 113.860 120.175 114.870 120.405 ;
        RECT 113.310 118.165 113.710 120.125 ;
        RECT 113.860 120.055 114.140 120.175 ;
        RECT 115.050 120.125 115.420 120.455 ;
        RECT 108.590 117.765 108.870 117.885 ;
        RECT 111.215 116.350 111.525 116.380 ;
        RECT 102.680 116.040 111.525 116.350 ;
        RECT 102.680 109.725 104.910 116.040 ;
        RECT 111.215 116.010 111.525 116.040 ;
        RECT 113.310 114.985 113.680 118.165 ;
        RECT 114.560 118.115 114.870 118.195 ;
        RECT 115.030 118.165 115.420 120.125 ;
        RECT 113.870 117.885 114.870 118.115 ;
        RECT 114.560 117.815 114.870 117.885 ;
        RECT 115.050 115.760 115.420 118.165 ;
        RECT 109.580 114.875 113.680 114.985 ;
        RECT 108.150 114.625 113.680 114.875 ;
        RECT 102.680 108.035 108.000 109.725 ;
        RECT 102.680 96.005 104.910 108.035 ;
        RECT 102.680 94.305 108.010 96.005 ;
        RECT 102.680 89.935 104.910 94.305 ;
        RECT 108.150 90.645 108.400 114.625 ;
        RECT 109.580 114.560 113.680 114.625 ;
        RECT 115.035 115.515 115.420 115.760 ;
        RECT 115.035 114.560 115.405 115.515 ;
        RECT 116.590 114.560 117.630 128.645 ;
        RECT 135.840 128.495 139.690 128.745 ;
        RECT 125.920 128.205 139.690 128.495 ;
        RECT 120.475 126.790 121.385 127.640 ;
        RECT 109.580 114.410 117.630 114.560 ;
        RECT 108.580 113.645 108.840 113.745 ;
        RECT 108.550 113.415 109.550 113.645 ;
        RECT 108.580 113.315 108.840 113.415 ;
        RECT 109.260 111.355 109.520 111.465 ;
        RECT 108.550 111.125 109.550 111.355 ;
        RECT 109.260 111.035 109.520 111.125 ;
        RECT 108.580 109.065 108.840 109.165 ;
        RECT 108.550 108.835 109.550 109.065 ;
        RECT 108.580 108.735 108.840 108.835 ;
        RECT 109.260 106.775 109.520 106.875 ;
        RECT 108.550 106.545 109.550 106.775 ;
        RECT 109.260 106.445 109.520 106.545 ;
        RECT 108.580 104.485 108.840 104.585 ;
        RECT 108.550 104.255 109.550 104.485 ;
        RECT 108.580 104.155 108.840 104.255 ;
        RECT 109.260 102.195 109.520 102.305 ;
        RECT 108.550 101.965 109.550 102.195 ;
        RECT 109.260 101.875 109.520 101.965 ;
        RECT 108.580 99.905 108.840 100.005 ;
        RECT 108.550 99.675 109.550 99.905 ;
        RECT 108.580 99.575 108.840 99.675 ;
        RECT 109.260 97.615 109.520 97.725 ;
        RECT 108.550 97.385 109.550 97.615 ;
        RECT 109.260 97.295 109.520 97.385 ;
        RECT 108.580 95.325 108.840 95.425 ;
        RECT 108.550 95.095 109.550 95.325 ;
        RECT 108.580 94.995 108.840 95.095 ;
        RECT 109.260 93.035 109.520 93.135 ;
        RECT 108.550 92.805 109.550 93.035 ;
        RECT 109.260 92.705 109.520 92.805 ;
        RECT 108.580 90.745 108.840 90.845 ;
        RECT 108.550 90.515 109.550 90.745 ;
        RECT 109.690 90.645 110.040 114.410 ;
        RECT 111.680 114.195 117.630 114.410 ;
        RECT 111.680 108.285 112.255 114.195 ;
        RECT 113.310 114.190 117.630 114.195 ;
        RECT 116.590 114.165 117.630 114.190 ;
        RECT 120.505 112.105 121.355 126.790 ;
        RECT 123.285 123.000 125.735 124.350 ;
        RECT 123.285 116.975 124.635 123.000 ;
        RECT 125.920 120.905 126.210 128.205 ;
        RECT 127.040 126.845 127.340 126.945 ;
        RECT 126.350 126.615 127.350 126.845 ;
        RECT 127.040 126.525 127.340 126.615 ;
        RECT 126.390 126.255 126.690 126.365 ;
        RECT 126.350 126.025 127.350 126.255 ;
        RECT 126.390 125.915 126.690 126.025 ;
        RECT 127.040 125.665 127.340 125.765 ;
        RECT 126.350 125.435 127.350 125.665 ;
        RECT 127.040 125.345 127.340 125.435 ;
        RECT 126.390 125.075 126.690 125.185 ;
        RECT 126.350 124.845 127.350 125.075 ;
        RECT 126.390 124.735 126.690 124.845 ;
        RECT 127.040 124.485 127.340 124.585 ;
        RECT 126.350 124.255 127.350 124.485 ;
        RECT 127.040 124.165 127.340 124.255 ;
        RECT 126.390 123.895 126.690 124.005 ;
        RECT 126.350 123.665 127.350 123.895 ;
        RECT 126.390 123.555 126.690 123.665 ;
        RECT 127.040 123.305 127.340 123.405 ;
        RECT 126.350 123.075 127.350 123.305 ;
        RECT 127.040 122.985 127.340 123.075 ;
        RECT 126.390 122.715 126.690 122.825 ;
        RECT 126.350 122.485 127.350 122.715 ;
        RECT 126.390 122.375 126.690 122.485 ;
        RECT 127.040 122.125 127.340 122.225 ;
        RECT 126.350 121.895 127.350 122.125 ;
        RECT 127.040 121.805 127.340 121.895 ;
        RECT 126.390 121.535 126.690 121.645 ;
        RECT 126.350 121.305 127.350 121.535 ;
        RECT 126.390 121.195 126.690 121.305 ;
        RECT 127.040 120.945 127.340 121.045 ;
        RECT 126.350 120.715 127.350 120.945 ;
        RECT 127.500 120.905 127.790 128.205 ;
        RECT 128.000 120.905 128.290 128.205 ;
        RECT 129.140 126.845 129.440 126.945 ;
        RECT 128.440 126.615 129.440 126.845 ;
        RECT 129.140 126.525 129.440 126.615 ;
        RECT 128.470 126.255 128.770 126.365 ;
        RECT 128.440 126.025 129.440 126.255 ;
        RECT 128.470 125.915 128.770 126.025 ;
        RECT 129.140 125.665 129.440 125.765 ;
        RECT 128.440 125.435 129.440 125.665 ;
        RECT 129.140 125.345 129.440 125.435 ;
        RECT 128.470 125.075 128.770 125.185 ;
        RECT 128.440 124.845 129.440 125.075 ;
        RECT 128.470 124.735 128.770 124.845 ;
        RECT 129.140 124.485 129.440 124.585 ;
        RECT 128.440 124.255 129.440 124.485 ;
        RECT 129.140 124.165 129.440 124.255 ;
        RECT 128.470 123.895 128.770 124.005 ;
        RECT 128.440 123.665 129.440 123.895 ;
        RECT 128.470 123.555 128.770 123.665 ;
        RECT 129.140 123.305 129.440 123.405 ;
        RECT 128.440 123.075 129.440 123.305 ;
        RECT 129.140 122.985 129.440 123.075 ;
        RECT 128.470 122.715 128.770 122.825 ;
        RECT 128.440 122.485 129.440 122.715 ;
        RECT 128.470 122.375 128.770 122.485 ;
        RECT 129.140 122.125 129.440 122.225 ;
        RECT 128.440 121.895 129.440 122.125 ;
        RECT 129.140 121.805 129.440 121.895 ;
        RECT 128.470 121.535 128.770 121.645 ;
        RECT 128.440 121.305 129.440 121.535 ;
        RECT 128.470 121.195 128.770 121.305 ;
        RECT 129.140 120.945 129.440 121.045 ;
        RECT 128.440 120.715 129.440 120.945 ;
        RECT 129.580 120.905 129.870 128.205 ;
        RECT 130.100 120.905 130.390 128.205 ;
        RECT 131.210 126.845 131.510 126.945 ;
        RECT 130.530 126.615 131.530 126.845 ;
        RECT 131.210 126.525 131.510 126.615 ;
        RECT 130.550 126.255 130.850 126.375 ;
        RECT 130.530 126.025 131.530 126.255 ;
        RECT 130.550 125.925 130.850 126.025 ;
        RECT 131.220 125.665 131.520 125.765 ;
        RECT 130.530 125.435 131.530 125.665 ;
        RECT 131.220 125.345 131.520 125.435 ;
        RECT 130.550 125.075 130.850 125.185 ;
        RECT 130.530 124.845 131.530 125.075 ;
        RECT 130.550 124.735 130.850 124.845 ;
        RECT 131.220 124.485 131.520 124.575 ;
        RECT 130.530 124.255 131.530 124.485 ;
        RECT 131.220 124.155 131.520 124.255 ;
        RECT 130.550 123.895 130.850 124.005 ;
        RECT 130.530 123.665 131.530 123.895 ;
        RECT 130.550 123.555 130.850 123.665 ;
        RECT 131.220 123.305 131.520 123.405 ;
        RECT 130.530 123.075 131.530 123.305 ;
        RECT 131.220 122.985 131.520 123.075 ;
        RECT 130.550 122.715 130.850 122.825 ;
        RECT 130.530 122.485 131.530 122.715 ;
        RECT 130.550 122.375 130.850 122.485 ;
        RECT 131.220 122.125 131.520 122.225 ;
        RECT 130.530 121.895 131.530 122.125 ;
        RECT 131.220 121.805 131.520 121.895 ;
        RECT 130.550 121.535 130.850 121.635 ;
        RECT 130.530 121.305 131.530 121.535 ;
        RECT 130.550 121.185 130.850 121.305 ;
        RECT 131.220 120.945 131.520 121.045 ;
        RECT 130.530 120.715 131.530 120.945 ;
        RECT 131.690 120.905 131.980 128.205 ;
        RECT 132.180 120.905 132.470 128.205 ;
        RECT 133.310 126.845 133.610 126.945 ;
        RECT 132.620 126.615 133.620 126.845 ;
        RECT 133.310 126.525 133.610 126.615 ;
        RECT 132.650 126.255 132.950 126.375 ;
        RECT 132.620 126.025 133.620 126.255 ;
        RECT 132.650 125.925 132.950 126.025 ;
        RECT 133.310 125.665 133.610 125.765 ;
        RECT 132.620 125.435 133.620 125.665 ;
        RECT 133.310 125.345 133.610 125.435 ;
        RECT 132.650 125.075 132.950 125.185 ;
        RECT 132.620 124.845 133.620 125.075 ;
        RECT 132.650 124.735 132.950 124.845 ;
        RECT 133.310 124.485 133.610 124.585 ;
        RECT 132.620 124.255 133.620 124.485 ;
        RECT 133.310 124.165 133.610 124.255 ;
        RECT 132.650 123.895 132.950 124.005 ;
        RECT 132.620 123.665 133.620 123.895 ;
        RECT 132.650 123.555 132.950 123.665 ;
        RECT 133.310 123.305 133.610 123.405 ;
        RECT 132.620 123.075 133.620 123.305 ;
        RECT 133.310 122.985 133.610 123.075 ;
        RECT 132.650 122.715 132.950 122.825 ;
        RECT 132.620 122.485 133.620 122.715 ;
        RECT 132.650 122.375 132.950 122.485 ;
        RECT 133.310 122.125 133.610 122.225 ;
        RECT 132.620 121.895 133.620 122.125 ;
        RECT 133.310 121.805 133.610 121.895 ;
        RECT 132.650 121.535 132.950 121.645 ;
        RECT 132.620 121.305 133.620 121.535 ;
        RECT 132.650 121.195 132.950 121.305 ;
        RECT 133.310 120.945 133.610 121.035 ;
        RECT 132.620 120.715 133.620 120.945 ;
        RECT 133.770 120.905 134.060 128.205 ;
        RECT 134.260 120.905 134.550 128.205 ;
        RECT 135.840 128.020 139.690 128.205 ;
        RECT 145.860 128.105 146.140 128.195 ;
        RECT 135.400 126.845 135.700 126.935 ;
        RECT 134.710 126.615 135.710 126.845 ;
        RECT 135.400 126.515 135.700 126.615 ;
        RECT 134.720 126.255 135.020 126.365 ;
        RECT 134.710 126.025 135.710 126.255 ;
        RECT 134.720 125.915 135.020 126.025 ;
        RECT 135.400 125.665 135.700 125.765 ;
        RECT 134.710 125.435 135.710 125.665 ;
        RECT 135.400 125.345 135.700 125.435 ;
        RECT 134.730 125.075 135.030 125.185 ;
        RECT 134.710 124.845 135.710 125.075 ;
        RECT 134.730 124.735 135.030 124.845 ;
        RECT 135.400 124.485 135.700 124.585 ;
        RECT 134.710 124.255 135.710 124.485 ;
        RECT 135.400 124.165 135.700 124.255 ;
        RECT 134.730 123.895 135.030 124.005 ;
        RECT 134.710 123.665 135.710 123.895 ;
        RECT 134.730 123.555 135.030 123.665 ;
        RECT 135.400 123.305 135.700 123.405 ;
        RECT 134.710 123.075 135.710 123.305 ;
        RECT 135.400 122.985 135.700 123.075 ;
        RECT 134.730 122.715 135.030 122.835 ;
        RECT 134.710 122.485 135.710 122.715 ;
        RECT 134.730 122.385 135.030 122.485 ;
        RECT 135.400 122.125 135.700 122.225 ;
        RECT 134.710 121.895 135.710 122.125 ;
        RECT 135.400 121.805 135.700 121.895 ;
        RECT 134.730 121.535 135.030 121.645 ;
        RECT 134.710 121.305 135.710 121.535 ;
        RECT 134.730 121.195 135.030 121.305 ;
        RECT 135.400 120.945 135.700 121.045 ;
        RECT 134.710 120.715 135.710 120.945 ;
        RECT 135.850 120.905 136.140 128.020 ;
        RECT 137.750 127.885 139.690 128.020 ;
        RECT 127.040 120.625 127.340 120.715 ;
        RECT 129.140 120.625 129.440 120.715 ;
        RECT 131.220 120.625 131.520 120.715 ;
        RECT 133.310 120.615 133.610 120.715 ;
        RECT 135.400 120.625 135.700 120.715 ;
        RECT 144.710 120.185 145.010 127.885 ;
        RECT 145.185 127.875 146.185 128.105 ;
        RECT 145.860 127.785 146.140 127.875 ;
        RECT 145.230 126.815 145.530 126.915 ;
        RECT 145.185 126.585 146.185 126.815 ;
        RECT 145.230 126.495 145.530 126.585 ;
        RECT 145.870 125.525 146.150 125.625 ;
        RECT 145.185 125.295 146.185 125.525 ;
        RECT 145.870 125.215 146.150 125.295 ;
        RECT 145.230 124.235 145.530 124.335 ;
        RECT 145.185 124.005 146.185 124.235 ;
        RECT 145.230 123.915 145.530 124.005 ;
        RECT 145.880 122.945 146.160 123.035 ;
        RECT 145.185 122.715 146.185 122.945 ;
        RECT 145.880 122.625 146.160 122.715 ;
        RECT 145.230 121.655 145.530 121.755 ;
        RECT 145.185 121.425 146.185 121.655 ;
        RECT 145.230 121.335 145.530 121.425 ;
        RECT 145.170 120.390 145.500 120.660 ;
        RECT 145.200 120.185 145.470 120.390 ;
        RECT 146.350 120.185 146.650 127.885 ;
        RECT 149.010 125.475 151.240 129.035 ;
        RECT 146.810 124.015 151.240 125.475 ;
        RECT 144.710 119.655 146.650 120.185 ;
        RECT 127.050 119.305 127.340 119.405 ;
        RECT 129.150 119.305 129.440 119.405 ;
        RECT 131.230 119.305 131.520 119.405 ;
        RECT 133.310 119.305 133.600 119.405 ;
        RECT 135.400 119.305 135.690 119.405 ;
        RECT 123.220 115.550 125.740 116.975 ;
        RECT 116.550 112.090 121.355 112.105 ;
        RECT 116.550 111.910 124.985 112.090 ;
        RECT 116.550 111.810 125.530 111.910 ;
        RECT 125.920 111.810 126.210 119.095 ;
        RECT 126.350 119.075 127.350 119.305 ;
        RECT 127.050 118.985 127.340 119.075 ;
        RECT 126.400 118.715 126.700 118.805 ;
        RECT 126.350 118.485 127.350 118.715 ;
        RECT 126.400 118.405 126.700 118.485 ;
        RECT 127.050 118.125 127.340 118.225 ;
        RECT 126.350 117.895 127.350 118.125 ;
        RECT 127.050 117.805 127.340 117.895 ;
        RECT 126.400 117.535 126.700 117.625 ;
        RECT 126.350 117.305 127.350 117.535 ;
        RECT 126.400 117.225 126.700 117.305 ;
        RECT 127.050 116.945 127.340 117.045 ;
        RECT 126.350 116.715 127.350 116.945 ;
        RECT 127.050 116.625 127.340 116.715 ;
        RECT 126.400 116.355 126.700 116.445 ;
        RECT 126.350 116.125 127.350 116.355 ;
        RECT 126.400 116.045 126.700 116.125 ;
        RECT 127.050 115.765 127.340 115.865 ;
        RECT 126.350 115.535 127.350 115.765 ;
        RECT 127.050 115.445 127.340 115.535 ;
        RECT 126.400 115.175 126.700 115.255 ;
        RECT 126.350 114.945 127.350 115.175 ;
        RECT 126.400 114.855 126.700 114.945 ;
        RECT 127.050 114.585 127.340 114.695 ;
        RECT 126.350 114.355 127.350 114.585 ;
        RECT 127.050 114.275 127.340 114.355 ;
        RECT 126.400 113.995 126.700 114.085 ;
        RECT 126.350 113.765 127.350 113.995 ;
        RECT 126.400 113.685 126.700 113.765 ;
        RECT 127.050 113.405 127.340 113.505 ;
        RECT 126.350 113.175 127.350 113.405 ;
        RECT 127.050 113.085 127.340 113.175 ;
        RECT 127.500 111.810 127.790 119.065 ;
        RECT 128.000 111.810 128.290 119.095 ;
        RECT 128.440 119.075 129.440 119.305 ;
        RECT 129.150 118.985 129.440 119.075 ;
        RECT 128.490 118.715 128.790 118.805 ;
        RECT 128.440 118.485 129.440 118.715 ;
        RECT 128.490 118.405 128.790 118.485 ;
        RECT 129.150 118.125 129.440 118.225 ;
        RECT 128.440 117.895 129.440 118.125 ;
        RECT 129.150 117.805 129.440 117.895 ;
        RECT 128.490 117.535 128.790 117.625 ;
        RECT 128.440 117.305 129.440 117.535 ;
        RECT 128.490 117.225 128.790 117.305 ;
        RECT 129.150 116.945 129.440 117.045 ;
        RECT 128.440 116.715 129.440 116.945 ;
        RECT 129.150 116.625 129.440 116.715 ;
        RECT 128.490 116.355 128.790 116.445 ;
        RECT 128.440 116.125 129.440 116.355 ;
        RECT 128.490 116.045 128.790 116.125 ;
        RECT 129.150 115.765 129.440 115.865 ;
        RECT 128.440 115.535 129.440 115.765 ;
        RECT 129.150 115.445 129.440 115.535 ;
        RECT 128.490 115.175 128.790 115.265 ;
        RECT 128.440 114.945 129.440 115.175 ;
        RECT 128.490 114.865 128.790 114.945 ;
        RECT 129.150 114.585 129.440 114.685 ;
        RECT 128.440 114.355 129.440 114.585 ;
        RECT 129.150 114.265 129.440 114.355 ;
        RECT 128.490 113.995 128.790 114.085 ;
        RECT 128.440 113.765 129.440 113.995 ;
        RECT 128.490 113.685 128.790 113.765 ;
        RECT 129.150 113.405 129.440 113.505 ;
        RECT 128.440 113.175 129.440 113.405 ;
        RECT 129.150 113.085 129.440 113.175 ;
        RECT 129.580 111.810 129.870 119.095 ;
        RECT 130.100 111.810 130.390 119.095 ;
        RECT 130.530 119.075 131.530 119.305 ;
        RECT 131.230 118.985 131.520 119.075 ;
        RECT 130.570 118.715 130.870 118.805 ;
        RECT 130.530 118.485 131.530 118.715 ;
        RECT 130.570 118.405 130.870 118.485 ;
        RECT 131.230 118.125 131.520 118.225 ;
        RECT 130.530 117.895 131.530 118.125 ;
        RECT 131.230 117.805 131.520 117.895 ;
        RECT 130.570 117.535 130.870 117.625 ;
        RECT 130.530 117.305 131.530 117.535 ;
        RECT 130.570 117.225 130.870 117.305 ;
        RECT 131.230 116.945 131.520 117.035 ;
        RECT 130.530 116.715 131.530 116.945 ;
        RECT 131.230 116.615 131.520 116.715 ;
        RECT 130.570 116.355 130.870 116.445 ;
        RECT 130.530 116.125 131.530 116.355 ;
        RECT 130.570 116.045 130.870 116.125 ;
        RECT 131.230 115.765 131.520 115.865 ;
        RECT 130.530 115.535 131.530 115.765 ;
        RECT 131.230 115.445 131.520 115.535 ;
        RECT 130.570 115.175 130.870 115.265 ;
        RECT 130.530 114.945 131.530 115.175 ;
        RECT 130.570 114.865 130.870 114.945 ;
        RECT 131.230 114.585 131.520 114.685 ;
        RECT 130.530 114.355 131.530 114.585 ;
        RECT 131.230 114.265 131.520 114.355 ;
        RECT 130.570 113.995 130.870 114.085 ;
        RECT 130.530 113.765 131.530 113.995 ;
        RECT 130.570 113.685 130.870 113.765 ;
        RECT 131.240 113.405 131.530 113.505 ;
        RECT 130.530 113.175 131.530 113.405 ;
        RECT 131.240 113.085 131.530 113.175 ;
        RECT 131.690 111.810 131.980 119.095 ;
        RECT 132.180 111.810 132.470 119.095 ;
        RECT 132.620 119.075 133.620 119.305 ;
        RECT 133.310 118.985 133.600 119.075 ;
        RECT 132.630 118.715 132.930 118.805 ;
        RECT 132.620 118.485 133.620 118.715 ;
        RECT 132.630 118.405 132.930 118.485 ;
        RECT 133.310 118.125 133.600 118.225 ;
        RECT 132.620 117.895 133.620 118.125 ;
        RECT 133.310 117.805 133.600 117.895 ;
        RECT 132.630 117.535 132.930 117.625 ;
        RECT 132.620 117.305 133.620 117.535 ;
        RECT 132.630 117.225 132.930 117.305 ;
        RECT 133.310 116.945 133.600 117.045 ;
        RECT 132.620 116.715 133.620 116.945 ;
        RECT 133.310 116.625 133.600 116.715 ;
        RECT 132.630 116.355 132.930 116.445 ;
        RECT 132.620 116.125 133.620 116.355 ;
        RECT 132.630 116.045 132.930 116.125 ;
        RECT 133.310 115.765 133.600 115.865 ;
        RECT 132.620 115.535 133.620 115.765 ;
        RECT 133.310 115.445 133.600 115.535 ;
        RECT 132.630 115.175 132.930 115.265 ;
        RECT 132.620 114.945 133.620 115.175 ;
        RECT 132.630 114.865 132.930 114.945 ;
        RECT 133.310 114.585 133.600 114.685 ;
        RECT 132.620 114.355 133.620 114.585 ;
        RECT 133.310 114.265 133.600 114.355 ;
        RECT 132.630 113.995 132.930 114.085 ;
        RECT 132.620 113.765 133.620 113.995 ;
        RECT 132.630 113.685 132.930 113.765 ;
        RECT 133.310 113.405 133.600 113.505 ;
        RECT 132.620 113.175 133.620 113.405 ;
        RECT 133.310 113.085 133.600 113.175 ;
        RECT 133.770 111.810 134.060 119.095 ;
        RECT 134.260 111.810 134.550 119.095 ;
        RECT 134.710 119.075 135.710 119.305 ;
        RECT 135.400 118.985 135.690 119.075 ;
        RECT 134.730 118.715 135.030 118.805 ;
        RECT 134.710 118.485 135.710 118.715 ;
        RECT 134.730 118.405 135.030 118.485 ;
        RECT 135.400 118.125 135.690 118.225 ;
        RECT 134.710 117.895 135.710 118.125 ;
        RECT 135.400 117.805 135.690 117.895 ;
        RECT 134.730 117.535 135.030 117.625 ;
        RECT 134.710 117.305 135.710 117.535 ;
        RECT 134.730 117.225 135.030 117.305 ;
        RECT 135.400 116.945 135.690 117.045 ;
        RECT 134.710 116.715 135.710 116.945 ;
        RECT 135.400 116.625 135.690 116.715 ;
        RECT 134.730 116.355 135.030 116.445 ;
        RECT 134.710 116.125 135.710 116.355 ;
        RECT 134.730 116.045 135.030 116.125 ;
        RECT 135.400 115.765 135.690 115.865 ;
        RECT 134.710 115.535 135.710 115.765 ;
        RECT 135.400 115.445 135.690 115.535 ;
        RECT 134.730 115.175 135.030 115.265 ;
        RECT 134.710 114.945 135.710 115.175 ;
        RECT 134.730 114.865 135.030 114.945 ;
        RECT 135.400 114.585 135.690 114.685 ;
        RECT 134.710 114.355 135.710 114.585 ;
        RECT 135.400 114.265 135.690 114.355 ;
        RECT 134.730 113.995 135.030 114.085 ;
        RECT 134.710 113.765 135.710 113.995 ;
        RECT 134.730 113.685 135.030 113.765 ;
        RECT 135.400 113.405 135.690 113.505 ;
        RECT 134.710 113.175 135.710 113.405 ;
        RECT 135.400 113.085 135.690 113.175 ;
        RECT 135.850 111.810 136.140 119.095 ;
        RECT 116.550 111.520 136.140 111.810 ;
        RECT 144.710 111.795 145.010 119.655 ;
        RECT 145.190 118.325 145.490 118.415 ;
        RECT 145.155 118.095 146.155 118.325 ;
        RECT 145.190 117.995 145.490 118.095 ;
        RECT 145.880 117.035 146.160 117.135 ;
        RECT 145.155 116.805 146.160 117.035 ;
        RECT 145.880 116.725 146.160 116.805 ;
        RECT 145.190 115.745 145.490 115.845 ;
        RECT 145.155 115.515 146.155 115.745 ;
        RECT 145.190 115.425 145.490 115.515 ;
        RECT 145.880 114.455 146.160 114.545 ;
        RECT 145.155 114.225 146.160 114.455 ;
        RECT 145.880 114.135 146.160 114.225 ;
        RECT 145.190 113.165 145.490 113.255 ;
        RECT 145.155 112.935 146.155 113.165 ;
        RECT 145.190 112.835 145.490 112.935 ;
        RECT 145.880 111.875 146.160 111.965 ;
        RECT 145.155 111.645 146.160 111.875 ;
        RECT 146.350 111.795 146.650 119.655 ;
        RECT 149.010 115.655 151.240 124.015 ;
        RECT 146.800 114.195 151.240 115.655 ;
        RECT 145.880 111.555 146.160 111.645 ;
        RECT 116.550 111.415 125.530 111.520 ;
        RECT 125.920 111.505 126.210 111.520 ;
        RECT 127.500 111.475 127.790 111.520 ;
        RECT 128.000 111.505 128.290 111.520 ;
        RECT 129.580 111.505 129.870 111.520 ;
        RECT 130.100 111.505 130.390 111.520 ;
        RECT 131.690 111.505 131.980 111.520 ;
        RECT 132.180 111.505 132.470 111.520 ;
        RECT 133.770 111.505 134.060 111.520 ;
        RECT 134.260 111.505 134.550 111.520 ;
        RECT 135.850 111.505 136.140 111.520 ;
        RECT 116.550 111.240 124.985 111.415 ;
        RECT 147.690 110.715 148.165 110.745 ;
        RECT 149.010 110.715 151.240 114.195 ;
        RECT 147.690 110.240 151.240 110.715 ;
        RECT 147.690 110.210 148.165 110.240 ;
        RECT 116.425 109.955 116.765 109.975 ;
        RECT 118.430 109.955 119.230 109.985 ;
        RECT 116.425 109.155 119.230 109.955 ;
        RECT 116.425 109.005 116.765 109.155 ;
        RECT 118.430 109.125 119.230 109.155 ;
        RECT 110.995 107.710 112.255 108.285 ;
        RECT 113.770 108.655 116.770 109.005 ;
        RECT 108.580 90.415 108.840 90.515 ;
        RECT 102.680 89.715 107.320 89.935 ;
        RECT 102.680 89.310 107.525 89.715 ;
        RECT 102.680 89.095 107.320 89.310 ;
        RECT 102.680 83.575 104.910 89.095 ;
        RECT 110.995 88.885 111.570 107.710 ;
        RECT 112.840 100.400 113.630 103.855 ;
        RECT 112.115 99.745 113.630 100.400 ;
        RECT 112.115 99.525 113.500 99.745 ;
        RECT 112.115 98.020 112.990 99.525 ;
        RECT 113.770 95.455 114.120 108.655 ;
        RECT 114.280 107.365 114.700 107.475 ;
        RECT 114.280 107.135 116.280 107.365 ;
        RECT 114.280 107.035 114.700 107.135 ;
        RECT 115.800 106.775 116.220 106.855 ;
        RECT 114.280 106.545 116.280 106.775 ;
        RECT 115.800 106.455 116.220 106.545 ;
        RECT 114.280 106.185 114.700 106.295 ;
        RECT 114.280 105.955 116.280 106.185 ;
        RECT 114.280 105.855 114.700 105.955 ;
        RECT 115.800 105.595 116.220 105.675 ;
        RECT 114.280 105.365 116.280 105.595 ;
        RECT 115.800 105.275 116.220 105.365 ;
        RECT 114.280 105.005 114.700 105.105 ;
        RECT 114.280 104.775 116.280 105.005 ;
        RECT 114.280 104.665 114.700 104.775 ;
        RECT 115.800 104.415 116.220 104.505 ;
        RECT 114.280 104.185 116.280 104.415 ;
        RECT 115.800 104.105 116.220 104.185 ;
        RECT 114.280 103.825 114.700 103.925 ;
        RECT 114.280 103.595 116.280 103.825 ;
        RECT 114.280 103.485 114.700 103.595 ;
        RECT 115.800 103.235 116.220 103.325 ;
        RECT 114.280 103.005 116.280 103.235 ;
        RECT 115.800 102.925 116.220 103.005 ;
        RECT 114.280 102.645 114.700 102.745 ;
        RECT 114.280 102.415 116.280 102.645 ;
        RECT 114.280 102.305 114.700 102.415 ;
        RECT 115.800 102.055 116.220 102.145 ;
        RECT 114.280 101.825 116.280 102.055 ;
        RECT 115.800 101.745 116.220 101.825 ;
        RECT 114.280 101.465 114.700 101.565 ;
        RECT 114.280 101.235 116.280 101.465 ;
        RECT 114.280 101.125 114.700 101.235 ;
        RECT 115.800 100.875 116.220 100.965 ;
        RECT 114.280 100.645 116.280 100.875 ;
        RECT 115.800 100.565 116.220 100.645 ;
        RECT 114.280 100.285 114.700 100.385 ;
        RECT 114.280 100.055 116.280 100.285 ;
        RECT 114.280 99.945 114.700 100.055 ;
        RECT 115.800 99.695 116.220 99.785 ;
        RECT 114.280 99.465 116.280 99.695 ;
        RECT 115.800 99.385 116.220 99.465 ;
        RECT 114.290 99.105 114.710 99.205 ;
        RECT 114.280 98.875 116.280 99.105 ;
        RECT 114.290 98.765 114.710 98.875 ;
        RECT 115.800 98.515 116.220 98.605 ;
        RECT 114.280 98.285 116.280 98.515 ;
        RECT 115.800 98.205 116.220 98.285 ;
        RECT 114.290 97.925 114.710 98.025 ;
        RECT 114.280 97.695 116.280 97.925 ;
        RECT 114.290 97.585 114.710 97.695 ;
        RECT 115.800 97.335 116.220 97.425 ;
        RECT 114.280 97.105 116.280 97.335 ;
        RECT 115.800 97.025 116.220 97.105 ;
        RECT 114.290 96.745 114.710 96.845 ;
        RECT 114.280 96.515 116.280 96.745 ;
        RECT 114.290 96.405 114.710 96.515 ;
        RECT 115.800 96.155 116.220 96.245 ;
        RECT 114.280 95.925 116.280 96.155 ;
        RECT 115.800 95.845 116.220 95.925 ;
        RECT 114.290 95.565 114.710 95.665 ;
        RECT 114.280 95.335 116.280 95.565 ;
        RECT 116.420 95.455 116.770 108.655 ;
        RECT 123.760 107.755 124.190 107.865 ;
        RECT 127.400 107.755 127.830 107.865 ;
        RECT 131.150 107.755 131.580 107.865 ;
        RECT 134.790 107.755 135.220 107.865 ;
        RECT 138.500 107.755 138.930 107.865 ;
        RECT 142.140 107.755 142.570 107.865 ;
        RECT 145.830 107.755 146.260 107.865 ;
        RECT 114.290 95.225 114.710 95.335 ;
        RECT 110.990 88.295 113.640 88.885 ;
        RECT 108.160 88.055 113.640 88.295 ;
        RECT 102.680 81.855 108.020 83.575 ;
        RECT 102.680 69.595 104.910 81.855 ;
        RECT 102.680 67.865 108.010 69.595 ;
        RECT 102.680 63.670 104.910 67.865 ;
        RECT 108.160 64.345 108.400 88.055 ;
        RECT 108.550 87.325 108.930 87.465 ;
        RECT 108.550 87.095 109.560 87.325 ;
        RECT 108.550 86.995 108.930 87.095 ;
        RECT 109.200 85.035 109.570 85.155 ;
        RECT 108.560 84.805 109.570 85.035 ;
        RECT 109.200 84.665 109.570 84.805 ;
        RECT 108.550 82.745 108.930 82.865 ;
        RECT 108.550 82.515 109.560 82.745 ;
        RECT 108.550 82.395 108.930 82.515 ;
        RECT 109.200 80.455 109.570 80.585 ;
        RECT 108.560 80.225 109.570 80.455 ;
        RECT 109.200 80.095 109.570 80.225 ;
        RECT 108.550 78.165 108.930 78.285 ;
        RECT 108.550 77.935 109.560 78.165 ;
        RECT 108.550 77.815 108.930 77.935 ;
        RECT 109.200 75.875 109.570 76.005 ;
        RECT 108.560 75.645 109.570 75.875 ;
        RECT 109.200 75.515 109.570 75.645 ;
        RECT 108.550 73.585 108.930 73.705 ;
        RECT 108.550 73.355 109.560 73.585 ;
        RECT 108.550 73.235 108.930 73.355 ;
        RECT 109.200 71.295 109.570 71.435 ;
        RECT 108.560 71.065 109.570 71.295 ;
        RECT 109.200 70.945 109.570 71.065 ;
        RECT 108.550 69.005 108.930 69.125 ;
        RECT 108.550 68.775 109.560 69.005 ;
        RECT 108.550 68.655 108.930 68.775 ;
        RECT 109.200 66.715 109.570 66.835 ;
        RECT 108.560 66.485 109.570 66.715 ;
        RECT 109.200 66.345 109.570 66.485 ;
        RECT 108.550 64.425 108.930 64.545 ;
        RECT 108.550 64.195 109.560 64.425 ;
        RECT 109.720 64.345 109.960 88.055 ;
        RECT 108.550 64.075 108.930 64.195 ;
        RECT 102.680 62.945 107.555 63.670 ;
        RECT 102.680 57.715 104.910 62.945 ;
        RECT 112.560 62.765 113.635 88.055 ;
        RECT 117.880 80.155 118.960 80.185 ;
        RECT 121.250 80.155 121.500 107.535 ;
        RECT 121.695 107.525 124.195 107.755 ;
        RECT 123.760 107.425 124.190 107.525 ;
        RECT 121.700 106.465 122.210 106.585 ;
        RECT 121.695 106.235 124.195 106.465 ;
        RECT 121.700 106.115 122.210 106.235 ;
        RECT 123.760 105.175 124.190 105.285 ;
        RECT 121.695 104.945 124.195 105.175 ;
        RECT 123.760 104.845 124.190 104.945 ;
        RECT 121.700 103.885 122.210 104.005 ;
        RECT 121.695 103.655 124.195 103.885 ;
        RECT 121.700 103.535 122.210 103.655 ;
        RECT 123.760 102.595 124.190 102.695 ;
        RECT 121.695 102.365 124.195 102.595 ;
        RECT 123.760 102.255 124.190 102.365 ;
        RECT 121.700 101.305 122.210 101.415 ;
        RECT 121.695 101.075 124.195 101.305 ;
        RECT 121.700 100.945 122.210 101.075 ;
        RECT 123.760 100.015 124.190 100.125 ;
        RECT 121.695 99.785 124.195 100.015 ;
        RECT 123.760 99.685 124.190 99.785 ;
        RECT 121.660 98.725 122.170 98.855 ;
        RECT 121.660 98.495 124.195 98.725 ;
        RECT 121.660 98.385 122.170 98.495 ;
        RECT 123.770 97.435 124.200 97.545 ;
        RECT 121.695 97.205 124.200 97.435 ;
        RECT 123.770 97.105 124.200 97.205 ;
        RECT 121.700 96.145 122.210 96.265 ;
        RECT 121.695 95.915 124.195 96.145 ;
        RECT 121.700 95.795 122.210 95.915 ;
        RECT 123.770 94.855 124.200 94.955 ;
        RECT 121.695 94.625 124.200 94.855 ;
        RECT 123.770 94.515 124.200 94.625 ;
        RECT 121.700 93.565 122.210 93.685 ;
        RECT 121.695 93.335 124.195 93.565 ;
        RECT 121.700 93.215 122.210 93.335 ;
        RECT 123.770 92.275 124.200 92.385 ;
        RECT 121.695 92.045 124.200 92.275 ;
        RECT 123.770 91.945 124.200 92.045 ;
        RECT 121.690 90.985 122.200 91.105 ;
        RECT 121.690 90.755 124.195 90.985 ;
        RECT 121.690 90.635 122.200 90.755 ;
        RECT 123.770 89.695 124.200 89.795 ;
        RECT 121.695 89.465 124.200 89.695 ;
        RECT 123.770 89.355 124.200 89.465 ;
        RECT 121.680 88.405 122.190 88.525 ;
        RECT 121.680 88.175 124.195 88.405 ;
        RECT 121.680 88.055 122.190 88.175 ;
        RECT 123.770 87.115 124.200 87.225 ;
        RECT 121.695 86.885 124.200 87.115 ;
        RECT 123.770 86.785 124.200 86.885 ;
        RECT 121.690 85.825 122.200 85.945 ;
        RECT 121.690 85.595 124.195 85.825 ;
        RECT 121.690 85.475 122.200 85.595 ;
        RECT 123.770 84.535 124.200 84.645 ;
        RECT 121.695 84.305 124.200 84.535 ;
        RECT 123.770 84.205 124.200 84.305 ;
        RECT 121.690 83.245 122.200 83.365 ;
        RECT 121.690 83.015 124.195 83.245 ;
        RECT 121.690 82.895 122.200 83.015 ;
        RECT 123.770 81.955 124.200 82.055 ;
        RECT 121.695 81.725 124.200 81.955 ;
        RECT 123.770 81.615 124.200 81.725 ;
        RECT 124.400 80.155 124.650 107.535 ;
        RECT 124.940 80.155 125.190 107.545 ;
        RECT 125.375 107.525 127.875 107.755 ;
        RECT 127.400 107.425 127.830 107.525 ;
        RECT 125.350 106.465 125.860 106.585 ;
        RECT 125.350 106.235 127.875 106.465 ;
        RECT 125.350 106.115 125.860 106.235 ;
        RECT 127.400 105.175 127.830 105.285 ;
        RECT 125.375 104.945 127.875 105.175 ;
        RECT 127.400 104.845 127.830 104.945 ;
        RECT 125.370 103.885 125.880 104.005 ;
        RECT 125.370 103.655 127.875 103.885 ;
        RECT 125.370 103.535 125.880 103.655 ;
        RECT 127.400 102.595 127.830 102.705 ;
        RECT 125.375 102.365 127.875 102.595 ;
        RECT 127.400 102.265 127.830 102.365 ;
        RECT 125.350 101.305 125.860 101.425 ;
        RECT 125.350 101.075 127.875 101.305 ;
        RECT 125.350 100.955 125.860 101.075 ;
        RECT 127.400 100.015 127.830 100.125 ;
        RECT 125.375 99.785 127.875 100.015 ;
        RECT 127.400 99.685 127.830 99.785 ;
        RECT 125.370 98.725 125.880 98.845 ;
        RECT 125.370 98.495 127.875 98.725 ;
        RECT 125.370 98.375 125.880 98.495 ;
        RECT 127.400 97.435 127.830 97.545 ;
        RECT 125.375 97.205 127.875 97.435 ;
        RECT 127.400 97.105 127.830 97.205 ;
        RECT 125.390 96.145 125.900 96.255 ;
        RECT 125.375 95.915 127.875 96.145 ;
        RECT 125.390 95.785 125.900 95.915 ;
        RECT 127.400 94.855 127.830 94.965 ;
        RECT 125.375 94.625 127.875 94.855 ;
        RECT 127.400 94.525 127.830 94.625 ;
        RECT 125.370 93.565 125.880 93.685 ;
        RECT 125.370 93.335 127.875 93.565 ;
        RECT 125.370 93.215 125.880 93.335 ;
        RECT 127.400 92.275 127.830 92.395 ;
        RECT 125.375 92.045 127.875 92.275 ;
        RECT 127.400 91.955 127.830 92.045 ;
        RECT 125.380 90.985 125.890 91.105 ;
        RECT 125.375 90.755 127.875 90.985 ;
        RECT 125.380 90.635 125.890 90.755 ;
        RECT 127.400 89.695 127.830 89.805 ;
        RECT 125.375 89.465 127.875 89.695 ;
        RECT 127.400 89.365 127.830 89.465 ;
        RECT 125.370 88.405 125.880 88.525 ;
        RECT 125.370 88.175 127.875 88.405 ;
        RECT 125.370 88.055 125.880 88.175 ;
        RECT 127.400 87.115 127.830 87.225 ;
        RECT 125.375 86.885 127.875 87.115 ;
        RECT 127.400 86.785 127.830 86.885 ;
        RECT 125.370 85.825 125.880 85.935 ;
        RECT 125.370 85.595 127.875 85.825 ;
        RECT 125.370 85.465 125.880 85.595 ;
        RECT 127.400 84.535 127.830 84.645 ;
        RECT 125.375 84.305 127.875 84.535 ;
        RECT 127.400 84.205 127.830 84.305 ;
        RECT 125.370 83.245 125.880 83.375 ;
        RECT 125.370 83.015 127.875 83.245 ;
        RECT 125.370 82.905 125.880 83.015 ;
        RECT 127.400 81.955 127.830 82.055 ;
        RECT 125.375 81.725 127.875 81.955 ;
        RECT 127.400 81.615 127.830 81.725 ;
        RECT 128.080 80.155 128.330 107.535 ;
        RECT 128.620 80.155 128.870 107.535 ;
        RECT 129.055 107.525 131.580 107.755 ;
        RECT 131.150 107.425 131.580 107.525 ;
        RECT 129.060 106.465 129.570 106.585 ;
        RECT 129.055 106.235 131.555 106.465 ;
        RECT 129.060 106.115 129.570 106.235 ;
        RECT 131.150 105.175 131.580 105.285 ;
        RECT 129.055 104.945 131.580 105.175 ;
        RECT 131.150 104.845 131.580 104.945 ;
        RECT 129.060 103.885 129.570 104.005 ;
        RECT 129.055 103.655 131.555 103.885 ;
        RECT 129.060 103.535 129.570 103.655 ;
        RECT 131.150 102.595 131.580 102.715 ;
        RECT 129.055 102.365 131.580 102.595 ;
        RECT 131.150 102.275 131.580 102.365 ;
        RECT 129.030 101.305 129.540 101.425 ;
        RECT 129.030 101.075 131.555 101.305 ;
        RECT 129.030 100.955 129.540 101.075 ;
        RECT 131.150 100.015 131.580 100.125 ;
        RECT 129.055 99.785 131.580 100.015 ;
        RECT 131.150 99.685 131.580 99.785 ;
        RECT 129.060 98.725 129.570 98.845 ;
        RECT 129.055 98.495 131.555 98.725 ;
        RECT 129.060 98.375 129.570 98.495 ;
        RECT 131.150 97.435 131.580 97.545 ;
        RECT 129.055 97.205 131.580 97.435 ;
        RECT 131.150 97.105 131.580 97.205 ;
        RECT 129.050 96.145 129.560 96.265 ;
        RECT 129.050 95.915 131.555 96.145 ;
        RECT 129.050 95.795 129.560 95.915 ;
        RECT 131.150 94.855 131.580 94.965 ;
        RECT 129.055 94.625 131.580 94.855 ;
        RECT 131.150 94.525 131.580 94.625 ;
        RECT 129.050 93.565 129.560 93.685 ;
        RECT 129.050 93.335 131.555 93.565 ;
        RECT 129.050 93.215 129.560 93.335 ;
        RECT 131.150 92.275 131.580 92.385 ;
        RECT 129.055 92.045 131.580 92.275 ;
        RECT 131.150 91.945 131.580 92.045 ;
        RECT 129.050 90.985 129.560 91.105 ;
        RECT 129.050 90.755 131.555 90.985 ;
        RECT 129.050 90.635 129.560 90.755 ;
        RECT 131.150 89.695 131.580 89.805 ;
        RECT 129.055 89.465 131.580 89.695 ;
        RECT 131.150 89.365 131.580 89.465 ;
        RECT 129.050 88.405 129.560 88.525 ;
        RECT 129.050 88.175 131.555 88.405 ;
        RECT 129.050 88.055 129.560 88.175 ;
        RECT 131.150 87.115 131.580 87.225 ;
        RECT 129.055 86.885 131.580 87.115 ;
        RECT 131.150 86.785 131.580 86.885 ;
        RECT 129.040 85.825 129.550 85.945 ;
        RECT 129.040 85.595 131.555 85.825 ;
        RECT 129.040 85.475 129.550 85.595 ;
        RECT 131.150 84.535 131.580 84.645 ;
        RECT 129.055 84.305 131.580 84.535 ;
        RECT 131.150 84.205 131.580 84.305 ;
        RECT 129.050 83.245 129.560 83.365 ;
        RECT 129.050 83.015 131.555 83.245 ;
        RECT 129.050 82.895 129.560 83.015 ;
        RECT 131.150 81.955 131.580 82.055 ;
        RECT 129.055 81.725 131.580 81.955 ;
        RECT 131.150 81.615 131.580 81.725 ;
        RECT 131.750 80.155 132.000 107.535 ;
        RECT 132.300 80.155 132.550 107.535 ;
        RECT 132.735 107.525 135.235 107.755 ;
        RECT 134.790 107.425 135.220 107.525 ;
        RECT 132.730 106.465 133.240 106.585 ;
        RECT 132.730 106.235 135.235 106.465 ;
        RECT 132.730 106.115 133.240 106.235 ;
        RECT 134.790 105.175 135.220 105.285 ;
        RECT 132.735 104.945 135.235 105.175 ;
        RECT 134.790 104.845 135.220 104.945 ;
        RECT 132.730 103.885 133.240 104.025 ;
        RECT 132.730 103.655 135.235 103.885 ;
        RECT 132.730 103.555 133.240 103.655 ;
        RECT 134.790 102.595 135.220 102.705 ;
        RECT 132.735 102.365 135.235 102.595 ;
        RECT 134.790 102.265 135.220 102.365 ;
        RECT 132.720 101.305 133.230 101.435 ;
        RECT 132.720 101.075 135.235 101.305 ;
        RECT 132.720 100.965 133.230 101.075 ;
        RECT 134.790 100.015 135.220 100.125 ;
        RECT 132.735 99.785 135.235 100.015 ;
        RECT 134.790 99.685 135.220 99.785 ;
        RECT 132.740 98.725 133.250 98.855 ;
        RECT 132.735 98.495 135.235 98.725 ;
        RECT 132.740 98.385 133.250 98.495 ;
        RECT 134.790 97.435 135.220 97.545 ;
        RECT 132.735 97.205 135.235 97.435 ;
        RECT 134.790 97.105 135.220 97.205 ;
        RECT 132.730 96.145 133.240 96.265 ;
        RECT 132.730 95.915 135.235 96.145 ;
        RECT 132.730 95.795 133.240 95.915 ;
        RECT 134.790 94.855 135.220 94.965 ;
        RECT 132.735 94.625 135.235 94.855 ;
        RECT 134.790 94.525 135.220 94.625 ;
        RECT 132.730 93.565 133.240 93.695 ;
        RECT 132.730 93.335 135.235 93.565 ;
        RECT 132.730 93.225 133.240 93.335 ;
        RECT 134.790 92.275 135.220 92.385 ;
        RECT 132.735 92.045 135.235 92.275 ;
        RECT 134.790 91.945 135.220 92.045 ;
        RECT 132.740 90.985 133.250 91.115 ;
        RECT 132.735 90.755 135.235 90.985 ;
        RECT 132.740 90.645 133.250 90.755 ;
        RECT 134.790 89.695 135.220 89.805 ;
        RECT 132.735 89.465 135.235 89.695 ;
        RECT 134.790 89.365 135.220 89.465 ;
        RECT 132.720 88.405 133.230 88.525 ;
        RECT 132.720 88.175 135.235 88.405 ;
        RECT 132.720 88.055 133.230 88.175 ;
        RECT 134.790 87.115 135.220 87.215 ;
        RECT 132.735 86.885 135.235 87.115 ;
        RECT 134.790 86.775 135.220 86.885 ;
        RECT 132.730 85.825 133.240 85.945 ;
        RECT 132.730 85.595 135.235 85.825 ;
        RECT 132.730 85.475 133.240 85.595 ;
        RECT 134.790 84.535 135.220 84.635 ;
        RECT 132.735 84.305 135.235 84.535 ;
        RECT 134.790 84.195 135.220 84.305 ;
        RECT 132.740 83.245 133.250 83.365 ;
        RECT 132.735 83.015 135.235 83.245 ;
        RECT 132.740 82.895 133.250 83.015 ;
        RECT 134.790 81.955 135.220 82.055 ;
        RECT 132.735 81.725 135.235 81.955 ;
        RECT 134.790 81.615 135.220 81.725 ;
        RECT 135.430 80.155 135.680 107.535 ;
        RECT 135.980 80.155 136.230 107.535 ;
        RECT 136.415 107.525 138.930 107.755 ;
        RECT 138.500 107.425 138.930 107.525 ;
        RECT 136.440 106.465 136.950 106.595 ;
        RECT 136.415 106.235 138.915 106.465 ;
        RECT 136.440 106.125 136.950 106.235 ;
        RECT 138.500 105.175 138.930 105.285 ;
        RECT 136.415 104.945 138.930 105.175 ;
        RECT 138.500 104.845 138.930 104.945 ;
        RECT 136.440 103.885 136.950 104.015 ;
        RECT 136.415 103.655 138.915 103.885 ;
        RECT 136.440 103.545 136.950 103.655 ;
        RECT 138.500 102.595 138.930 102.705 ;
        RECT 136.415 102.365 138.930 102.595 ;
        RECT 138.500 102.265 138.930 102.365 ;
        RECT 136.440 101.305 136.950 101.415 ;
        RECT 136.415 101.075 138.915 101.305 ;
        RECT 136.440 100.945 136.950 101.075 ;
        RECT 138.500 100.015 138.930 100.125 ;
        RECT 136.415 99.785 138.930 100.015 ;
        RECT 138.500 99.685 138.930 99.785 ;
        RECT 136.440 98.725 136.950 98.855 ;
        RECT 136.415 98.495 138.915 98.725 ;
        RECT 136.440 98.385 136.950 98.495 ;
        RECT 138.500 97.435 138.930 97.545 ;
        RECT 136.415 97.205 138.930 97.435 ;
        RECT 138.500 97.105 138.930 97.205 ;
        RECT 136.440 96.145 136.950 96.265 ;
        RECT 136.415 95.915 138.915 96.145 ;
        RECT 136.440 95.795 136.950 95.915 ;
        RECT 138.500 94.855 138.930 94.965 ;
        RECT 136.415 94.625 138.930 94.855 ;
        RECT 138.500 94.525 138.930 94.625 ;
        RECT 136.440 93.565 136.950 93.705 ;
        RECT 136.415 93.335 138.915 93.565 ;
        RECT 136.440 93.235 136.950 93.335 ;
        RECT 138.500 92.275 138.930 92.385 ;
        RECT 136.415 92.045 138.930 92.275 ;
        RECT 138.500 91.945 138.930 92.045 ;
        RECT 136.440 90.985 136.950 91.105 ;
        RECT 136.415 90.755 138.915 90.985 ;
        RECT 136.440 90.635 136.950 90.755 ;
        RECT 138.500 89.695 138.930 89.805 ;
        RECT 136.415 89.465 138.930 89.695 ;
        RECT 138.500 89.365 138.930 89.465 ;
        RECT 136.440 88.405 136.950 88.515 ;
        RECT 136.415 88.175 138.915 88.405 ;
        RECT 136.440 88.045 136.950 88.175 ;
        RECT 138.500 87.115 138.930 87.225 ;
        RECT 136.415 86.885 138.930 87.115 ;
        RECT 138.500 86.785 138.930 86.885 ;
        RECT 136.440 85.825 136.950 85.945 ;
        RECT 136.415 85.595 138.915 85.825 ;
        RECT 136.440 85.475 136.950 85.595 ;
        RECT 138.500 84.535 138.930 84.645 ;
        RECT 136.415 84.305 138.930 84.535 ;
        RECT 138.500 84.205 138.930 84.305 ;
        RECT 136.440 83.245 136.950 83.365 ;
        RECT 136.415 83.015 138.915 83.245 ;
        RECT 136.440 82.895 136.950 83.015 ;
        RECT 138.500 81.955 138.930 82.065 ;
        RECT 136.415 81.725 138.930 81.955 ;
        RECT 138.500 81.625 138.930 81.725 ;
        RECT 139.110 80.155 139.360 107.535 ;
        RECT 139.660 80.155 139.910 107.535 ;
        RECT 140.095 107.525 142.595 107.755 ;
        RECT 142.140 107.425 142.570 107.525 ;
        RECT 140.110 106.465 140.620 106.595 ;
        RECT 140.095 106.235 142.595 106.465 ;
        RECT 140.110 106.125 140.620 106.235 ;
        RECT 142.140 105.175 142.570 105.285 ;
        RECT 140.095 104.945 142.595 105.175 ;
        RECT 142.140 104.845 142.570 104.945 ;
        RECT 140.110 103.885 140.620 104.015 ;
        RECT 140.095 103.655 142.595 103.885 ;
        RECT 140.110 103.545 140.620 103.655 ;
        RECT 142.140 102.595 142.570 102.695 ;
        RECT 140.095 102.365 142.595 102.595 ;
        RECT 142.140 102.255 142.570 102.365 ;
        RECT 140.110 101.305 140.620 101.415 ;
        RECT 140.095 101.075 142.595 101.305 ;
        RECT 140.110 100.945 140.620 101.075 ;
        RECT 142.140 100.015 142.570 100.125 ;
        RECT 140.095 99.785 142.595 100.015 ;
        RECT 142.140 99.685 142.570 99.785 ;
        RECT 140.110 98.725 140.620 98.855 ;
        RECT 140.095 98.495 142.595 98.725 ;
        RECT 140.110 98.385 140.620 98.495 ;
        RECT 142.140 97.435 142.570 97.545 ;
        RECT 140.095 97.205 142.595 97.435 ;
        RECT 142.140 97.105 142.570 97.205 ;
        RECT 140.110 96.145 140.620 96.265 ;
        RECT 140.095 95.915 142.595 96.145 ;
        RECT 140.110 95.795 140.620 95.915 ;
        RECT 142.140 94.855 142.570 94.965 ;
        RECT 140.095 94.625 142.595 94.855 ;
        RECT 142.140 94.525 142.570 94.625 ;
        RECT 140.110 93.565 140.620 93.695 ;
        RECT 140.095 93.335 142.595 93.565 ;
        RECT 140.110 93.225 140.620 93.335 ;
        RECT 142.140 92.275 142.570 92.385 ;
        RECT 140.095 92.045 142.595 92.275 ;
        RECT 142.140 91.945 142.570 92.045 ;
        RECT 140.110 90.985 140.620 91.105 ;
        RECT 140.095 90.755 142.595 90.985 ;
        RECT 140.110 90.635 140.620 90.755 ;
        RECT 142.150 89.695 142.580 89.805 ;
        RECT 140.095 89.465 142.595 89.695 ;
        RECT 142.150 89.365 142.580 89.465 ;
        RECT 140.110 88.405 140.620 88.515 ;
        RECT 140.095 88.175 142.595 88.405 ;
        RECT 140.110 88.045 140.620 88.175 ;
        RECT 142.150 87.115 142.580 87.225 ;
        RECT 140.095 86.885 142.595 87.115 ;
        RECT 142.150 86.785 142.580 86.885 ;
        RECT 140.110 85.825 140.620 85.935 ;
        RECT 140.095 85.595 142.595 85.825 ;
        RECT 140.110 85.465 140.620 85.595 ;
        RECT 142.150 84.535 142.580 84.645 ;
        RECT 140.095 84.305 142.595 84.535 ;
        RECT 142.150 84.205 142.580 84.305 ;
        RECT 140.110 83.245 140.620 83.355 ;
        RECT 140.095 83.015 142.595 83.245 ;
        RECT 140.110 82.885 140.620 83.015 ;
        RECT 142.150 81.955 142.580 82.055 ;
        RECT 140.095 81.725 142.595 81.955 ;
        RECT 142.150 81.615 142.580 81.725 ;
        RECT 142.780 80.155 143.030 107.535 ;
        RECT 143.330 80.155 143.580 107.535 ;
        RECT 143.775 107.525 146.275 107.755 ;
        RECT 145.830 107.425 146.260 107.525 ;
        RECT 143.790 106.465 144.300 106.585 ;
        RECT 143.775 106.235 146.275 106.465 ;
        RECT 143.790 106.115 144.300 106.235 ;
        RECT 145.830 105.175 146.260 105.275 ;
        RECT 143.775 104.945 146.275 105.175 ;
        RECT 145.830 104.835 146.260 104.945 ;
        RECT 143.790 103.885 144.300 104.005 ;
        RECT 143.775 103.655 146.275 103.885 ;
        RECT 143.790 103.535 144.300 103.655 ;
        RECT 145.830 102.595 146.260 102.695 ;
        RECT 143.775 102.365 146.275 102.595 ;
        RECT 145.830 102.255 146.260 102.365 ;
        RECT 143.790 101.305 144.300 101.425 ;
        RECT 143.775 101.075 146.275 101.305 ;
        RECT 143.790 100.955 144.300 101.075 ;
        RECT 145.830 100.015 146.260 100.115 ;
        RECT 143.775 99.785 146.275 100.015 ;
        RECT 145.830 99.675 146.260 99.785 ;
        RECT 143.790 98.725 144.300 98.845 ;
        RECT 143.775 98.495 146.275 98.725 ;
        RECT 143.790 98.375 144.300 98.495 ;
        RECT 145.830 97.435 146.260 97.535 ;
        RECT 143.775 97.205 146.275 97.435 ;
        RECT 145.830 97.095 146.260 97.205 ;
        RECT 143.790 96.145 144.300 96.265 ;
        RECT 143.775 95.915 146.275 96.145 ;
        RECT 143.790 95.795 144.300 95.915 ;
        RECT 145.830 94.855 146.260 94.955 ;
        RECT 143.775 94.625 146.275 94.855 ;
        RECT 145.830 94.515 146.260 94.625 ;
        RECT 143.790 93.565 144.300 93.685 ;
        RECT 143.775 93.335 146.275 93.565 ;
        RECT 143.790 93.215 144.300 93.335 ;
        RECT 145.830 92.275 146.260 92.375 ;
        RECT 143.775 92.045 146.275 92.275 ;
        RECT 145.830 91.935 146.260 92.045 ;
        RECT 143.790 90.985 144.300 91.115 ;
        RECT 143.775 90.755 146.275 90.985 ;
        RECT 143.790 90.645 144.300 90.755 ;
        RECT 145.830 89.695 146.260 89.795 ;
        RECT 143.775 89.465 146.275 89.695 ;
        RECT 145.830 89.355 146.260 89.465 ;
        RECT 143.800 88.405 144.310 88.525 ;
        RECT 143.775 88.175 146.275 88.405 ;
        RECT 143.800 88.055 144.310 88.175 ;
        RECT 145.830 87.115 146.260 87.225 ;
        RECT 143.775 86.885 146.275 87.115 ;
        RECT 145.830 86.785 146.260 86.885 ;
        RECT 143.800 85.825 144.310 85.945 ;
        RECT 143.775 85.595 146.275 85.825 ;
        RECT 143.800 85.475 144.310 85.595 ;
        RECT 145.830 84.535 146.260 84.635 ;
        RECT 143.775 84.305 146.275 84.535 ;
        RECT 145.830 84.195 146.260 84.305 ;
        RECT 143.820 83.245 144.330 83.355 ;
        RECT 143.775 83.015 146.275 83.245 ;
        RECT 143.820 82.885 144.330 83.015 ;
        RECT 145.830 81.955 146.260 82.055 ;
        RECT 143.775 81.725 146.275 81.955 ;
        RECT 145.830 81.615 146.260 81.725 ;
        RECT 146.470 80.155 146.720 107.545 ;
        RECT 149.010 106.595 151.240 110.240 ;
        RECT 146.880 104.575 151.240 106.595 ;
        RECT 149.010 85.715 151.240 104.575 ;
        RECT 146.870 83.695 151.240 85.715 ;
        RECT 117.880 79.075 146.720 80.155 ;
        RECT 147.450 79.950 148.125 79.980 ;
        RECT 149.010 79.950 151.240 83.695 ;
        RECT 147.450 79.275 151.240 79.950 ;
        RECT 147.450 79.245 148.125 79.275 ;
        RECT 117.880 79.045 118.960 79.075 ;
        RECT 110.575 62.345 113.635 62.765 ;
        RECT 108.170 62.115 113.635 62.345 ;
        RECT 102.660 55.985 108.010 57.715 ;
        RECT 102.660 55.975 107.530 55.985 ;
        RECT 102.680 43.655 104.910 55.975 ;
        RECT 102.680 41.915 108.010 43.655 ;
        RECT 102.680 36.935 104.910 41.915 ;
        RECT 108.170 38.545 108.400 62.115 ;
        RECT 108.570 61.515 108.910 61.635 ;
        RECT 108.560 61.285 109.560 61.515 ;
        RECT 108.570 61.175 108.910 61.285 ;
        RECT 109.200 59.225 109.520 59.345 ;
        RECT 108.560 58.995 109.560 59.225 ;
        RECT 109.200 58.885 109.520 58.995 ;
        RECT 108.570 56.935 108.910 57.045 ;
        RECT 108.560 56.705 109.560 56.935 ;
        RECT 108.570 56.585 108.910 56.705 ;
        RECT 109.200 54.645 109.520 54.775 ;
        RECT 108.560 54.415 109.560 54.645 ;
        RECT 109.200 54.315 109.520 54.415 ;
        RECT 108.570 52.355 108.910 52.485 ;
        RECT 108.560 52.125 109.560 52.355 ;
        RECT 108.570 52.025 108.910 52.125 ;
        RECT 109.200 50.065 109.520 50.185 ;
        RECT 108.560 49.835 109.560 50.065 ;
        RECT 109.200 49.725 109.520 49.835 ;
        RECT 108.570 47.775 108.910 47.905 ;
        RECT 108.560 47.545 109.560 47.775 ;
        RECT 108.570 47.445 108.910 47.545 ;
        RECT 109.200 45.485 109.520 45.605 ;
        RECT 108.560 45.255 109.560 45.485 ;
        RECT 109.200 45.145 109.520 45.255 ;
        RECT 108.570 43.195 108.910 43.315 ;
        RECT 108.560 42.965 109.560 43.195 ;
        RECT 108.570 42.855 108.910 42.965 ;
        RECT 109.200 40.905 109.520 41.025 ;
        RECT 108.560 40.675 109.560 40.905 ;
        RECT 109.200 40.565 109.520 40.675 ;
        RECT 108.570 38.615 108.910 38.735 ;
        RECT 108.560 38.385 109.560 38.615 ;
        RECT 109.720 38.545 109.950 62.115 ;
        RECT 110.575 61.690 113.635 62.115 ;
        RECT 110.825 52.300 111.935 53.350 ;
        RECT 110.855 49.550 111.905 52.300 ;
        RECT 112.560 49.880 113.635 61.690 ;
        RECT 111.075 47.755 111.665 49.550 ;
        RECT 112.555 48.870 114.710 49.880 ;
        RECT 111.075 43.235 111.670 47.755 ;
        RECT 113.700 45.615 114.710 48.870 ;
        RECT 113.250 45.605 114.710 45.615 ;
        RECT 113.250 45.335 115.090 45.605 ;
        RECT 111.075 39.595 113.040 43.235 ;
        RECT 108.570 38.275 108.910 38.385 ;
        RECT 111.075 38.145 111.665 39.595 ;
        RECT 113.250 39.165 113.520 45.335 ;
        RECT 113.720 43.815 114.050 43.935 ;
        RECT 113.670 43.585 114.670 43.815 ;
        RECT 113.720 43.475 114.050 43.585 ;
        RECT 114.280 41.525 114.610 41.645 ;
        RECT 113.670 41.295 114.670 41.525 ;
        RECT 114.280 41.195 114.610 41.295 ;
        RECT 113.720 39.235 114.050 39.345 ;
        RECT 113.670 39.005 114.670 39.235 ;
        RECT 114.820 39.165 115.090 45.335 ;
        RECT 116.730 43.665 117.780 53.380 ;
        RECT 121.250 51.545 121.500 79.075 ;
        RECT 123.770 77.395 124.200 77.505 ;
        RECT 121.695 77.165 124.200 77.395 ;
        RECT 123.770 77.065 124.200 77.165 ;
        RECT 121.680 76.105 122.200 76.255 ;
        RECT 121.680 75.875 124.195 76.105 ;
        RECT 121.680 75.755 122.200 75.875 ;
        RECT 123.770 74.815 124.200 74.915 ;
        RECT 121.695 74.585 124.200 74.815 ;
        RECT 123.770 74.475 124.200 74.585 ;
        RECT 121.680 73.525 122.200 73.665 ;
        RECT 121.680 73.295 124.195 73.525 ;
        RECT 121.680 73.165 122.200 73.295 ;
        RECT 123.770 72.235 124.200 72.345 ;
        RECT 121.695 72.005 124.200 72.235 ;
        RECT 123.770 71.905 124.200 72.005 ;
        RECT 121.670 70.945 122.190 71.075 ;
        RECT 121.670 70.715 124.195 70.945 ;
        RECT 121.670 70.575 122.190 70.715 ;
        RECT 123.770 69.655 124.200 69.765 ;
        RECT 121.695 69.425 124.200 69.655 ;
        RECT 123.770 69.325 124.200 69.425 ;
        RECT 121.690 68.365 122.210 68.505 ;
        RECT 121.690 68.135 124.195 68.365 ;
        RECT 121.690 68.005 122.210 68.135 ;
        RECT 123.770 67.075 124.200 67.185 ;
        RECT 121.695 66.845 124.200 67.075 ;
        RECT 123.770 66.745 124.200 66.845 ;
        RECT 121.700 65.785 122.220 65.925 ;
        RECT 121.695 65.555 124.195 65.785 ;
        RECT 121.700 65.425 122.220 65.555 ;
        RECT 123.770 64.495 124.200 64.605 ;
        RECT 121.695 64.265 124.200 64.495 ;
        RECT 123.770 64.165 124.200 64.265 ;
        RECT 121.680 63.205 122.200 63.345 ;
        RECT 121.680 62.975 124.195 63.205 ;
        RECT 121.680 62.845 122.200 62.975 ;
        RECT 123.770 61.915 124.200 62.025 ;
        RECT 121.695 61.685 124.200 61.915 ;
        RECT 123.770 61.585 124.200 61.685 ;
        RECT 121.690 60.625 122.210 60.745 ;
        RECT 121.690 60.395 124.195 60.625 ;
        RECT 121.690 60.245 122.210 60.395 ;
        RECT 123.770 59.335 124.200 59.445 ;
        RECT 121.695 59.105 124.200 59.335 ;
        RECT 123.770 59.005 124.200 59.105 ;
        RECT 121.690 58.045 122.210 58.185 ;
        RECT 121.690 57.815 124.195 58.045 ;
        RECT 121.690 57.685 122.210 57.815 ;
        RECT 123.770 56.755 124.200 56.865 ;
        RECT 121.695 56.525 124.200 56.755 ;
        RECT 123.770 56.425 124.200 56.525 ;
        RECT 121.700 55.465 122.220 55.595 ;
        RECT 121.695 55.235 124.195 55.465 ;
        RECT 121.700 55.095 122.220 55.235 ;
        RECT 123.770 54.175 124.200 54.285 ;
        RECT 121.695 53.945 124.200 54.175 ;
        RECT 123.770 53.845 124.200 53.945 ;
        RECT 121.700 52.885 122.220 53.015 ;
        RECT 121.695 52.655 124.195 52.885 ;
        RECT 121.700 52.515 122.220 52.655 ;
        RECT 123.770 51.595 124.200 51.705 ;
        RECT 121.695 51.365 124.200 51.595 ;
        RECT 124.400 51.545 124.650 79.075 ;
        RECT 124.940 51.555 125.190 79.075 ;
        RECT 127.400 77.395 127.830 77.505 ;
        RECT 125.375 77.165 127.875 77.395 ;
        RECT 127.400 77.065 127.830 77.165 ;
        RECT 125.370 76.105 125.890 76.245 ;
        RECT 125.370 75.875 127.875 76.105 ;
        RECT 125.370 75.745 125.890 75.875 ;
        RECT 127.410 74.815 127.840 74.925 ;
        RECT 125.375 74.585 127.875 74.815 ;
        RECT 127.410 74.485 127.840 74.585 ;
        RECT 125.350 73.525 125.870 73.655 ;
        RECT 125.350 73.295 127.875 73.525 ;
        RECT 125.350 73.155 125.870 73.295 ;
        RECT 127.410 72.235 127.840 72.345 ;
        RECT 125.375 72.005 127.875 72.235 ;
        RECT 127.410 71.905 127.840 72.005 ;
        RECT 125.370 70.945 125.890 71.085 ;
        RECT 125.370 70.715 127.875 70.945 ;
        RECT 125.370 70.585 125.890 70.715 ;
        RECT 127.410 69.655 127.840 69.765 ;
        RECT 125.375 69.425 127.875 69.655 ;
        RECT 127.410 69.325 127.840 69.425 ;
        RECT 125.370 68.365 125.890 68.505 ;
        RECT 125.370 68.135 127.875 68.365 ;
        RECT 125.370 68.005 125.890 68.135 ;
        RECT 127.410 67.075 127.840 67.185 ;
        RECT 125.375 66.845 127.875 67.075 ;
        RECT 127.410 66.745 127.840 66.845 ;
        RECT 125.350 65.785 125.870 65.915 ;
        RECT 125.350 65.555 127.875 65.785 ;
        RECT 125.350 65.415 125.870 65.555 ;
        RECT 127.410 64.495 127.840 64.605 ;
        RECT 125.375 64.265 127.875 64.495 ;
        RECT 127.410 64.165 127.840 64.265 ;
        RECT 125.370 63.205 125.890 63.335 ;
        RECT 125.370 62.975 127.875 63.205 ;
        RECT 125.370 62.835 125.890 62.975 ;
        RECT 127.410 61.915 127.840 62.025 ;
        RECT 125.375 61.685 127.875 61.915 ;
        RECT 127.410 61.585 127.840 61.685 ;
        RECT 125.390 60.625 125.910 60.755 ;
        RECT 125.375 60.395 127.875 60.625 ;
        RECT 125.390 60.255 125.910 60.395 ;
        RECT 127.410 59.335 127.840 59.445 ;
        RECT 125.375 59.105 127.875 59.335 ;
        RECT 127.410 59.005 127.840 59.105 ;
        RECT 125.370 58.045 125.890 58.185 ;
        RECT 125.370 57.815 127.875 58.045 ;
        RECT 125.370 57.685 125.890 57.815 ;
        RECT 127.410 56.755 127.840 56.865 ;
        RECT 125.375 56.525 127.875 56.755 ;
        RECT 127.410 56.425 127.840 56.525 ;
        RECT 125.380 55.465 125.900 55.605 ;
        RECT 125.375 55.235 127.875 55.465 ;
        RECT 125.380 55.105 125.900 55.235 ;
        RECT 127.410 54.175 127.840 54.285 ;
        RECT 125.375 53.945 127.875 54.175 ;
        RECT 127.410 53.845 127.840 53.945 ;
        RECT 125.370 52.885 125.890 53.025 ;
        RECT 125.370 52.655 127.875 52.885 ;
        RECT 125.370 52.525 125.890 52.655 ;
        RECT 127.410 51.595 127.840 51.705 ;
        RECT 125.375 51.365 127.875 51.595 ;
        RECT 128.080 51.545 128.330 79.075 ;
        RECT 128.620 51.545 128.870 79.075 ;
        RECT 131.150 77.395 131.580 77.505 ;
        RECT 129.055 77.165 131.580 77.395 ;
        RECT 131.150 77.065 131.580 77.165 ;
        RECT 129.060 76.105 129.580 76.245 ;
        RECT 129.055 75.875 131.555 76.105 ;
        RECT 129.060 75.745 129.580 75.875 ;
        RECT 131.150 74.815 131.580 74.935 ;
        RECT 129.055 74.585 131.580 74.815 ;
        RECT 131.150 74.495 131.580 74.585 ;
        RECT 129.040 73.525 129.560 73.655 ;
        RECT 129.040 73.295 131.555 73.525 ;
        RECT 129.040 73.155 129.560 73.295 ;
        RECT 131.150 72.235 131.580 72.345 ;
        RECT 129.055 72.005 131.580 72.235 ;
        RECT 131.150 71.905 131.580 72.005 ;
        RECT 129.060 70.945 129.580 71.075 ;
        RECT 129.055 70.715 131.555 70.945 ;
        RECT 129.060 70.575 129.580 70.715 ;
        RECT 131.150 69.655 131.580 69.765 ;
        RECT 129.055 69.425 131.580 69.655 ;
        RECT 131.150 69.325 131.580 69.425 ;
        RECT 129.050 68.365 129.570 68.495 ;
        RECT 129.050 68.135 131.555 68.365 ;
        RECT 129.050 67.995 129.570 68.135 ;
        RECT 131.150 67.075 131.580 67.185 ;
        RECT 129.055 66.845 131.580 67.075 ;
        RECT 131.150 66.745 131.580 66.845 ;
        RECT 129.050 65.785 129.570 65.935 ;
        RECT 129.050 65.555 131.555 65.785 ;
        RECT 129.050 65.435 129.570 65.555 ;
        RECT 131.150 64.495 131.580 64.595 ;
        RECT 129.055 64.265 131.580 64.495 ;
        RECT 131.150 64.155 131.580 64.265 ;
        RECT 129.050 63.205 129.570 63.335 ;
        RECT 129.050 62.975 131.555 63.205 ;
        RECT 129.050 62.835 129.570 62.975 ;
        RECT 131.150 61.915 131.580 62.035 ;
        RECT 129.055 61.685 131.580 61.915 ;
        RECT 131.150 61.595 131.580 61.685 ;
        RECT 129.060 60.625 129.580 60.755 ;
        RECT 129.055 60.395 131.555 60.625 ;
        RECT 129.060 60.255 129.580 60.395 ;
        RECT 131.150 59.335 131.580 59.445 ;
        RECT 129.055 59.105 131.580 59.335 ;
        RECT 131.150 59.005 131.580 59.105 ;
        RECT 129.040 58.045 129.560 58.195 ;
        RECT 129.040 57.815 131.555 58.045 ;
        RECT 129.040 57.695 129.560 57.815 ;
        RECT 131.150 56.755 131.580 56.875 ;
        RECT 129.055 56.525 131.580 56.755 ;
        RECT 131.150 56.435 131.580 56.525 ;
        RECT 129.050 55.465 129.570 55.595 ;
        RECT 129.050 55.235 131.555 55.465 ;
        RECT 129.050 55.095 129.570 55.235 ;
        RECT 131.150 54.175 131.580 54.285 ;
        RECT 129.055 53.945 131.580 54.175 ;
        RECT 131.150 53.845 131.580 53.945 ;
        RECT 129.050 52.885 129.570 53.035 ;
        RECT 129.050 52.655 131.555 52.885 ;
        RECT 129.050 52.535 129.570 52.655 ;
        RECT 131.150 51.595 131.580 51.705 ;
        RECT 129.055 51.365 131.580 51.595 ;
        RECT 131.750 51.545 132.000 79.075 ;
        RECT 132.300 51.545 132.550 79.075 ;
        RECT 134.790 77.395 135.220 77.505 ;
        RECT 132.735 77.165 135.235 77.395 ;
        RECT 134.790 77.065 135.220 77.165 ;
        RECT 132.740 76.105 133.260 76.245 ;
        RECT 132.735 75.875 135.235 76.105 ;
        RECT 132.740 75.745 133.260 75.875 ;
        RECT 134.790 74.815 135.220 74.925 ;
        RECT 132.735 74.585 135.235 74.815 ;
        RECT 134.790 74.485 135.220 74.585 ;
        RECT 132.740 73.525 133.260 73.655 ;
        RECT 132.735 73.295 135.235 73.525 ;
        RECT 132.740 73.155 133.260 73.295 ;
        RECT 134.790 72.235 135.220 72.345 ;
        RECT 132.735 72.005 135.235 72.235 ;
        RECT 134.790 71.905 135.220 72.005 ;
        RECT 132.740 70.945 133.260 71.085 ;
        RECT 132.735 70.715 135.235 70.945 ;
        RECT 132.740 70.585 133.260 70.715 ;
        RECT 134.790 69.655 135.220 69.765 ;
        RECT 132.735 69.425 135.235 69.655 ;
        RECT 134.790 69.325 135.220 69.425 ;
        RECT 132.740 68.365 133.260 68.495 ;
        RECT 132.735 68.135 135.235 68.365 ;
        RECT 132.740 67.995 133.260 68.135 ;
        RECT 134.790 67.075 135.220 67.185 ;
        RECT 132.735 66.845 135.235 67.075 ;
        RECT 134.790 66.745 135.220 66.845 ;
        RECT 132.740 65.785 133.260 65.935 ;
        RECT 132.735 65.555 135.235 65.785 ;
        RECT 132.740 65.435 133.260 65.555 ;
        RECT 134.790 64.495 135.220 64.605 ;
        RECT 132.735 64.265 135.235 64.495 ;
        RECT 134.790 64.165 135.220 64.265 ;
        RECT 132.730 63.205 133.250 63.335 ;
        RECT 132.730 62.975 135.235 63.205 ;
        RECT 132.730 62.835 133.250 62.975 ;
        RECT 134.790 61.915 135.220 62.025 ;
        RECT 132.735 61.685 135.235 61.915 ;
        RECT 134.790 61.585 135.220 61.685 ;
        RECT 132.740 60.625 133.260 60.755 ;
        RECT 132.735 60.395 135.235 60.625 ;
        RECT 132.740 60.255 133.260 60.395 ;
        RECT 134.790 59.335 135.220 59.445 ;
        RECT 132.735 59.105 135.235 59.335 ;
        RECT 134.790 59.005 135.220 59.105 ;
        RECT 132.740 58.045 133.260 58.165 ;
        RECT 132.735 57.815 135.235 58.045 ;
        RECT 132.740 57.665 133.260 57.815 ;
        RECT 134.790 56.755 135.220 56.865 ;
        RECT 132.735 56.525 135.235 56.755 ;
        RECT 134.790 56.425 135.220 56.525 ;
        RECT 132.740 55.465 133.260 55.595 ;
        RECT 132.735 55.235 135.235 55.465 ;
        RECT 132.740 55.095 133.260 55.235 ;
        RECT 134.790 54.175 135.220 54.285 ;
        RECT 132.735 53.945 135.235 54.175 ;
        RECT 134.790 53.845 135.220 53.945 ;
        RECT 132.740 52.885 133.260 53.025 ;
        RECT 132.735 52.655 135.235 52.885 ;
        RECT 132.740 52.525 133.260 52.655 ;
        RECT 134.790 51.595 135.220 51.695 ;
        RECT 132.735 51.365 135.235 51.595 ;
        RECT 135.430 51.545 135.680 79.075 ;
        RECT 135.980 51.545 136.230 79.075 ;
        RECT 138.490 77.395 138.920 77.495 ;
        RECT 136.415 77.165 138.920 77.395 ;
        RECT 138.490 77.055 138.920 77.165 ;
        RECT 136.410 76.105 136.930 76.245 ;
        RECT 136.410 75.875 138.915 76.105 ;
        RECT 136.410 75.745 136.930 75.875 ;
        RECT 138.490 74.815 138.920 74.935 ;
        RECT 136.415 74.585 138.920 74.815 ;
        RECT 138.490 74.495 138.920 74.585 ;
        RECT 136.400 73.525 136.920 73.665 ;
        RECT 136.400 73.295 138.915 73.525 ;
        RECT 136.400 73.165 136.920 73.295 ;
        RECT 138.490 72.235 138.920 72.345 ;
        RECT 136.415 72.005 138.920 72.235 ;
        RECT 138.490 71.905 138.920 72.005 ;
        RECT 136.410 70.945 136.930 71.075 ;
        RECT 136.410 70.715 138.915 70.945 ;
        RECT 136.410 70.575 136.930 70.715 ;
        RECT 138.490 69.655 138.920 69.765 ;
        RECT 136.415 69.425 138.920 69.655 ;
        RECT 138.490 69.325 138.920 69.425 ;
        RECT 136.400 68.365 136.920 68.495 ;
        RECT 136.400 68.135 138.915 68.365 ;
        RECT 136.400 67.995 136.920 68.135 ;
        RECT 138.490 67.075 138.920 67.185 ;
        RECT 136.415 66.845 138.920 67.075 ;
        RECT 138.490 66.745 138.920 66.845 ;
        RECT 136.400 65.785 136.920 65.915 ;
        RECT 136.400 65.555 138.915 65.785 ;
        RECT 136.400 65.415 136.920 65.555 ;
        RECT 138.490 64.495 138.920 64.605 ;
        RECT 136.415 64.265 138.920 64.495 ;
        RECT 138.490 64.165 138.920 64.265 ;
        RECT 136.410 63.205 136.930 63.325 ;
        RECT 136.410 62.975 138.915 63.205 ;
        RECT 136.410 62.825 136.930 62.975 ;
        RECT 138.490 61.915 138.920 62.025 ;
        RECT 136.415 61.685 138.920 61.915 ;
        RECT 138.490 61.585 138.920 61.685 ;
        RECT 136.420 60.625 136.940 60.755 ;
        RECT 136.415 60.395 138.915 60.625 ;
        RECT 136.420 60.255 136.940 60.395 ;
        RECT 138.490 59.335 138.920 59.445 ;
        RECT 136.415 59.105 138.920 59.335 ;
        RECT 138.490 59.005 138.920 59.105 ;
        RECT 136.420 58.045 136.940 58.185 ;
        RECT 136.415 57.815 138.915 58.045 ;
        RECT 136.420 57.685 136.940 57.815 ;
        RECT 138.490 56.755 138.920 56.865 ;
        RECT 136.415 56.525 138.920 56.755 ;
        RECT 138.490 56.425 138.920 56.525 ;
        RECT 136.410 55.465 136.930 55.605 ;
        RECT 136.410 55.235 138.915 55.465 ;
        RECT 136.410 55.105 136.930 55.235 ;
        RECT 138.490 54.175 138.920 54.285 ;
        RECT 136.415 53.945 138.920 54.175 ;
        RECT 138.490 53.845 138.920 53.945 ;
        RECT 136.420 52.885 136.940 53.015 ;
        RECT 136.415 52.655 138.915 52.885 ;
        RECT 136.420 52.515 136.940 52.655 ;
        RECT 138.490 51.595 138.920 51.705 ;
        RECT 136.415 51.365 138.920 51.595 ;
        RECT 139.110 51.545 139.360 79.075 ;
        RECT 139.660 51.545 139.910 79.075 ;
        RECT 142.150 77.395 142.580 77.495 ;
        RECT 140.095 77.165 142.595 77.395 ;
        RECT 142.150 77.055 142.580 77.165 ;
        RECT 140.100 76.105 140.620 76.245 ;
        RECT 140.095 75.875 142.595 76.105 ;
        RECT 140.100 75.745 140.620 75.875 ;
        RECT 142.150 74.815 142.580 74.925 ;
        RECT 140.095 74.585 142.595 74.815 ;
        RECT 142.150 74.485 142.580 74.585 ;
        RECT 140.080 73.525 140.600 73.655 ;
        RECT 140.080 73.295 142.595 73.525 ;
        RECT 140.080 73.155 140.600 73.295 ;
        RECT 142.150 72.235 142.580 72.345 ;
        RECT 140.095 72.005 142.595 72.235 ;
        RECT 142.150 71.905 142.580 72.005 ;
        RECT 140.090 70.945 140.610 71.075 ;
        RECT 140.090 70.715 142.595 70.945 ;
        RECT 140.090 70.575 140.610 70.715 ;
        RECT 142.150 69.655 142.580 69.755 ;
        RECT 140.095 69.425 142.595 69.655 ;
        RECT 142.150 69.315 142.580 69.425 ;
        RECT 140.080 68.365 140.600 68.495 ;
        RECT 140.080 68.135 142.595 68.365 ;
        RECT 140.080 67.995 140.600 68.135 ;
        RECT 142.150 67.075 142.580 67.195 ;
        RECT 140.095 66.845 142.595 67.075 ;
        RECT 142.150 66.755 142.580 66.845 ;
        RECT 140.110 65.785 140.630 65.905 ;
        RECT 140.095 65.555 142.595 65.785 ;
        RECT 140.110 65.405 140.630 65.555 ;
        RECT 142.130 64.495 142.560 64.605 ;
        RECT 140.095 64.265 142.595 64.495 ;
        RECT 142.130 64.165 142.560 64.265 ;
        RECT 140.090 63.205 140.610 63.335 ;
        RECT 140.090 62.975 142.595 63.205 ;
        RECT 140.090 62.835 140.610 62.975 ;
        RECT 142.130 61.915 142.560 62.025 ;
        RECT 140.095 61.685 142.595 61.915 ;
        RECT 142.130 61.585 142.560 61.685 ;
        RECT 140.080 60.625 140.600 60.755 ;
        RECT 140.080 60.395 142.595 60.625 ;
        RECT 140.080 60.255 140.600 60.395 ;
        RECT 142.130 59.335 142.560 59.455 ;
        RECT 140.095 59.105 142.595 59.335 ;
        RECT 142.130 59.015 142.560 59.105 ;
        RECT 140.100 58.045 140.620 58.175 ;
        RECT 140.095 57.815 142.595 58.045 ;
        RECT 140.100 57.675 140.620 57.815 ;
        RECT 142.130 56.755 142.560 56.865 ;
        RECT 140.095 56.525 142.595 56.755 ;
        RECT 142.130 56.425 142.560 56.525 ;
        RECT 140.100 55.465 140.620 55.605 ;
        RECT 140.095 55.235 142.595 55.465 ;
        RECT 140.100 55.105 140.620 55.235 ;
        RECT 142.130 54.175 142.560 54.275 ;
        RECT 140.095 53.945 142.595 54.175 ;
        RECT 142.130 53.835 142.560 53.945 ;
        RECT 140.100 52.885 140.620 53.015 ;
        RECT 140.095 52.655 142.595 52.885 ;
        RECT 140.100 52.515 140.620 52.655 ;
        RECT 142.130 51.595 142.560 51.695 ;
        RECT 140.095 51.365 142.595 51.595 ;
        RECT 142.780 51.545 143.030 79.075 ;
        RECT 143.330 51.545 143.580 79.075 ;
        RECT 145.830 77.395 146.260 77.495 ;
        RECT 143.775 77.165 146.275 77.395 ;
        RECT 145.830 77.055 146.260 77.165 ;
        RECT 143.780 76.105 144.300 76.255 ;
        RECT 143.775 75.875 146.275 76.105 ;
        RECT 143.780 75.755 144.300 75.875 ;
        RECT 145.830 74.815 146.260 74.925 ;
        RECT 143.775 74.585 146.275 74.815 ;
        RECT 145.830 74.485 146.260 74.585 ;
        RECT 143.780 73.525 144.300 73.655 ;
        RECT 143.775 73.295 146.275 73.525 ;
        RECT 143.780 73.155 144.300 73.295 ;
        RECT 145.830 72.235 146.260 72.345 ;
        RECT 143.775 72.005 146.275 72.235 ;
        RECT 145.830 71.905 146.260 72.005 ;
        RECT 143.780 70.945 144.300 71.065 ;
        RECT 143.775 70.715 146.275 70.945 ;
        RECT 143.780 70.565 144.300 70.715 ;
        RECT 145.830 69.655 146.260 69.765 ;
        RECT 143.775 69.425 146.275 69.655 ;
        RECT 145.830 69.325 146.260 69.425 ;
        RECT 143.760 68.365 144.280 68.485 ;
        RECT 143.760 68.135 146.275 68.365 ;
        RECT 143.760 67.985 144.280 68.135 ;
        RECT 145.830 67.075 146.260 67.175 ;
        RECT 143.775 66.845 146.275 67.075 ;
        RECT 145.830 66.735 146.260 66.845 ;
        RECT 143.780 65.785 144.300 65.915 ;
        RECT 143.775 65.555 146.275 65.785 ;
        RECT 143.780 65.415 144.300 65.555 ;
        RECT 145.830 64.495 146.260 64.605 ;
        RECT 143.775 64.265 146.275 64.495 ;
        RECT 145.830 64.165 146.260 64.265 ;
        RECT 143.790 63.205 144.310 63.335 ;
        RECT 143.775 62.975 146.275 63.205 ;
        RECT 143.790 62.835 144.310 62.975 ;
        RECT 145.830 61.915 146.260 62.015 ;
        RECT 143.775 61.685 146.275 61.915 ;
        RECT 145.830 61.575 146.260 61.685 ;
        RECT 143.790 60.625 144.310 60.765 ;
        RECT 143.775 60.395 146.275 60.625 ;
        RECT 143.790 60.265 144.310 60.395 ;
        RECT 145.830 59.335 146.260 59.445 ;
        RECT 143.775 59.105 146.275 59.335 ;
        RECT 145.830 59.005 146.260 59.105 ;
        RECT 143.780 58.045 144.300 58.165 ;
        RECT 143.775 57.815 146.275 58.045 ;
        RECT 143.780 57.665 144.300 57.815 ;
        RECT 145.830 56.755 146.260 56.855 ;
        RECT 143.775 56.525 146.275 56.755 ;
        RECT 145.830 56.415 146.260 56.525 ;
        RECT 143.770 55.465 144.290 55.585 ;
        RECT 143.770 55.235 146.275 55.465 ;
        RECT 143.770 55.085 144.290 55.235 ;
        RECT 145.830 54.175 146.260 54.285 ;
        RECT 143.775 53.945 146.275 54.175 ;
        RECT 145.830 53.845 146.260 53.945 ;
        RECT 143.780 52.885 144.300 53.015 ;
        RECT 143.775 52.655 146.275 52.885 ;
        RECT 143.780 52.515 144.300 52.655 ;
        RECT 145.830 51.595 146.260 51.695 ;
        RECT 143.775 51.365 146.275 51.595 ;
        RECT 146.470 51.555 146.720 79.075 ;
        RECT 149.010 76.245 151.240 79.275 ;
        RECT 146.890 74.225 151.240 76.245 ;
        RECT 149.010 55.415 151.240 74.225 ;
        RECT 146.880 53.395 151.240 55.415 ;
        RECT 123.770 51.265 124.200 51.365 ;
        RECT 127.410 51.265 127.840 51.365 ;
        RECT 131.150 51.265 131.580 51.365 ;
        RECT 134.790 51.255 135.220 51.365 ;
        RECT 138.490 51.265 138.920 51.365 ;
        RECT 142.130 51.255 142.560 51.365 ;
        RECT 145.830 51.255 146.260 51.365 ;
        RECT 131.150 45.895 131.880 48.710 ;
        RECT 129.190 45.815 131.880 45.895 ;
        RECT 140.555 47.860 146.430 48.090 ;
        RECT 140.555 45.835 140.785 47.860 ;
        RECT 141.310 47.280 141.965 47.310 ;
        RECT 143.590 47.280 144.245 47.860 ;
        RECT 141.310 47.245 144.245 47.280 ;
        RECT 141.310 46.625 144.250 47.245 ;
        RECT 141.310 46.595 141.965 46.625 ;
        RECT 143.700 46.085 144.250 46.625 ;
        RECT 141.060 46.025 145.940 46.085 ;
        RECT 122.860 45.185 123.140 45.195 ;
        RECT 123.380 45.185 123.660 45.195 ;
        RECT 127.940 45.185 128.220 45.715 ;
        RECT 118.280 44.905 128.220 45.185 ;
        RECT 116.730 39.335 118.070 43.665 ;
        RECT 118.280 39.515 118.560 44.905 ;
        RECT 118.770 43.995 119.190 44.095 ;
        RECT 118.710 43.765 122.710 43.995 ;
        RECT 118.770 43.675 119.190 43.765 ;
        RECT 122.220 43.515 122.640 43.605 ;
        RECT 118.710 43.285 122.710 43.515 ;
        RECT 122.220 43.185 122.640 43.285 ;
        RECT 118.770 43.035 119.190 43.135 ;
        RECT 118.710 42.805 122.710 43.035 ;
        RECT 118.770 42.715 119.190 42.805 ;
        RECT 122.220 42.555 122.640 42.655 ;
        RECT 118.710 42.325 122.710 42.555 ;
        RECT 122.220 42.235 122.640 42.325 ;
        RECT 118.770 42.075 119.190 42.175 ;
        RECT 118.710 41.845 122.710 42.075 ;
        RECT 118.770 41.755 119.190 41.845 ;
        RECT 122.220 41.595 122.640 41.695 ;
        RECT 118.710 41.365 122.710 41.595 ;
        RECT 122.220 41.275 122.640 41.365 ;
        RECT 118.770 41.115 119.190 41.205 ;
        RECT 118.710 40.885 122.710 41.115 ;
        RECT 118.770 40.785 119.190 40.885 ;
        RECT 122.220 40.635 122.640 40.735 ;
        RECT 118.710 40.405 122.710 40.635 ;
        RECT 122.220 40.315 122.640 40.405 ;
        RECT 118.770 40.155 119.190 40.255 ;
        RECT 118.710 39.925 122.710 40.155 ;
        RECT 118.770 39.835 119.190 39.925 ;
        RECT 122.220 39.675 122.640 39.775 ;
        RECT 118.710 39.445 122.710 39.675 ;
        RECT 122.220 39.355 122.640 39.445 ;
        RECT 118.770 39.195 119.190 39.305 ;
        RECT 113.720 38.885 114.050 39.005 ;
        RECT 118.710 38.965 122.710 39.195 ;
        RECT 122.860 39.085 123.140 44.905 ;
        RECT 123.380 39.085 123.660 44.905 ;
        RECT 123.860 43.995 124.280 44.085 ;
        RECT 123.800 43.765 127.800 43.995 ;
        RECT 123.860 43.665 124.280 43.765 ;
        RECT 127.310 43.515 127.730 43.615 ;
        RECT 123.800 43.285 127.800 43.515 ;
        RECT 127.310 43.195 127.730 43.285 ;
        RECT 123.860 43.035 124.280 43.135 ;
        RECT 123.800 42.805 127.800 43.035 ;
        RECT 123.860 42.715 124.280 42.805 ;
        RECT 127.310 42.555 127.730 42.655 ;
        RECT 123.800 42.325 127.800 42.555 ;
        RECT 127.310 42.235 127.730 42.325 ;
        RECT 123.860 42.075 124.280 42.165 ;
        RECT 123.800 41.845 127.800 42.075 ;
        RECT 123.860 41.745 124.280 41.845 ;
        RECT 127.310 41.595 127.730 41.695 ;
        RECT 123.800 41.365 127.800 41.595 ;
        RECT 127.310 41.275 127.730 41.365 ;
        RECT 123.860 41.115 124.280 41.215 ;
        RECT 123.800 40.885 127.800 41.115 ;
        RECT 123.860 40.795 124.280 40.885 ;
        RECT 127.310 40.635 127.730 40.735 ;
        RECT 123.800 40.405 127.800 40.635 ;
        RECT 127.310 40.315 127.730 40.405 ;
        RECT 123.860 40.155 124.280 40.255 ;
        RECT 123.800 39.925 127.800 40.155 ;
        RECT 123.860 39.835 124.280 39.925 ;
        RECT 127.310 39.675 127.730 39.775 ;
        RECT 123.800 39.445 127.800 39.675 ;
        RECT 127.940 39.525 128.220 44.905 ;
        RECT 129.190 45.085 137.050 45.815 ;
        RECT 129.190 44.895 131.420 45.085 ;
        RECT 127.310 39.355 127.730 39.445 ;
        RECT 123.860 39.195 124.280 39.295 ;
        RECT 123.800 38.965 127.800 39.195 ;
        RECT 118.770 38.885 119.190 38.965 ;
        RECT 123.860 38.875 124.280 38.965 ;
        RECT 111.075 37.625 113.320 38.145 ;
        RECT 102.680 36.170 108.105 36.935 ;
        RECT 102.680 34.415 104.910 36.170 ;
        RECT 111.075 34.610 111.665 37.625 ;
        RECT 114.300 37.445 114.620 38.095 ;
        RECT 114.260 37.425 115.370 37.445 ;
        RECT 116.595 37.425 117.270 37.570 ;
        RECT 114.260 37.045 117.270 37.425 ;
        RECT 115.090 37.040 117.270 37.045 ;
        RECT 116.595 35.335 117.270 37.040 ;
        RECT 118.645 35.335 119.330 38.075 ;
        RECT 123.250 35.335 124.250 35.415 ;
        RECT 116.595 34.660 124.250 35.335 ;
        RECT 129.190 35.230 130.190 44.895 ;
        RECT 131.150 39.045 131.410 44.895 ;
        RECT 131.650 43.935 132.060 44.005 ;
        RECT 131.595 43.705 136.595 43.935 ;
        RECT 131.650 43.635 132.060 43.705 ;
        RECT 136.090 43.455 136.500 43.525 ;
        RECT 131.595 43.225 136.595 43.455 ;
        RECT 136.090 43.145 136.500 43.225 ;
        RECT 131.650 42.975 132.060 43.045 ;
        RECT 131.595 42.745 136.595 42.975 ;
        RECT 131.650 42.675 132.060 42.745 ;
        RECT 136.090 42.495 136.500 42.575 ;
        RECT 131.595 42.265 136.595 42.495 ;
        RECT 136.090 42.195 136.500 42.265 ;
        RECT 131.650 42.015 132.060 42.085 ;
        RECT 131.595 41.785 136.595 42.015 ;
        RECT 131.650 41.715 132.060 41.785 ;
        RECT 136.090 41.535 136.500 41.615 ;
        RECT 131.595 41.305 136.595 41.535 ;
        RECT 136.090 41.235 136.500 41.305 ;
        RECT 131.650 41.055 132.060 41.125 ;
        RECT 131.595 40.825 136.595 41.055 ;
        RECT 131.650 40.755 132.060 40.825 ;
        RECT 136.090 40.575 136.500 40.655 ;
        RECT 131.595 40.345 136.595 40.575 ;
        RECT 136.090 40.275 136.500 40.345 ;
        RECT 131.650 40.095 132.060 40.165 ;
        RECT 131.595 39.865 136.595 40.095 ;
        RECT 131.650 39.795 132.060 39.865 ;
        RECT 136.090 39.615 136.500 39.695 ;
        RECT 131.595 39.385 136.595 39.615 ;
        RECT 136.090 39.315 136.500 39.385 ;
        RECT 131.650 39.135 132.060 39.205 ;
        RECT 131.595 38.905 136.595 39.135 ;
        RECT 136.790 39.045 137.050 45.085 ;
        RECT 140.550 45.745 140.785 45.835 ;
        RECT 140.995 45.795 145.995 46.025 ;
        RECT 141.060 45.775 145.940 45.795 ;
        RECT 140.550 44.785 140.790 45.745 ;
        RECT 137.300 42.985 138.020 42.995 ;
        RECT 137.260 41.765 138.020 42.985 ;
        RECT 137.260 41.005 139.030 41.765 ;
        RECT 137.260 39.965 138.020 41.005 ;
        RECT 137.260 39.955 137.980 39.965 ;
        RECT 131.650 38.835 132.060 38.905 ;
        RECT 138.270 35.595 139.030 41.005 ;
        RECT 140.550 39.195 140.785 44.785 ;
        RECT 141.040 44.735 145.930 44.805 ;
        RECT 140.995 44.505 145.995 44.735 ;
        RECT 141.040 44.465 145.930 44.505 ;
        RECT 143.430 43.105 144.550 44.465 ;
        RECT 143.430 41.985 145.310 43.105 ;
        RECT 143.430 40.625 144.550 41.985 ;
        RECT 141.020 40.615 145.910 40.625 ;
        RECT 141.020 40.565 145.930 40.615 ;
        RECT 140.985 40.335 145.985 40.565 ;
        RECT 141.020 40.305 145.930 40.335 ;
        RECT 141.020 40.285 145.910 40.305 ;
        RECT 146.200 40.285 146.430 47.860 ;
        RECT 149.010 45.835 151.240 53.395 ;
        RECT 146.620 44.645 151.240 45.835 ;
        RECT 146.980 43.105 148.100 43.135 ;
        RECT 149.010 43.105 151.240 44.645 ;
        RECT 146.980 41.985 151.240 43.105 ;
        RECT 146.980 41.955 148.100 41.985 ;
        RECT 149.010 40.375 151.240 41.985 ;
        RECT 146.190 39.325 146.430 40.285 ;
        RECT 141.040 39.275 146.010 39.305 ;
        RECT 140.555 36.890 140.785 39.195 ;
        RECT 140.985 39.045 146.010 39.275 ;
        RECT 141.040 38.985 146.010 39.045 ;
        RECT 146.195 39.195 146.430 39.325 ;
        RECT 143.700 37.395 144.260 38.985 ;
        RECT 146.195 36.890 146.425 39.195 ;
        RECT 146.600 39.185 151.240 40.375 ;
        RECT 140.555 36.660 146.425 36.890 ;
        RECT 114.710 34.610 115.395 34.640 ;
        RECT 111.075 34.415 115.395 34.610 ;
        RECT 123.250 34.415 124.250 34.660 ;
        RECT 102.680 34.105 115.395 34.415 ;
        RECT 102.690 33.925 115.395 34.105 ;
        RECT 102.690 33.830 111.665 33.925 ;
        RECT 114.710 33.895 115.395 33.925 ;
        RECT 123.360 32.540 124.165 34.415 ;
        RECT 129.120 34.395 130.190 35.230 ;
        RECT 123.330 31.735 124.195 32.540 ;
        RECT 129.120 31.235 130.040 34.395 ;
        RECT 149.010 34.005 151.240 39.185 ;
      LAYER via ;
        RECT 103.150 160.830 104.650 162.330 ;
        RECT 149.350 161.110 150.850 162.610 ;
        RECT 118.165 147.805 119.055 148.695 ;
        RECT 138.730 147.745 139.585 148.600 ;
        RECT 104.290 140.835 104.740 142.035 ;
        RECT 108.580 140.735 108.860 141.085 ;
        RECT 111.250 142.670 111.885 143.305 ;
        RECT 118.235 143.810 119.085 144.660 ;
        RECT 131.955 143.275 132.985 144.305 ;
        RECT 108.590 136.145 108.870 136.495 ;
        RECT 108.590 131.575 108.870 131.925 ;
        RECT 108.590 126.985 108.870 127.335 ;
        RECT 108.590 122.415 108.870 122.765 ;
        RECT 108.590 117.815 108.870 118.165 ;
        RECT 114.570 140.755 114.880 141.035 ;
        RECT 113.860 138.425 114.140 138.775 ;
        RECT 116.535 138.625 117.280 139.370 ;
        RECT 114.570 136.175 114.880 136.455 ;
        RECT 113.860 133.845 114.140 134.195 ;
        RECT 114.570 131.595 114.880 131.875 ;
        RECT 113.870 129.275 114.150 129.625 ;
        RECT 146.920 143.275 147.950 144.305 ;
        RECT 114.570 127.015 114.880 127.295 ;
        RECT 113.860 124.685 114.140 125.035 ;
        RECT 114.550 122.445 114.860 122.725 ;
        RECT 113.860 120.105 114.140 120.455 ;
        RECT 111.215 116.040 111.525 116.350 ;
        RECT 114.560 117.865 114.870 118.145 ;
        RECT 120.505 126.790 121.355 127.640 ;
        RECT 108.580 113.365 108.840 113.695 ;
        RECT 109.260 111.085 109.520 111.415 ;
        RECT 108.580 108.785 108.840 109.115 ;
        RECT 109.260 106.495 109.520 106.825 ;
        RECT 108.580 104.205 108.840 104.535 ;
        RECT 109.260 101.925 109.520 102.255 ;
        RECT 108.580 99.625 108.840 99.955 ;
        RECT 109.260 97.345 109.520 97.675 ;
        RECT 108.580 95.045 108.840 95.375 ;
        RECT 109.260 92.755 109.520 93.085 ;
        RECT 108.580 90.465 108.840 90.795 ;
        RECT 127.040 126.575 127.340 126.895 ;
        RECT 126.390 125.965 126.690 126.315 ;
        RECT 127.040 125.395 127.340 125.715 ;
        RECT 126.390 124.785 126.690 125.135 ;
        RECT 127.040 124.215 127.340 124.535 ;
        RECT 126.390 123.605 126.690 123.955 ;
        RECT 127.040 123.035 127.340 123.355 ;
        RECT 126.390 122.425 126.690 122.775 ;
        RECT 127.040 121.855 127.340 122.175 ;
        RECT 126.390 121.245 126.690 121.595 ;
        RECT 127.040 120.675 127.340 120.995 ;
        RECT 129.140 126.575 129.440 126.895 ;
        RECT 128.470 125.965 128.770 126.315 ;
        RECT 129.140 125.395 129.440 125.715 ;
        RECT 128.470 124.785 128.770 125.135 ;
        RECT 129.140 124.215 129.440 124.535 ;
        RECT 128.470 123.605 128.770 123.955 ;
        RECT 129.140 123.035 129.440 123.355 ;
        RECT 128.470 122.425 128.770 122.775 ;
        RECT 129.140 121.855 129.440 122.175 ;
        RECT 128.470 121.245 128.770 121.595 ;
        RECT 129.140 120.675 129.440 120.995 ;
        RECT 131.210 126.575 131.510 126.895 ;
        RECT 130.550 125.975 130.850 126.325 ;
        RECT 131.220 125.395 131.520 125.715 ;
        RECT 130.550 124.785 130.850 125.135 ;
        RECT 131.220 124.205 131.520 124.525 ;
        RECT 130.550 123.605 130.850 123.955 ;
        RECT 131.220 123.035 131.520 123.355 ;
        RECT 130.550 122.425 130.850 122.775 ;
        RECT 131.220 121.855 131.520 122.175 ;
        RECT 130.550 121.235 130.850 121.585 ;
        RECT 131.220 120.675 131.520 120.995 ;
        RECT 133.310 126.575 133.610 126.895 ;
        RECT 132.650 125.975 132.950 126.325 ;
        RECT 133.310 125.395 133.610 125.715 ;
        RECT 132.650 124.785 132.950 125.135 ;
        RECT 133.310 124.215 133.610 124.535 ;
        RECT 132.650 123.605 132.950 123.955 ;
        RECT 133.310 123.035 133.610 123.355 ;
        RECT 132.650 122.425 132.950 122.775 ;
        RECT 133.310 121.855 133.610 122.175 ;
        RECT 132.650 121.245 132.950 121.595 ;
        RECT 133.310 120.665 133.610 120.985 ;
        RECT 135.400 126.565 135.700 126.885 ;
        RECT 134.720 125.965 135.020 126.315 ;
        RECT 135.400 125.395 135.700 125.715 ;
        RECT 134.730 124.785 135.030 125.135 ;
        RECT 135.400 124.215 135.700 124.535 ;
        RECT 134.730 123.605 135.030 123.955 ;
        RECT 135.400 123.035 135.700 123.355 ;
        RECT 134.730 122.435 135.030 122.785 ;
        RECT 135.400 121.855 135.700 122.175 ;
        RECT 134.730 121.245 135.030 121.595 ;
        RECT 135.400 120.675 135.700 120.995 ;
        RECT 145.860 127.835 146.140 128.145 ;
        RECT 145.230 126.545 145.530 126.865 ;
        RECT 145.870 125.265 146.150 125.575 ;
        RECT 145.230 123.965 145.530 124.285 ;
        RECT 145.880 122.675 146.160 122.985 ;
        RECT 145.230 121.385 145.530 121.705 ;
        RECT 145.200 120.390 145.470 120.660 ;
        RECT 123.250 115.550 124.675 116.975 ;
        RECT 116.580 111.240 117.445 112.105 ;
        RECT 127.050 119.035 127.340 119.355 ;
        RECT 126.400 118.455 126.700 118.755 ;
        RECT 127.050 117.855 127.340 118.175 ;
        RECT 126.400 117.275 126.700 117.575 ;
        RECT 127.050 116.675 127.340 116.995 ;
        RECT 126.400 116.095 126.700 116.395 ;
        RECT 127.050 115.495 127.340 115.815 ;
        RECT 126.400 114.905 126.700 115.205 ;
        RECT 127.050 114.325 127.340 114.645 ;
        RECT 126.400 113.735 126.700 114.035 ;
        RECT 127.050 113.135 127.340 113.455 ;
        RECT 129.150 119.035 129.440 119.355 ;
        RECT 128.490 118.455 128.790 118.755 ;
        RECT 129.150 117.855 129.440 118.175 ;
        RECT 128.490 117.275 128.790 117.575 ;
        RECT 129.150 116.675 129.440 116.995 ;
        RECT 128.490 116.095 128.790 116.395 ;
        RECT 129.150 115.495 129.440 115.815 ;
        RECT 128.490 114.915 128.790 115.215 ;
        RECT 129.150 114.315 129.440 114.635 ;
        RECT 128.490 113.735 128.790 114.035 ;
        RECT 129.150 113.135 129.440 113.455 ;
        RECT 131.230 119.035 131.520 119.355 ;
        RECT 130.570 118.455 130.870 118.755 ;
        RECT 131.230 117.855 131.520 118.175 ;
        RECT 130.570 117.275 130.870 117.575 ;
        RECT 131.230 116.665 131.520 116.985 ;
        RECT 130.570 116.095 130.870 116.395 ;
        RECT 131.230 115.495 131.520 115.815 ;
        RECT 130.570 114.915 130.870 115.215 ;
        RECT 131.230 114.315 131.520 114.635 ;
        RECT 130.570 113.735 130.870 114.035 ;
        RECT 131.240 113.135 131.530 113.455 ;
        RECT 133.310 119.035 133.600 119.355 ;
        RECT 132.630 118.455 132.930 118.755 ;
        RECT 133.310 117.855 133.600 118.175 ;
        RECT 132.630 117.275 132.930 117.575 ;
        RECT 133.310 116.675 133.600 116.995 ;
        RECT 132.630 116.095 132.930 116.395 ;
        RECT 133.310 115.495 133.600 115.815 ;
        RECT 132.630 114.915 132.930 115.215 ;
        RECT 133.310 114.315 133.600 114.635 ;
        RECT 132.630 113.735 132.930 114.035 ;
        RECT 133.310 113.135 133.600 113.455 ;
        RECT 135.400 119.035 135.690 119.355 ;
        RECT 134.730 118.455 135.030 118.755 ;
        RECT 135.400 117.855 135.690 118.175 ;
        RECT 134.730 117.275 135.030 117.575 ;
        RECT 135.400 116.675 135.690 116.995 ;
        RECT 134.730 116.095 135.030 116.395 ;
        RECT 135.400 115.495 135.690 115.815 ;
        RECT 134.730 114.915 135.030 115.215 ;
        RECT 135.400 114.315 135.690 114.635 ;
        RECT 134.730 113.735 135.030 114.035 ;
        RECT 135.400 113.135 135.690 113.455 ;
        RECT 145.190 118.045 145.490 118.365 ;
        RECT 145.880 116.775 146.160 117.085 ;
        RECT 145.190 115.475 145.490 115.795 ;
        RECT 145.880 114.185 146.160 114.495 ;
        RECT 145.190 112.885 145.490 113.205 ;
        RECT 145.880 111.605 146.160 111.915 ;
        RECT 118.430 109.155 119.230 109.955 ;
        RECT 107.180 89.340 107.525 89.685 ;
        RECT 112.115 98.050 112.990 98.925 ;
        RECT 114.280 107.085 114.700 107.425 ;
        RECT 115.800 106.505 116.220 106.805 ;
        RECT 114.280 105.905 114.700 106.245 ;
        RECT 115.800 105.325 116.220 105.625 ;
        RECT 114.280 104.715 114.700 105.055 ;
        RECT 115.800 104.155 116.220 104.455 ;
        RECT 114.280 103.535 114.700 103.875 ;
        RECT 115.800 102.975 116.220 103.275 ;
        RECT 114.280 102.355 114.700 102.695 ;
        RECT 115.800 101.795 116.220 102.095 ;
        RECT 114.280 101.175 114.700 101.515 ;
        RECT 115.800 100.615 116.220 100.915 ;
        RECT 114.280 99.995 114.700 100.335 ;
        RECT 115.800 99.435 116.220 99.735 ;
        RECT 114.290 98.815 114.710 99.155 ;
        RECT 115.800 98.255 116.220 98.555 ;
        RECT 114.290 97.635 114.710 97.975 ;
        RECT 115.800 97.075 116.220 97.375 ;
        RECT 114.290 96.455 114.710 96.795 ;
        RECT 115.800 95.895 116.220 96.195 ;
        RECT 114.290 95.275 114.710 95.615 ;
        RECT 108.550 87.045 108.930 87.415 ;
        RECT 109.200 84.715 109.570 85.105 ;
        RECT 108.550 82.445 108.930 82.815 ;
        RECT 109.200 80.145 109.570 80.535 ;
        RECT 108.550 77.865 108.930 78.235 ;
        RECT 109.200 75.565 109.570 75.955 ;
        RECT 108.550 73.285 108.930 73.655 ;
        RECT 109.200 70.995 109.570 71.385 ;
        RECT 108.550 68.705 108.930 69.075 ;
        RECT 109.200 66.395 109.570 66.785 ;
        RECT 108.550 64.125 108.930 64.495 ;
        RECT 107.005 63.125 107.375 63.495 ;
        RECT 123.760 107.475 124.190 107.815 ;
        RECT 121.700 106.165 122.210 106.535 ;
        RECT 123.760 104.895 124.190 105.235 ;
        RECT 121.700 103.585 122.210 103.955 ;
        RECT 123.760 102.305 124.190 102.645 ;
        RECT 121.700 100.995 122.210 101.365 ;
        RECT 123.760 99.735 124.190 100.075 ;
        RECT 121.660 98.435 122.170 98.805 ;
        RECT 123.770 97.155 124.200 97.495 ;
        RECT 121.700 95.845 122.210 96.215 ;
        RECT 123.770 94.565 124.200 94.905 ;
        RECT 121.700 93.265 122.210 93.635 ;
        RECT 123.770 91.995 124.200 92.335 ;
        RECT 121.690 90.685 122.200 91.055 ;
        RECT 123.770 89.405 124.200 89.745 ;
        RECT 121.680 88.105 122.190 88.475 ;
        RECT 123.770 86.835 124.200 87.175 ;
        RECT 121.690 85.525 122.200 85.895 ;
        RECT 123.770 84.255 124.200 84.595 ;
        RECT 121.690 82.945 122.200 83.315 ;
        RECT 123.770 81.665 124.200 82.005 ;
        RECT 127.400 107.475 127.830 107.815 ;
        RECT 125.350 106.165 125.860 106.535 ;
        RECT 127.400 104.895 127.830 105.235 ;
        RECT 125.370 103.585 125.880 103.955 ;
        RECT 127.400 102.315 127.830 102.655 ;
        RECT 125.350 101.005 125.860 101.375 ;
        RECT 127.400 99.735 127.830 100.075 ;
        RECT 125.370 98.425 125.880 98.795 ;
        RECT 127.400 97.155 127.830 97.495 ;
        RECT 125.390 95.835 125.900 96.205 ;
        RECT 127.400 94.575 127.830 94.915 ;
        RECT 125.370 93.265 125.880 93.635 ;
        RECT 127.400 92.005 127.830 92.345 ;
        RECT 125.380 90.685 125.890 91.055 ;
        RECT 127.400 89.415 127.830 89.755 ;
        RECT 125.370 88.105 125.880 88.475 ;
        RECT 127.400 86.835 127.830 87.175 ;
        RECT 125.370 85.515 125.880 85.885 ;
        RECT 127.400 84.255 127.830 84.595 ;
        RECT 125.370 82.955 125.880 83.325 ;
        RECT 127.400 81.665 127.830 82.005 ;
        RECT 131.150 107.475 131.580 107.815 ;
        RECT 129.060 106.165 129.570 106.535 ;
        RECT 131.150 104.895 131.580 105.235 ;
        RECT 129.060 103.585 129.570 103.955 ;
        RECT 131.150 102.325 131.580 102.665 ;
        RECT 129.030 101.005 129.540 101.375 ;
        RECT 131.150 99.735 131.580 100.075 ;
        RECT 129.060 98.425 129.570 98.795 ;
        RECT 131.150 97.155 131.580 97.495 ;
        RECT 129.050 95.845 129.560 96.215 ;
        RECT 131.150 94.575 131.580 94.915 ;
        RECT 129.050 93.265 129.560 93.635 ;
        RECT 131.150 91.995 131.580 92.335 ;
        RECT 129.050 90.685 129.560 91.055 ;
        RECT 131.150 89.415 131.580 89.755 ;
        RECT 129.050 88.105 129.560 88.475 ;
        RECT 131.150 86.835 131.580 87.175 ;
        RECT 129.040 85.525 129.550 85.895 ;
        RECT 131.150 84.255 131.580 84.595 ;
        RECT 129.050 82.945 129.560 83.315 ;
        RECT 131.150 81.665 131.580 82.005 ;
        RECT 134.790 107.475 135.220 107.815 ;
        RECT 132.730 106.165 133.240 106.535 ;
        RECT 134.790 104.895 135.220 105.235 ;
        RECT 132.730 103.605 133.240 103.975 ;
        RECT 134.790 102.315 135.220 102.655 ;
        RECT 132.720 101.015 133.230 101.385 ;
        RECT 134.790 99.735 135.220 100.075 ;
        RECT 132.740 98.435 133.250 98.805 ;
        RECT 134.790 97.155 135.220 97.495 ;
        RECT 132.730 95.845 133.240 96.215 ;
        RECT 134.790 94.575 135.220 94.915 ;
        RECT 132.730 93.275 133.240 93.645 ;
        RECT 134.790 91.995 135.220 92.335 ;
        RECT 132.740 90.695 133.250 91.065 ;
        RECT 134.790 89.415 135.220 89.755 ;
        RECT 132.720 88.105 133.230 88.475 ;
        RECT 134.790 86.825 135.220 87.165 ;
        RECT 132.730 85.525 133.240 85.895 ;
        RECT 134.790 84.245 135.220 84.585 ;
        RECT 132.740 82.945 133.250 83.315 ;
        RECT 134.790 81.665 135.220 82.005 ;
        RECT 138.500 107.475 138.930 107.815 ;
        RECT 136.440 106.175 136.950 106.545 ;
        RECT 138.500 104.895 138.930 105.235 ;
        RECT 136.440 103.595 136.950 103.965 ;
        RECT 138.500 102.315 138.930 102.655 ;
        RECT 136.440 100.995 136.950 101.365 ;
        RECT 138.500 99.735 138.930 100.075 ;
        RECT 136.440 98.435 136.950 98.805 ;
        RECT 138.500 97.155 138.930 97.495 ;
        RECT 136.440 95.845 136.950 96.215 ;
        RECT 138.500 94.575 138.930 94.915 ;
        RECT 136.440 93.285 136.950 93.655 ;
        RECT 138.500 91.995 138.930 92.335 ;
        RECT 136.440 90.685 136.950 91.055 ;
        RECT 138.500 89.415 138.930 89.755 ;
        RECT 136.440 88.095 136.950 88.465 ;
        RECT 138.500 86.835 138.930 87.175 ;
        RECT 136.440 85.525 136.950 85.895 ;
        RECT 138.500 84.255 138.930 84.595 ;
        RECT 136.440 82.945 136.950 83.315 ;
        RECT 138.500 81.675 138.930 82.015 ;
        RECT 142.140 107.475 142.570 107.815 ;
        RECT 140.110 106.175 140.620 106.545 ;
        RECT 142.140 104.895 142.570 105.235 ;
        RECT 140.110 103.595 140.620 103.965 ;
        RECT 142.140 102.305 142.570 102.645 ;
        RECT 140.110 100.995 140.620 101.365 ;
        RECT 142.140 99.735 142.570 100.075 ;
        RECT 140.110 98.435 140.620 98.805 ;
        RECT 142.140 97.155 142.570 97.495 ;
        RECT 140.110 95.845 140.620 96.215 ;
        RECT 142.140 94.575 142.570 94.915 ;
        RECT 140.110 93.275 140.620 93.645 ;
        RECT 142.140 91.995 142.570 92.335 ;
        RECT 140.110 90.685 140.620 91.055 ;
        RECT 142.150 89.415 142.580 89.755 ;
        RECT 140.110 88.095 140.620 88.465 ;
        RECT 142.150 86.835 142.580 87.175 ;
        RECT 140.110 85.515 140.620 85.885 ;
        RECT 142.150 84.255 142.580 84.595 ;
        RECT 140.110 82.935 140.620 83.305 ;
        RECT 142.150 81.665 142.580 82.005 ;
        RECT 145.830 107.475 146.260 107.815 ;
        RECT 143.790 106.165 144.300 106.535 ;
        RECT 145.830 104.885 146.260 105.225 ;
        RECT 143.790 103.585 144.300 103.955 ;
        RECT 145.830 102.305 146.260 102.645 ;
        RECT 143.790 101.005 144.300 101.375 ;
        RECT 145.830 99.725 146.260 100.065 ;
        RECT 143.790 98.425 144.300 98.795 ;
        RECT 145.830 97.145 146.260 97.485 ;
        RECT 143.790 95.845 144.300 96.215 ;
        RECT 145.830 94.565 146.260 94.905 ;
        RECT 143.790 93.265 144.300 93.635 ;
        RECT 145.830 91.985 146.260 92.325 ;
        RECT 143.790 90.695 144.300 91.065 ;
        RECT 145.830 89.405 146.260 89.745 ;
        RECT 143.800 88.105 144.310 88.475 ;
        RECT 145.830 86.835 146.260 87.175 ;
        RECT 143.800 85.525 144.310 85.895 ;
        RECT 145.830 84.245 146.260 84.585 ;
        RECT 143.820 82.935 144.330 83.305 ;
        RECT 145.830 81.665 146.260 82.005 ;
        RECT 108.570 61.225 108.910 61.585 ;
        RECT 109.200 58.935 109.520 59.295 ;
        RECT 108.570 56.635 108.910 56.995 ;
        RECT 109.200 54.365 109.520 54.725 ;
        RECT 108.570 52.075 108.910 52.435 ;
        RECT 109.200 49.775 109.520 50.135 ;
        RECT 108.570 47.495 108.910 47.855 ;
        RECT 109.200 45.195 109.520 45.555 ;
        RECT 108.570 42.905 108.910 43.265 ;
        RECT 109.200 40.615 109.520 40.975 ;
        RECT 108.570 38.325 108.910 38.685 ;
        RECT 110.855 52.300 111.905 53.350 ;
        RECT 116.730 52.300 117.780 53.350 ;
        RECT 113.720 43.525 114.050 43.885 ;
        RECT 114.280 41.245 114.610 41.595 ;
        RECT 113.720 38.935 114.050 39.295 ;
        RECT 123.770 77.115 124.200 77.455 ;
        RECT 121.680 75.805 122.200 76.205 ;
        RECT 123.770 74.525 124.200 74.865 ;
        RECT 121.680 73.215 122.200 73.615 ;
        RECT 123.770 71.955 124.200 72.295 ;
        RECT 121.670 70.625 122.190 71.025 ;
        RECT 123.770 69.375 124.200 69.715 ;
        RECT 121.690 68.055 122.210 68.455 ;
        RECT 123.770 66.795 124.200 67.135 ;
        RECT 121.700 65.475 122.220 65.875 ;
        RECT 123.770 64.215 124.200 64.555 ;
        RECT 121.680 62.895 122.200 63.295 ;
        RECT 123.770 61.635 124.200 61.975 ;
        RECT 121.690 60.295 122.210 60.695 ;
        RECT 123.770 59.055 124.200 59.395 ;
        RECT 121.690 57.735 122.210 58.135 ;
        RECT 123.770 56.475 124.200 56.815 ;
        RECT 121.700 55.145 122.220 55.545 ;
        RECT 123.770 53.895 124.200 54.235 ;
        RECT 121.700 52.565 122.220 52.965 ;
        RECT 123.770 51.315 124.200 51.655 ;
        RECT 127.400 77.115 127.830 77.455 ;
        RECT 125.370 75.795 125.890 76.195 ;
        RECT 127.410 74.535 127.840 74.875 ;
        RECT 125.350 73.205 125.870 73.605 ;
        RECT 127.410 71.955 127.840 72.295 ;
        RECT 125.370 70.635 125.890 71.035 ;
        RECT 127.410 69.375 127.840 69.715 ;
        RECT 125.370 68.055 125.890 68.455 ;
        RECT 127.410 66.795 127.840 67.135 ;
        RECT 125.350 65.465 125.870 65.865 ;
        RECT 127.410 64.215 127.840 64.555 ;
        RECT 125.370 62.885 125.890 63.285 ;
        RECT 127.410 61.635 127.840 61.975 ;
        RECT 125.390 60.305 125.910 60.705 ;
        RECT 127.410 59.055 127.840 59.395 ;
        RECT 125.370 57.735 125.890 58.135 ;
        RECT 127.410 56.475 127.840 56.815 ;
        RECT 125.380 55.155 125.900 55.555 ;
        RECT 127.410 53.895 127.840 54.235 ;
        RECT 125.370 52.575 125.890 52.975 ;
        RECT 127.410 51.315 127.840 51.655 ;
        RECT 131.150 77.115 131.580 77.455 ;
        RECT 129.060 75.795 129.580 76.195 ;
        RECT 131.150 74.545 131.580 74.885 ;
        RECT 129.040 73.205 129.560 73.605 ;
        RECT 131.150 71.955 131.580 72.295 ;
        RECT 129.060 70.625 129.580 71.025 ;
        RECT 131.150 69.375 131.580 69.715 ;
        RECT 129.050 68.045 129.570 68.445 ;
        RECT 131.150 66.795 131.580 67.135 ;
        RECT 129.050 65.485 129.570 65.885 ;
        RECT 131.150 64.205 131.580 64.545 ;
        RECT 129.050 62.885 129.570 63.285 ;
        RECT 131.150 61.645 131.580 61.985 ;
        RECT 129.060 60.305 129.580 60.705 ;
        RECT 131.150 59.055 131.580 59.395 ;
        RECT 129.040 57.745 129.560 58.145 ;
        RECT 131.150 56.485 131.580 56.825 ;
        RECT 129.050 55.145 129.570 55.545 ;
        RECT 131.150 53.895 131.580 54.235 ;
        RECT 129.050 52.585 129.570 52.985 ;
        RECT 131.150 51.315 131.580 51.655 ;
        RECT 134.790 77.115 135.220 77.455 ;
        RECT 132.740 75.795 133.260 76.195 ;
        RECT 134.790 74.535 135.220 74.875 ;
        RECT 132.740 73.205 133.260 73.605 ;
        RECT 134.790 71.955 135.220 72.295 ;
        RECT 132.740 70.635 133.260 71.035 ;
        RECT 134.790 69.375 135.220 69.715 ;
        RECT 132.740 68.045 133.260 68.445 ;
        RECT 134.790 66.795 135.220 67.135 ;
        RECT 132.740 65.485 133.260 65.885 ;
        RECT 134.790 64.215 135.220 64.555 ;
        RECT 132.730 62.885 133.250 63.285 ;
        RECT 134.790 61.635 135.220 61.975 ;
        RECT 132.740 60.305 133.260 60.705 ;
        RECT 134.790 59.055 135.220 59.395 ;
        RECT 132.740 57.715 133.260 58.115 ;
        RECT 134.790 56.475 135.220 56.815 ;
        RECT 132.740 55.145 133.260 55.545 ;
        RECT 134.790 53.895 135.220 54.235 ;
        RECT 132.740 52.575 133.260 52.975 ;
        RECT 134.790 51.305 135.220 51.645 ;
        RECT 138.490 77.105 138.920 77.445 ;
        RECT 136.410 75.795 136.930 76.195 ;
        RECT 138.490 74.545 138.920 74.885 ;
        RECT 136.400 73.215 136.920 73.615 ;
        RECT 138.490 71.955 138.920 72.295 ;
        RECT 136.410 70.625 136.930 71.025 ;
        RECT 138.490 69.375 138.920 69.715 ;
        RECT 136.400 68.045 136.920 68.445 ;
        RECT 138.490 66.795 138.920 67.135 ;
        RECT 136.400 65.465 136.920 65.865 ;
        RECT 138.490 64.215 138.920 64.555 ;
        RECT 136.410 62.875 136.930 63.275 ;
        RECT 138.490 61.635 138.920 61.975 ;
        RECT 136.420 60.305 136.940 60.705 ;
        RECT 138.490 59.055 138.920 59.395 ;
        RECT 136.420 57.735 136.940 58.135 ;
        RECT 138.490 56.475 138.920 56.815 ;
        RECT 136.410 55.155 136.930 55.555 ;
        RECT 138.490 53.895 138.920 54.235 ;
        RECT 136.420 52.565 136.940 52.965 ;
        RECT 138.490 51.315 138.920 51.655 ;
        RECT 142.150 77.105 142.580 77.445 ;
        RECT 140.100 75.795 140.620 76.195 ;
        RECT 142.150 74.535 142.580 74.875 ;
        RECT 140.080 73.205 140.600 73.605 ;
        RECT 142.150 71.955 142.580 72.295 ;
        RECT 140.090 70.625 140.610 71.025 ;
        RECT 142.150 69.365 142.580 69.705 ;
        RECT 140.080 68.045 140.600 68.445 ;
        RECT 142.150 66.805 142.580 67.145 ;
        RECT 140.110 65.455 140.630 65.855 ;
        RECT 142.130 64.215 142.560 64.555 ;
        RECT 140.090 62.885 140.610 63.285 ;
        RECT 142.130 61.635 142.560 61.975 ;
        RECT 140.080 60.305 140.600 60.705 ;
        RECT 142.130 59.065 142.560 59.405 ;
        RECT 140.100 57.725 140.620 58.125 ;
        RECT 142.130 56.475 142.560 56.815 ;
        RECT 140.100 55.155 140.620 55.555 ;
        RECT 142.130 53.885 142.560 54.225 ;
        RECT 140.100 52.565 140.620 52.965 ;
        RECT 142.130 51.305 142.560 51.645 ;
        RECT 145.830 77.105 146.260 77.445 ;
        RECT 143.780 75.805 144.300 76.205 ;
        RECT 145.830 74.535 146.260 74.875 ;
        RECT 143.780 73.205 144.300 73.605 ;
        RECT 145.830 71.955 146.260 72.295 ;
        RECT 143.780 70.615 144.300 71.015 ;
        RECT 145.830 69.375 146.260 69.715 ;
        RECT 143.760 68.035 144.280 68.435 ;
        RECT 145.830 66.785 146.260 67.125 ;
        RECT 143.780 65.465 144.300 65.865 ;
        RECT 145.830 64.215 146.260 64.555 ;
        RECT 143.790 62.885 144.310 63.285 ;
        RECT 145.830 61.625 146.260 61.965 ;
        RECT 143.790 60.315 144.310 60.715 ;
        RECT 145.830 59.055 146.260 59.395 ;
        RECT 143.780 57.715 144.300 58.115 ;
        RECT 145.830 56.465 146.260 56.805 ;
        RECT 143.770 55.135 144.290 55.535 ;
        RECT 145.830 53.895 146.260 54.235 ;
        RECT 143.780 52.565 144.300 52.965 ;
        RECT 145.830 51.305 146.260 51.645 ;
        RECT 131.150 47.950 131.880 48.680 ;
        RECT 127.940 45.405 128.220 45.685 ;
        RECT 118.770 43.725 119.190 44.045 ;
        RECT 122.220 43.235 122.640 43.555 ;
        RECT 118.770 42.765 119.190 43.085 ;
        RECT 122.220 42.285 122.640 42.605 ;
        RECT 118.770 41.805 119.190 42.125 ;
        RECT 122.220 41.325 122.640 41.645 ;
        RECT 118.770 40.835 119.190 41.155 ;
        RECT 122.220 40.365 122.640 40.685 ;
        RECT 118.770 39.885 119.190 40.205 ;
        RECT 122.220 39.405 122.640 39.725 ;
        RECT 118.770 38.935 119.190 39.255 ;
        RECT 123.860 43.715 124.280 44.035 ;
        RECT 127.310 43.245 127.730 43.565 ;
        RECT 123.860 42.765 124.280 43.085 ;
        RECT 127.310 42.285 127.730 42.605 ;
        RECT 123.860 41.795 124.280 42.115 ;
        RECT 127.310 41.325 127.730 41.645 ;
        RECT 123.860 40.845 124.280 41.165 ;
        RECT 127.310 40.365 127.730 40.685 ;
        RECT 123.860 39.885 124.280 40.205 ;
        RECT 127.310 39.405 127.730 39.725 ;
        RECT 123.860 38.925 124.280 39.245 ;
        RECT 112.900 37.725 113.220 38.045 ;
        RECT 114.300 37.745 114.620 38.065 ;
        RECT 107.545 36.380 107.895 36.730 ;
        RECT 118.770 37.520 119.200 37.950 ;
        RECT 131.650 43.685 132.060 43.955 ;
        RECT 136.090 43.195 136.500 43.475 ;
        RECT 131.650 42.725 132.060 42.995 ;
        RECT 136.090 42.245 136.500 42.525 ;
        RECT 131.650 41.765 132.060 42.035 ;
        RECT 136.090 41.285 136.500 41.565 ;
        RECT 131.650 40.805 132.060 41.075 ;
        RECT 136.090 40.325 136.500 40.605 ;
        RECT 131.650 39.845 132.060 40.115 ;
        RECT 136.090 39.365 136.500 39.645 ;
        RECT 131.650 38.885 132.060 39.155 ;
        RECT 144.160 41.985 145.280 43.105 ;
        RECT 143.700 37.425 144.260 37.985 ;
        RECT 138.270 35.625 139.030 36.385 ;
        RECT 114.710 33.925 115.395 34.610 ;
        RECT 149.345 34.670 150.030 35.355 ;
        RECT 123.360 31.735 124.165 32.540 ;
        RECT 129.210 31.325 129.955 32.070 ;
      LAYER met2 ;
        RECT 149.350 168.635 150.850 168.660 ;
        RECT 149.330 167.185 150.870 168.635 ;
        RECT 103.150 165.045 104.650 165.070 ;
        RECT 103.130 163.595 104.670 165.045 ;
        RECT 103.150 160.800 104.650 163.595 ;
        RECT 149.350 161.080 150.850 167.185 ;
        RECT 118.165 149.910 119.055 149.935 ;
        RECT 118.145 149.070 119.075 149.910 ;
        RECT 138.730 149.855 139.585 149.880 ;
        RECT 118.165 147.775 119.055 149.070 ;
        RECT 138.710 149.050 139.605 149.855 ;
        RECT 138.730 147.715 139.585 149.050 ;
        RECT 111.250 143.305 111.885 143.335 ;
        RECT 116.535 143.305 117.280 143.360 ;
        RECT 111.250 142.670 117.280 143.305 ;
        RECT 111.250 142.640 111.885 142.670 ;
        RECT 104.370 142.175 108.830 142.475 ;
        RECT 104.370 142.035 104.670 142.175 ;
        RECT 104.240 140.835 104.790 142.035 ;
        RECT 108.530 141.085 108.830 142.175 ;
        RECT 108.530 140.735 108.910 141.085 ;
        RECT 108.530 136.495 108.830 140.735 ;
        RECT 113.830 138.775 114.140 141.135 ;
        RECT 114.560 141.035 114.880 141.125 ;
        RECT 114.520 140.755 114.930 141.035 ;
        RECT 113.810 138.425 114.190 138.775 ;
        RECT 108.530 136.145 108.920 136.495 ;
        RECT 108.530 131.925 108.830 136.145 ;
        RECT 113.830 134.195 114.140 138.425 ;
        RECT 114.560 136.455 114.880 140.755 ;
        RECT 116.535 138.595 117.280 142.670 ;
        RECT 114.520 136.175 114.930 136.455 ;
        RECT 113.810 133.845 114.190 134.195 ;
        RECT 108.530 131.575 108.920 131.925 ;
        RECT 108.530 127.335 108.830 131.575 ;
        RECT 113.830 129.625 114.140 133.845 ;
        RECT 114.560 131.875 114.880 136.175 ;
        RECT 114.520 131.595 114.930 131.875 ;
        RECT 113.820 129.275 114.200 129.625 ;
        RECT 108.530 126.985 108.920 127.335 ;
        RECT 108.530 122.765 108.830 126.985 ;
        RECT 113.830 125.035 114.140 129.275 ;
        RECT 114.560 127.295 114.880 131.595 ;
        RECT 118.235 127.640 119.085 144.690 ;
        RECT 146.920 144.305 147.950 144.335 ;
        RECT 131.925 143.275 147.950 144.305 ;
        RECT 146.920 143.245 147.950 143.275 ;
        RECT 126.370 129.545 126.650 129.580 ;
        RECT 120.505 127.640 121.355 127.670 ;
        RECT 114.520 127.015 114.930 127.295 ;
        RECT 113.810 124.685 114.190 125.035 ;
        RECT 108.530 122.415 108.920 122.765 ;
        RECT 108.530 118.165 108.830 122.415 ;
        RECT 113.830 120.455 114.140 124.685 ;
        RECT 114.560 122.725 114.880 127.015 ;
        RECT 118.235 126.855 121.355 127.640 ;
        RECT 118.245 126.790 121.355 126.855 ;
        RECT 120.505 126.760 121.355 126.790 ;
        RECT 126.360 127.555 126.660 129.545 ;
        RECT 141.085 129.510 144.145 129.710 ;
        RECT 141.085 129.200 145.490 129.510 ;
        RECT 141.085 129.000 144.145 129.200 ;
        RECT 127.095 128.890 135.740 128.960 ;
        RECT 141.085 128.890 141.795 129.000 ;
        RECT 127.095 128.670 141.795 128.890 ;
        RECT 127.095 127.795 127.385 128.670 ;
        RECT 127.080 127.570 127.385 127.795 ;
        RECT 126.360 126.315 126.650 127.555 ;
        RECT 127.080 126.895 127.370 127.570 ;
        RECT 128.370 127.445 128.790 127.855 ;
        RECT 126.990 126.575 127.390 126.895 ;
        RECT 126.340 125.965 126.740 126.315 ;
        RECT 126.360 125.135 126.650 125.965 ;
        RECT 127.080 125.715 127.370 126.575 ;
        RECT 128.430 126.315 128.720 127.445 ;
        RECT 129.180 126.895 129.470 128.670 ;
        RECT 130.450 127.445 130.870 127.855 ;
        RECT 129.090 126.575 129.490 126.895 ;
        RECT 128.420 125.965 128.820 126.315 ;
        RECT 126.990 125.395 127.390 125.715 ;
        RECT 126.340 124.785 126.740 125.135 ;
        RECT 126.360 123.955 126.650 124.785 ;
        RECT 127.080 124.535 127.370 125.395 ;
        RECT 128.430 125.135 128.720 125.965 ;
        RECT 129.180 125.715 129.470 126.575 ;
        RECT 130.520 126.325 130.810 127.445 ;
        RECT 131.250 126.895 131.540 128.670 ;
        RECT 132.570 127.445 132.990 127.855 ;
        RECT 131.160 126.575 131.560 126.895 ;
        RECT 130.500 125.975 130.900 126.325 ;
        RECT 129.090 125.395 129.490 125.715 ;
        RECT 128.420 124.785 128.820 125.135 ;
        RECT 126.990 124.215 127.390 124.535 ;
        RECT 126.340 123.605 126.740 123.955 ;
        RECT 126.360 122.775 126.650 123.605 ;
        RECT 127.080 123.355 127.370 124.215 ;
        RECT 128.430 123.955 128.720 124.785 ;
        RECT 129.180 124.535 129.470 125.395 ;
        RECT 130.520 125.135 130.810 125.975 ;
        RECT 131.250 125.715 131.540 126.575 ;
        RECT 132.620 126.325 132.910 127.445 ;
        RECT 133.350 126.895 133.640 128.670 ;
        RECT 135.450 128.180 141.795 128.670 ;
        RECT 134.650 127.445 135.070 127.855 ;
        RECT 133.260 126.575 133.660 126.895 ;
        RECT 132.600 125.975 133.000 126.325 ;
        RECT 131.170 125.395 131.570 125.715 ;
        RECT 130.500 124.785 130.900 125.135 ;
        RECT 129.090 124.215 129.490 124.535 ;
        RECT 128.420 123.605 128.820 123.955 ;
        RECT 126.990 123.035 127.390 123.355 ;
        RECT 114.500 122.445 114.910 122.725 ;
        RECT 113.810 120.105 114.190 120.455 ;
        RECT 108.530 117.815 108.920 118.165 ;
        RECT 108.530 117.735 108.830 117.815 ;
        RECT 113.830 116.350 114.140 120.105 ;
        RECT 114.560 118.145 114.880 122.445 ;
        RECT 126.340 122.425 126.740 122.775 ;
        RECT 126.360 121.595 126.650 122.425 ;
        RECT 127.080 122.175 127.370 123.035 ;
        RECT 128.430 122.775 128.720 123.605 ;
        RECT 129.180 123.355 129.470 124.215 ;
        RECT 130.520 123.955 130.810 124.785 ;
        RECT 131.250 124.525 131.540 125.395 ;
        RECT 132.620 125.135 132.910 125.975 ;
        RECT 133.350 125.715 133.640 126.575 ;
        RECT 134.710 126.315 135.000 127.445 ;
        RECT 135.450 126.885 135.740 128.180 ;
        RECT 135.350 126.565 135.750 126.885 ;
        RECT 145.200 126.865 145.470 129.200 ;
        RECT 145.810 129.035 148.190 129.495 ;
        RECT 145.810 128.725 146.270 129.035 ;
        RECT 145.900 128.145 146.180 128.725 ;
        RECT 145.810 127.835 146.190 128.145 ;
        RECT 134.670 125.965 135.070 126.315 ;
        RECT 133.260 125.395 133.660 125.715 ;
        RECT 132.600 124.785 133.000 125.135 ;
        RECT 131.170 124.205 131.570 124.525 ;
        RECT 130.500 123.605 130.900 123.955 ;
        RECT 129.090 123.035 129.490 123.355 ;
        RECT 128.420 122.425 128.820 122.775 ;
        RECT 126.990 121.855 127.390 122.175 ;
        RECT 126.340 121.245 126.740 121.595 ;
        RECT 126.360 120.675 126.650 121.245 ;
        RECT 127.080 120.995 127.370 121.855 ;
        RECT 128.430 121.595 128.720 122.425 ;
        RECT 129.180 122.175 129.470 123.035 ;
        RECT 130.520 122.775 130.810 123.605 ;
        RECT 131.250 123.355 131.540 124.205 ;
        RECT 132.620 123.955 132.910 124.785 ;
        RECT 133.350 124.535 133.640 125.395 ;
        RECT 134.710 125.135 135.000 125.965 ;
        RECT 135.450 125.715 135.740 126.565 ;
        RECT 145.180 126.545 145.580 126.865 ;
        RECT 135.350 125.395 135.750 125.715 ;
        RECT 134.680 124.785 135.080 125.135 ;
        RECT 133.260 124.215 133.660 124.535 ;
        RECT 132.600 123.605 133.000 123.955 ;
        RECT 131.170 123.035 131.570 123.355 ;
        RECT 130.500 122.425 130.900 122.775 ;
        RECT 129.090 121.855 129.490 122.175 ;
        RECT 128.420 121.245 128.820 121.595 ;
        RECT 126.990 120.675 127.390 120.995 ;
        RECT 117.315 120.160 124.695 120.480 ;
        RECT 126.340 120.160 126.650 120.675 ;
        RECT 127.080 120.645 127.370 120.675 ;
        RECT 128.430 120.160 128.720 121.245 ;
        RECT 129.180 120.995 129.470 121.855 ;
        RECT 130.520 121.585 130.810 122.425 ;
        RECT 131.250 122.175 131.540 123.035 ;
        RECT 132.620 122.775 132.910 123.605 ;
        RECT 133.350 123.355 133.640 124.215 ;
        RECT 134.710 123.955 135.000 124.785 ;
        RECT 135.450 124.535 135.740 125.395 ;
        RECT 135.350 124.215 135.750 124.535 ;
        RECT 145.200 124.285 145.470 126.545 ;
        RECT 145.900 125.575 146.180 127.835 ;
        RECT 145.820 125.265 146.200 125.575 ;
        RECT 134.680 123.605 135.080 123.955 ;
        RECT 133.260 123.035 133.660 123.355 ;
        RECT 132.600 122.425 133.000 122.775 ;
        RECT 131.170 121.855 131.570 122.175 ;
        RECT 130.500 121.235 130.900 121.585 ;
        RECT 129.090 120.675 129.490 120.995 ;
        RECT 129.180 120.645 129.470 120.675 ;
        RECT 130.520 120.645 130.810 121.235 ;
        RECT 131.250 120.995 131.540 121.855 ;
        RECT 132.620 121.595 132.910 122.425 ;
        RECT 133.350 122.175 133.640 123.035 ;
        RECT 134.710 122.785 135.000 123.605 ;
        RECT 135.450 123.355 135.740 124.215 ;
        RECT 145.180 123.965 145.580 124.285 ;
        RECT 135.350 123.035 135.750 123.355 ;
        RECT 134.680 122.435 135.080 122.785 ;
        RECT 133.260 121.855 133.660 122.175 ;
        RECT 132.600 121.245 133.000 121.595 ;
        RECT 131.170 120.675 131.570 120.995 ;
        RECT 131.250 120.645 131.540 120.675 ;
        RECT 132.620 120.665 132.910 121.245 ;
        RECT 133.350 120.985 133.640 121.855 ;
        RECT 134.710 121.595 135.000 122.435 ;
        RECT 135.450 122.175 135.740 123.035 ;
        RECT 135.350 121.855 135.750 122.175 ;
        RECT 134.680 121.245 135.080 121.595 ;
        RECT 133.260 120.665 133.660 120.985 ;
        RECT 134.710 120.675 135.000 121.245 ;
        RECT 135.450 120.995 135.740 121.855 ;
        RECT 145.200 121.705 145.470 123.965 ;
        RECT 145.900 122.985 146.180 125.265 ;
        RECT 145.830 122.675 146.210 122.985 ;
        RECT 145.180 121.385 145.580 121.705 ;
        RECT 135.350 120.675 135.750 120.995 ;
        RECT 130.540 120.160 130.810 120.645 ;
        RECT 132.600 120.160 132.910 120.665 ;
        RECT 133.350 120.645 133.640 120.665 ;
        RECT 134.690 120.645 135.000 120.675 ;
        RECT 135.450 120.645 135.740 120.675 ;
        RECT 134.690 120.160 134.990 120.645 ;
        RECT 145.200 120.360 145.470 121.385 ;
        RECT 145.900 121.355 146.180 122.675 ;
        RECT 117.315 119.805 135.020 120.160 ;
        RECT 117.315 119.510 124.695 119.805 ;
        RECT 114.510 117.865 114.920 118.145 ;
        RECT 111.185 116.040 114.140 116.350 ;
        RECT 112.660 116.035 114.140 116.040 ;
        RECT 114.560 116.425 114.880 117.865 ;
        RECT 117.315 116.750 118.285 119.510 ;
        RECT 126.340 119.365 126.650 119.805 ;
        RECT 126.340 118.755 126.620 119.365 ;
        RECT 127.100 119.355 127.380 119.415 ;
        RECT 128.430 119.375 128.720 119.805 ;
        RECT 130.540 119.415 130.810 119.805 ;
        RECT 127.000 119.035 127.390 119.355 ;
        RECT 126.340 118.455 126.750 118.755 ;
        RECT 126.340 117.575 126.620 118.455 ;
        RECT 127.100 118.175 127.380 119.035 ;
        RECT 128.440 118.755 128.720 119.375 ;
        RECT 129.190 119.355 129.470 119.415 ;
        RECT 129.100 119.035 129.490 119.355 ;
        RECT 128.440 118.455 128.840 118.755 ;
        RECT 127.000 117.855 127.390 118.175 ;
        RECT 126.340 117.275 126.750 117.575 ;
        RECT 115.535 116.425 118.285 116.750 ;
        RECT 114.560 116.105 118.285 116.425 ;
        RECT 114.560 116.035 114.880 116.105 ;
        RECT 109.160 114.765 111.685 115.295 ;
        RECT 108.550 113.695 108.820 113.735 ;
        RECT 108.530 113.365 108.890 113.695 ;
        RECT 108.550 109.115 108.820 113.365 ;
        RECT 109.290 111.415 109.560 114.765 ;
        RECT 111.155 113.135 111.685 114.765 ;
        RECT 112.660 114.730 114.085 116.035 ;
        RECT 115.535 115.780 118.285 116.105 ;
        RECT 123.250 114.730 124.675 117.005 ;
        RECT 112.660 113.305 124.675 114.730 ;
        RECT 126.340 116.395 126.620 117.275 ;
        RECT 127.100 116.995 127.380 117.855 ;
        RECT 128.440 117.575 128.720 118.455 ;
        RECT 129.190 118.175 129.470 119.035 ;
        RECT 130.540 118.755 130.820 119.415 ;
        RECT 131.280 119.355 131.560 119.415 ;
        RECT 132.600 119.375 132.910 119.805 ;
        RECT 131.180 119.035 131.570 119.355 ;
        RECT 130.520 118.455 130.920 118.755 ;
        RECT 129.100 117.855 129.490 118.175 ;
        RECT 128.440 117.275 128.840 117.575 ;
        RECT 127.000 116.675 127.390 116.995 ;
        RECT 126.340 116.095 126.750 116.395 ;
        RECT 126.340 115.205 126.620 116.095 ;
        RECT 127.100 115.815 127.380 116.675 ;
        RECT 128.440 116.395 128.720 117.275 ;
        RECT 129.190 116.995 129.470 117.855 ;
        RECT 130.540 117.575 130.820 118.455 ;
        RECT 131.280 118.175 131.560 119.035 ;
        RECT 132.600 118.755 132.880 119.375 ;
        RECT 133.370 119.355 133.650 119.415 ;
        RECT 133.260 119.035 133.650 119.355 ;
        RECT 132.580 118.455 132.980 118.755 ;
        RECT 131.180 117.855 131.570 118.175 ;
        RECT 130.520 117.275 130.920 117.575 ;
        RECT 129.100 116.675 129.490 116.995 ;
        RECT 128.440 116.095 128.840 116.395 ;
        RECT 127.000 115.495 127.390 115.815 ;
        RECT 126.340 114.905 126.750 115.205 ;
        RECT 126.340 114.035 126.620 114.905 ;
        RECT 127.100 114.645 127.380 115.495 ;
        RECT 128.440 115.215 128.720 116.095 ;
        RECT 129.190 115.815 129.470 116.675 ;
        RECT 130.540 116.395 130.820 117.275 ;
        RECT 131.280 116.985 131.560 117.855 ;
        RECT 132.600 117.575 132.880 118.455 ;
        RECT 133.370 118.175 133.650 119.035 ;
        RECT 134.690 119.375 134.990 119.805 ;
        RECT 134.690 118.755 134.970 119.375 ;
        RECT 135.460 119.355 135.740 119.415 ;
        RECT 135.350 119.035 135.740 119.355 ;
        RECT 134.680 118.455 135.080 118.755 ;
        RECT 133.260 117.855 133.650 118.175 ;
        RECT 132.580 117.275 132.980 117.575 ;
        RECT 131.180 116.665 131.570 116.985 ;
        RECT 130.520 116.095 130.920 116.395 ;
        RECT 129.100 115.495 129.490 115.815 ;
        RECT 128.440 114.915 128.840 115.215 ;
        RECT 127.000 114.325 127.390 114.645 ;
        RECT 126.340 113.735 126.750 114.035 ;
        RECT 111.150 112.115 111.690 113.135 ;
        RECT 126.340 112.400 126.620 113.735 ;
        RECT 127.100 113.455 127.380 114.325 ;
        RECT 128.440 114.035 128.720 114.915 ;
        RECT 129.190 114.635 129.470 115.495 ;
        RECT 130.540 115.215 130.820 116.095 ;
        RECT 131.280 115.815 131.560 116.665 ;
        RECT 132.600 116.395 132.880 117.275 ;
        RECT 133.370 116.995 133.650 117.855 ;
        RECT 134.690 117.575 134.970 118.455 ;
        RECT 135.460 118.175 135.740 119.035 ;
        RECT 145.160 118.365 145.430 118.425 ;
        RECT 135.350 117.855 135.740 118.175 ;
        RECT 145.140 118.045 145.540 118.365 ;
        RECT 134.680 117.275 135.080 117.575 ;
        RECT 133.260 116.675 133.650 116.995 ;
        RECT 132.580 116.095 132.980 116.395 ;
        RECT 131.180 115.495 131.570 115.815 ;
        RECT 130.520 114.915 130.920 115.215 ;
        RECT 129.100 114.315 129.490 114.635 ;
        RECT 128.440 113.735 128.840 114.035 ;
        RECT 127.000 113.135 127.390 113.455 ;
        RECT 111.150 112.105 112.015 112.115 ;
        RECT 116.580 112.105 117.445 112.135 ;
        RECT 109.210 111.085 109.570 111.415 ;
        RECT 111.150 111.240 117.445 112.105 ;
        RECT 108.530 108.785 108.890 109.115 ;
        RECT 108.550 104.535 108.820 108.785 ;
        RECT 109.290 106.825 109.560 111.085 ;
        RECT 114.140 109.645 114.820 111.240 ;
        RECT 116.580 111.210 117.445 111.240 ;
        RECT 126.315 110.645 126.650 112.400 ;
        RECT 127.100 112.025 127.380 113.135 ;
        RECT 128.440 112.535 128.720 113.735 ;
        RECT 129.190 113.455 129.470 114.315 ;
        RECT 130.540 114.035 130.820 114.915 ;
        RECT 131.280 114.635 131.560 115.495 ;
        RECT 132.600 115.215 132.880 116.095 ;
        RECT 133.370 115.815 133.650 116.675 ;
        RECT 134.690 116.395 134.970 117.275 ;
        RECT 135.460 116.995 135.740 117.855 ;
        RECT 135.350 116.675 135.740 116.995 ;
        RECT 134.680 116.095 135.080 116.395 ;
        RECT 133.260 115.495 133.650 115.815 ;
        RECT 132.580 114.915 132.980 115.215 ;
        RECT 131.180 114.315 131.570 114.635 ;
        RECT 130.520 113.735 130.920 114.035 ;
        RECT 129.100 113.135 129.490 113.455 ;
        RECT 128.380 112.135 128.780 112.535 ;
        RECT 127.105 111.260 127.380 112.025 ;
        RECT 129.190 111.260 129.470 113.135 ;
        RECT 130.540 112.545 130.820 113.735 ;
        RECT 131.280 113.455 131.560 114.315 ;
        RECT 132.600 114.035 132.880 114.915 ;
        RECT 133.370 114.635 133.650 115.495 ;
        RECT 134.690 115.215 134.970 116.095 ;
        RECT 135.460 115.815 135.740 116.675 ;
        RECT 135.350 115.495 135.740 115.815 ;
        RECT 145.160 115.795 145.430 118.045 ;
        RECT 145.900 117.085 146.180 118.415 ;
        RECT 145.830 116.775 146.210 117.085 ;
        RECT 134.680 114.915 135.080 115.215 ;
        RECT 133.260 114.315 133.650 114.635 ;
        RECT 132.580 113.735 132.980 114.035 ;
        RECT 131.190 113.135 131.580 113.455 ;
        RECT 130.470 112.135 130.880 112.545 ;
        RECT 131.280 111.260 131.560 113.135 ;
        RECT 132.600 112.545 132.880 113.735 ;
        RECT 133.370 113.455 133.650 114.315 ;
        RECT 134.690 114.035 134.970 114.915 ;
        RECT 135.460 114.635 135.740 115.495 ;
        RECT 145.140 115.475 145.540 115.795 ;
        RECT 135.350 114.315 135.740 114.635 ;
        RECT 134.680 113.735 135.080 114.035 ;
        RECT 133.260 113.135 133.650 113.455 ;
        RECT 132.540 112.135 132.950 112.545 ;
        RECT 133.370 111.260 133.650 113.135 ;
        RECT 134.690 112.530 134.970 113.735 ;
        RECT 135.460 113.455 135.740 114.315 ;
        RECT 135.350 113.135 135.740 113.455 ;
        RECT 145.160 113.205 145.430 115.475 ;
        RECT 145.900 114.495 146.180 116.775 ;
        RECT 145.830 114.185 146.210 114.495 ;
        RECT 134.680 112.140 134.980 112.530 ;
        RECT 135.460 111.750 135.740 113.135 ;
        RECT 145.140 112.885 145.540 113.205 ;
        RECT 135.460 111.260 141.875 111.750 ;
        RECT 127.105 111.155 141.875 111.260 ;
        RECT 127.090 111.020 141.875 111.155 ;
        RECT 127.090 110.985 135.740 111.020 ;
        RECT 126.295 110.360 126.670 110.645 ;
        RECT 126.315 110.335 126.650 110.360 ;
        RECT 120.425 109.955 121.175 109.975 ;
        RECT 127.090 109.955 127.890 110.985 ;
        RECT 135.460 110.955 135.740 110.985 ;
        RECT 141.145 110.790 141.875 111.020 ;
        RECT 141.145 110.560 144.375 110.790 ;
        RECT 145.160 110.560 145.430 112.885 ;
        RECT 145.900 111.915 146.180 114.185 ;
        RECT 145.830 111.605 146.210 111.915 ;
        RECT 145.900 111.050 146.180 111.605 ;
        RECT 141.145 110.290 145.430 110.560 ;
        RECT 145.805 110.715 146.280 111.050 ;
        RECT 141.145 110.060 144.375 110.290 ;
        RECT 145.805 110.240 148.195 110.715 ;
        RECT 114.290 107.425 114.670 109.645 ;
        RECT 118.400 109.155 121.200 109.955 ;
        RECT 126.445 109.155 127.890 109.955 ;
        RECT 120.425 109.135 121.175 109.155 ;
        RECT 120.095 108.475 144.230 108.925 ;
        RECT 114.230 107.085 114.750 107.425 ;
        RECT 109.210 106.495 109.570 106.825 ;
        RECT 108.530 104.205 108.890 104.535 ;
        RECT 108.550 99.955 108.820 104.205 ;
        RECT 109.290 102.255 109.560 106.495 ;
        RECT 114.290 106.245 114.670 107.085 ;
        RECT 115.750 106.505 116.270 106.805 ;
        RECT 114.230 105.905 114.750 106.245 ;
        RECT 114.290 105.055 114.670 105.905 ;
        RECT 115.840 105.625 116.220 106.505 ;
        RECT 120.095 105.850 120.545 108.475 ;
        RECT 121.680 106.535 122.130 108.475 ;
        RECT 123.710 107.475 124.240 107.815 ;
        RECT 121.650 106.165 122.260 106.535 ;
        RECT 118.605 105.835 120.545 105.850 ;
        RECT 115.750 105.325 116.270 105.625 ;
        RECT 114.230 104.715 114.750 105.055 ;
        RECT 114.290 103.875 114.670 104.715 ;
        RECT 115.840 104.455 116.220 105.325 ;
        RECT 117.860 105.025 120.560 105.835 ;
        RECT 117.860 104.995 119.060 105.025 ;
        RECT 115.750 104.155 116.270 104.455 ;
        RECT 114.230 103.535 114.750 103.875 ;
        RECT 114.290 102.695 114.670 103.535 ;
        RECT 115.840 103.275 116.220 104.155 ;
        RECT 115.750 102.975 116.270 103.275 ;
        RECT 114.230 102.355 114.750 102.695 ;
        RECT 109.210 101.925 109.570 102.255 ;
        RECT 108.530 99.625 108.890 99.955 ;
        RECT 108.550 95.375 108.820 99.625 ;
        RECT 109.290 97.675 109.560 101.925 ;
        RECT 114.290 101.515 114.670 102.355 ;
        RECT 115.840 102.095 116.220 102.975 ;
        RECT 115.750 101.795 116.270 102.095 ;
        RECT 114.230 101.175 114.750 101.515 ;
        RECT 114.290 100.335 114.670 101.175 ;
        RECT 115.840 100.915 116.220 101.795 ;
        RECT 115.750 100.615 116.270 100.915 ;
        RECT 114.230 99.995 114.750 100.335 ;
        RECT 114.290 99.155 114.670 99.995 ;
        RECT 115.840 99.735 116.220 100.615 ;
        RECT 115.750 99.435 116.270 99.735 ;
        RECT 112.085 98.050 113.020 98.925 ;
        RECT 114.240 98.815 114.760 99.155 ;
        RECT 109.210 97.345 109.570 97.675 ;
        RECT 108.530 95.045 108.890 95.375 ;
        RECT 108.550 90.795 108.820 95.045 ;
        RECT 109.290 93.085 109.560 97.345 ;
        RECT 109.210 92.755 109.570 93.085 ;
        RECT 108.530 90.465 108.890 90.795 ;
        RECT 108.550 89.685 108.820 90.465 ;
        RECT 107.150 89.670 108.860 89.685 ;
        RECT 107.150 89.340 109.000 89.670 ;
        RECT 108.125 89.195 109.000 89.340 ;
        RECT 112.115 89.195 112.990 98.050 ;
        RECT 114.290 97.975 114.670 98.815 ;
        RECT 115.840 98.555 116.220 99.435 ;
        RECT 115.750 98.255 116.270 98.555 ;
        RECT 114.240 97.635 114.760 97.975 ;
        RECT 114.290 96.795 114.670 97.635 ;
        RECT 115.840 97.375 116.220 98.255 ;
        RECT 115.750 97.075 116.270 97.375 ;
        RECT 114.240 96.455 114.760 96.795 ;
        RECT 114.290 95.615 114.670 96.455 ;
        RECT 115.840 96.195 116.220 97.075 ;
        RECT 115.750 95.895 116.270 96.195 ;
        RECT 114.240 95.275 114.760 95.615 ;
        RECT 115.840 94.275 116.220 95.895 ;
        RECT 117.860 94.275 118.950 104.995 ;
        RECT 121.680 103.955 122.130 106.165 ;
        RECT 123.810 105.235 124.190 107.475 ;
        RECT 125.360 106.535 125.810 108.475 ;
        RECT 127.350 107.475 127.880 107.815 ;
        RECT 125.300 106.165 125.910 106.535 ;
        RECT 123.710 104.895 124.240 105.235 ;
        RECT 121.650 103.585 122.260 103.955 ;
        RECT 121.680 101.365 122.130 103.585 ;
        RECT 123.810 102.645 124.190 104.895 ;
        RECT 125.360 103.955 125.810 106.165 ;
        RECT 127.460 105.235 127.840 107.475 ;
        RECT 129.050 106.535 129.500 108.475 ;
        RECT 131.100 107.475 131.630 107.815 ;
        RECT 129.010 106.165 129.620 106.535 ;
        RECT 127.350 104.895 127.880 105.235 ;
        RECT 125.320 103.585 125.930 103.955 ;
        RECT 123.710 102.305 124.240 102.645 ;
        RECT 121.650 100.995 122.260 101.365 ;
        RECT 121.680 98.805 122.130 100.995 ;
        RECT 123.810 100.075 124.190 102.305 ;
        RECT 125.360 101.375 125.810 103.585 ;
        RECT 127.460 102.655 127.840 104.895 ;
        RECT 129.050 103.955 129.500 106.165 ;
        RECT 131.200 105.235 131.580 107.475 ;
        RECT 132.730 106.535 133.180 108.475 ;
        RECT 134.740 107.475 135.270 107.815 ;
        RECT 132.680 106.165 133.290 106.535 ;
        RECT 131.100 104.895 131.630 105.235 ;
        RECT 129.010 103.585 129.620 103.955 ;
        RECT 127.350 102.315 127.880 102.655 ;
        RECT 125.300 101.005 125.910 101.375 ;
        RECT 123.710 99.735 124.240 100.075 ;
        RECT 121.610 98.435 122.220 98.805 ;
        RECT 121.680 96.215 122.130 98.435 ;
        RECT 123.810 97.495 124.190 99.735 ;
        RECT 125.360 98.795 125.810 101.005 ;
        RECT 127.460 100.075 127.840 102.315 ;
        RECT 129.050 101.375 129.500 103.585 ;
        RECT 131.200 102.665 131.580 104.895 ;
        RECT 132.730 103.975 133.180 106.165 ;
        RECT 134.840 105.235 135.220 107.475 ;
        RECT 136.420 106.545 136.870 108.475 ;
        RECT 138.450 107.475 138.980 107.815 ;
        RECT 136.390 106.175 137.000 106.545 ;
        RECT 134.740 104.895 135.270 105.235 ;
        RECT 132.680 103.605 133.290 103.975 ;
        RECT 131.100 102.325 131.630 102.665 ;
        RECT 128.980 101.005 129.590 101.375 ;
        RECT 127.350 99.735 127.880 100.075 ;
        RECT 125.320 98.425 125.930 98.795 ;
        RECT 123.720 97.155 124.250 97.495 ;
        RECT 121.650 95.845 122.260 96.215 ;
        RECT 115.840 93.835 118.950 94.275 ;
        RECT 115.845 93.820 118.950 93.835 ;
        RECT 108.125 88.320 112.990 89.195 ;
        RECT 117.880 93.455 118.950 93.820 ;
        RECT 121.680 93.635 122.130 95.845 ;
        RECT 123.810 94.905 124.190 97.155 ;
        RECT 125.360 96.205 125.810 98.425 ;
        RECT 127.460 97.495 127.840 99.735 ;
        RECT 129.050 98.795 129.500 101.005 ;
        RECT 131.200 100.075 131.580 102.325 ;
        RECT 132.730 101.385 133.180 103.605 ;
        RECT 134.840 102.655 135.220 104.895 ;
        RECT 136.420 103.965 136.870 106.175 ;
        RECT 138.550 105.235 138.930 107.475 ;
        RECT 140.090 106.545 140.540 108.475 ;
        RECT 142.090 107.475 142.620 107.815 ;
        RECT 140.060 106.175 140.670 106.545 ;
        RECT 138.450 104.895 138.980 105.235 ;
        RECT 136.390 103.595 137.000 103.965 ;
        RECT 134.740 102.315 135.270 102.655 ;
        RECT 132.670 101.015 133.280 101.385 ;
        RECT 131.100 99.735 131.630 100.075 ;
        RECT 129.010 98.425 129.620 98.795 ;
        RECT 127.350 97.155 127.880 97.495 ;
        RECT 125.340 95.835 125.950 96.205 ;
        RECT 123.720 94.565 124.250 94.905 ;
        RECT 108.500 87.045 108.980 87.415 ;
        RECT 108.530 82.815 108.900 87.045 ;
        RECT 109.250 85.105 109.600 87.395 ;
        RECT 109.150 84.715 109.620 85.105 ;
        RECT 108.500 82.445 108.980 82.815 ;
        RECT 108.530 78.235 108.900 82.445 ;
        RECT 109.250 80.535 109.600 84.715 ;
        RECT 109.150 80.145 109.620 80.535 ;
        RECT 117.880 80.155 118.960 93.455 ;
        RECT 121.650 93.265 122.260 93.635 ;
        RECT 121.680 91.055 122.130 93.265 ;
        RECT 123.810 92.335 124.190 94.565 ;
        RECT 125.360 93.635 125.810 95.835 ;
        RECT 127.460 94.915 127.840 97.155 ;
        RECT 129.050 96.215 129.500 98.425 ;
        RECT 131.200 97.495 131.580 99.735 ;
        RECT 132.730 98.805 133.180 101.015 ;
        RECT 134.840 100.075 135.220 102.315 ;
        RECT 136.420 101.365 136.870 103.595 ;
        RECT 138.550 102.655 138.930 104.895 ;
        RECT 140.090 103.965 140.540 106.175 ;
        RECT 142.190 105.235 142.570 107.475 ;
        RECT 143.780 106.535 144.230 108.475 ;
        RECT 145.780 107.475 146.310 107.815 ;
        RECT 143.740 106.165 144.350 106.535 ;
        RECT 142.090 104.895 142.620 105.235 ;
        RECT 140.060 103.595 140.670 103.965 ;
        RECT 138.450 102.315 138.980 102.655 ;
        RECT 136.390 100.995 137.000 101.365 ;
        RECT 134.740 99.735 135.270 100.075 ;
        RECT 132.690 98.435 133.300 98.805 ;
        RECT 131.100 97.155 131.630 97.495 ;
        RECT 129.000 95.845 129.610 96.215 ;
        RECT 127.350 94.575 127.880 94.915 ;
        RECT 125.320 93.265 125.930 93.635 ;
        RECT 123.720 91.995 124.250 92.335 ;
        RECT 121.640 90.685 122.250 91.055 ;
        RECT 121.680 88.475 122.130 90.685 ;
        RECT 123.810 89.745 124.190 91.995 ;
        RECT 125.360 91.055 125.810 93.265 ;
        RECT 127.460 92.345 127.840 94.575 ;
        RECT 129.050 93.635 129.500 95.845 ;
        RECT 131.200 94.915 131.580 97.155 ;
        RECT 132.730 96.215 133.180 98.435 ;
        RECT 134.840 97.495 135.220 99.735 ;
        RECT 136.420 98.805 136.870 100.995 ;
        RECT 138.550 100.075 138.930 102.315 ;
        RECT 140.090 101.365 140.540 103.595 ;
        RECT 142.190 102.645 142.570 104.895 ;
        RECT 143.780 103.955 144.230 106.165 ;
        RECT 145.880 105.225 146.260 107.475 ;
        RECT 145.780 104.885 146.310 105.225 ;
        RECT 143.740 103.585 144.350 103.955 ;
        RECT 142.090 102.305 142.620 102.645 ;
        RECT 140.060 100.995 140.670 101.365 ;
        RECT 138.450 99.735 138.980 100.075 ;
        RECT 136.390 98.435 137.000 98.805 ;
        RECT 134.740 97.155 135.270 97.495 ;
        RECT 132.680 95.845 133.290 96.215 ;
        RECT 131.100 94.575 131.630 94.915 ;
        RECT 129.000 93.265 129.610 93.635 ;
        RECT 127.350 92.005 127.880 92.345 ;
        RECT 125.330 90.685 125.940 91.055 ;
        RECT 123.720 89.405 124.250 89.745 ;
        RECT 121.630 88.105 122.240 88.475 ;
        RECT 121.680 85.895 122.130 88.105 ;
        RECT 123.810 87.175 124.190 89.405 ;
        RECT 125.360 88.475 125.810 90.685 ;
        RECT 127.460 89.755 127.840 92.005 ;
        RECT 129.050 91.055 129.500 93.265 ;
        RECT 131.200 92.335 131.580 94.575 ;
        RECT 132.730 93.645 133.180 95.845 ;
        RECT 134.840 94.915 135.220 97.155 ;
        RECT 136.420 96.215 136.870 98.435 ;
        RECT 138.550 97.495 138.930 99.735 ;
        RECT 140.090 98.805 140.540 100.995 ;
        RECT 142.190 100.075 142.570 102.305 ;
        RECT 143.780 101.375 144.230 103.585 ;
        RECT 145.880 102.645 146.260 104.885 ;
        RECT 145.780 102.305 146.310 102.645 ;
        RECT 143.740 101.005 144.350 101.375 ;
        RECT 142.090 99.735 142.620 100.075 ;
        RECT 140.060 98.435 140.670 98.805 ;
        RECT 138.450 97.155 138.980 97.495 ;
        RECT 136.390 95.845 137.000 96.215 ;
        RECT 134.740 94.575 135.270 94.915 ;
        RECT 132.680 93.275 133.290 93.645 ;
        RECT 131.100 91.995 131.630 92.335 ;
        RECT 129.000 90.685 129.610 91.055 ;
        RECT 127.350 89.415 127.880 89.755 ;
        RECT 125.320 88.105 125.930 88.475 ;
        RECT 123.720 86.835 124.250 87.175 ;
        RECT 121.640 85.525 122.250 85.895 ;
        RECT 121.680 83.315 122.130 85.525 ;
        RECT 123.810 84.595 124.190 86.835 ;
        RECT 125.360 85.885 125.810 88.105 ;
        RECT 127.460 87.175 127.840 89.415 ;
        RECT 129.050 88.475 129.500 90.685 ;
        RECT 131.200 89.755 131.580 91.995 ;
        RECT 132.730 91.065 133.180 93.275 ;
        RECT 134.840 92.335 135.220 94.575 ;
        RECT 136.420 93.655 136.870 95.845 ;
        RECT 138.550 94.915 138.930 97.155 ;
        RECT 140.090 96.215 140.540 98.435 ;
        RECT 142.190 97.495 142.570 99.735 ;
        RECT 143.780 98.795 144.230 101.005 ;
        RECT 145.880 100.065 146.260 102.305 ;
        RECT 145.780 99.725 146.310 100.065 ;
        RECT 143.740 98.425 144.350 98.795 ;
        RECT 142.090 97.155 142.620 97.495 ;
        RECT 140.060 95.845 140.670 96.215 ;
        RECT 138.450 94.575 138.980 94.915 ;
        RECT 136.390 93.285 137.000 93.655 ;
        RECT 134.740 91.995 135.270 92.335 ;
        RECT 132.690 90.695 133.300 91.065 ;
        RECT 131.100 89.415 131.630 89.755 ;
        RECT 129.000 88.105 129.610 88.475 ;
        RECT 127.350 86.835 127.880 87.175 ;
        RECT 125.320 85.515 125.930 85.885 ;
        RECT 123.720 84.255 124.250 84.595 ;
        RECT 121.640 82.945 122.250 83.315 ;
        RECT 121.680 81.535 122.130 82.945 ;
        RECT 123.810 82.005 124.190 84.255 ;
        RECT 125.360 83.325 125.810 85.515 ;
        RECT 127.460 84.595 127.840 86.835 ;
        RECT 129.050 85.895 129.500 88.105 ;
        RECT 131.200 87.175 131.580 89.415 ;
        RECT 132.730 88.475 133.180 90.695 ;
        RECT 134.840 89.755 135.220 91.995 ;
        RECT 136.420 91.055 136.870 93.285 ;
        RECT 138.550 92.335 138.930 94.575 ;
        RECT 140.090 93.645 140.540 95.845 ;
        RECT 142.190 94.915 142.570 97.155 ;
        RECT 143.780 96.215 144.230 98.425 ;
        RECT 145.880 97.485 146.260 99.725 ;
        RECT 145.780 97.145 146.310 97.485 ;
        RECT 143.740 95.845 144.350 96.215 ;
        RECT 142.090 94.575 142.620 94.915 ;
        RECT 140.060 93.275 140.670 93.645 ;
        RECT 138.450 91.995 138.980 92.335 ;
        RECT 136.390 90.685 137.000 91.055 ;
        RECT 134.740 89.415 135.270 89.755 ;
        RECT 132.670 88.105 133.280 88.475 ;
        RECT 131.100 86.835 131.630 87.175 ;
        RECT 128.990 85.525 129.600 85.895 ;
        RECT 127.350 84.255 127.880 84.595 ;
        RECT 125.320 82.955 125.930 83.325 ;
        RECT 123.720 81.665 124.250 82.005 ;
        RECT 123.810 80.825 124.190 81.665 ;
        RECT 125.360 81.535 125.810 82.955 ;
        RECT 127.460 82.005 127.840 84.255 ;
        RECT 129.050 83.315 129.500 85.525 ;
        RECT 131.200 84.595 131.580 86.835 ;
        RECT 132.730 85.895 133.180 88.105 ;
        RECT 134.840 87.165 135.220 89.415 ;
        RECT 136.420 88.465 136.870 90.685 ;
        RECT 138.550 89.755 138.930 91.995 ;
        RECT 140.090 91.055 140.540 93.275 ;
        RECT 142.190 92.335 142.570 94.575 ;
        RECT 143.780 93.635 144.230 95.845 ;
        RECT 145.880 94.905 146.260 97.145 ;
        RECT 145.780 94.565 146.310 94.905 ;
        RECT 143.740 93.265 144.350 93.635 ;
        RECT 142.090 91.995 142.620 92.335 ;
        RECT 140.060 90.685 140.670 91.055 ;
        RECT 138.450 89.415 138.980 89.755 ;
        RECT 136.390 88.095 137.000 88.465 ;
        RECT 134.740 86.825 135.270 87.165 ;
        RECT 132.680 85.525 133.290 85.895 ;
        RECT 131.100 84.255 131.630 84.595 ;
        RECT 129.000 82.945 129.610 83.315 ;
        RECT 127.350 81.665 127.880 82.005 ;
        RECT 127.460 80.825 127.840 81.665 ;
        RECT 129.050 81.545 129.500 82.945 ;
        RECT 131.200 82.005 131.580 84.255 ;
        RECT 132.730 83.315 133.180 85.525 ;
        RECT 134.840 84.585 135.220 86.825 ;
        RECT 136.420 85.895 136.870 88.095 ;
        RECT 138.550 87.175 138.930 89.415 ;
        RECT 140.090 88.465 140.540 90.685 ;
        RECT 142.190 89.755 142.570 91.995 ;
        RECT 143.780 91.065 144.230 93.265 ;
        RECT 145.880 92.325 146.260 94.565 ;
        RECT 145.780 91.985 146.310 92.325 ;
        RECT 143.740 90.695 144.350 91.065 ;
        RECT 142.100 89.415 142.630 89.755 ;
        RECT 140.060 88.095 140.670 88.465 ;
        RECT 138.450 86.835 138.980 87.175 ;
        RECT 136.390 85.525 137.000 85.895 ;
        RECT 134.740 84.245 135.270 84.585 ;
        RECT 132.690 82.945 133.300 83.315 ;
        RECT 131.100 81.665 131.630 82.005 ;
        RECT 131.200 80.825 131.580 81.665 ;
        RECT 132.730 81.545 133.180 82.945 ;
        RECT 134.840 82.005 135.220 84.245 ;
        RECT 136.420 83.315 136.870 85.525 ;
        RECT 138.550 84.595 138.930 86.835 ;
        RECT 140.090 85.885 140.540 88.095 ;
        RECT 142.190 87.175 142.570 89.415 ;
        RECT 143.780 88.475 144.230 90.695 ;
        RECT 145.880 89.745 146.260 91.985 ;
        RECT 145.780 89.405 146.310 89.745 ;
        RECT 143.750 88.105 144.360 88.475 ;
        RECT 142.100 86.835 142.630 87.175 ;
        RECT 140.060 85.515 140.670 85.885 ;
        RECT 138.450 84.255 138.980 84.595 ;
        RECT 136.390 82.945 137.000 83.315 ;
        RECT 134.740 81.665 135.270 82.005 ;
        RECT 134.840 80.825 135.220 81.665 ;
        RECT 136.420 81.545 136.870 82.945 ;
        RECT 138.550 82.015 138.930 84.255 ;
        RECT 140.090 83.305 140.540 85.515 ;
        RECT 142.190 84.595 142.570 86.835 ;
        RECT 143.780 85.895 144.230 88.105 ;
        RECT 145.880 87.175 146.260 89.405 ;
        RECT 145.780 86.835 146.310 87.175 ;
        RECT 143.750 85.525 144.360 85.895 ;
        RECT 142.100 84.255 142.630 84.595 ;
        RECT 140.060 82.935 140.670 83.305 ;
        RECT 138.450 81.675 138.980 82.015 ;
        RECT 138.550 80.825 138.930 81.675 ;
        RECT 140.090 81.545 140.540 82.935 ;
        RECT 142.190 82.005 142.570 84.255 ;
        RECT 143.780 83.305 144.230 85.525 ;
        RECT 145.880 84.585 146.260 86.835 ;
        RECT 145.780 84.245 146.310 84.585 ;
        RECT 143.770 82.935 144.380 83.305 ;
        RECT 142.100 81.665 142.630 82.005 ;
        RECT 142.190 80.825 142.570 81.665 ;
        RECT 143.780 81.555 144.230 82.935 ;
        RECT 145.880 82.005 146.260 84.245 ;
        RECT 145.780 81.665 146.310 82.005 ;
        RECT 145.880 80.825 146.260 81.665 ;
        RECT 123.810 80.445 146.260 80.825 ;
        RECT 108.500 77.865 108.980 78.235 ;
        RECT 108.530 73.655 108.900 77.865 ;
        RECT 109.250 75.955 109.600 80.145 ;
        RECT 117.850 79.075 118.990 80.155 ;
        RECT 123.810 78.785 124.190 80.445 ;
        RECT 127.460 78.785 127.840 80.445 ;
        RECT 131.200 78.785 131.580 80.445 ;
        RECT 123.810 78.750 131.580 78.785 ;
        RECT 134.840 78.750 135.220 80.445 ;
        RECT 138.550 78.750 138.930 80.445 ;
        RECT 142.190 78.750 142.570 80.445 ;
        RECT 145.880 79.950 146.260 80.445 ;
        RECT 145.735 79.275 148.155 79.950 ;
        RECT 145.880 78.750 146.260 79.275 ;
        RECT 123.810 78.405 146.260 78.750 ;
        RECT 121.690 76.205 122.150 77.495 ;
        RECT 123.810 77.455 124.190 78.405 ;
        RECT 123.720 77.115 124.250 77.455 ;
        RECT 109.150 75.565 109.620 75.955 ;
        RECT 121.630 75.805 122.250 76.205 ;
        RECT 108.500 73.285 108.980 73.655 ;
        RECT 108.530 69.075 108.900 73.285 ;
        RECT 109.250 71.385 109.600 75.565 ;
        RECT 121.690 73.615 122.150 75.805 ;
        RECT 123.810 74.865 124.190 77.115 ;
        RECT 125.370 76.195 125.830 77.495 ;
        RECT 127.460 77.455 127.840 78.405 ;
        RECT 131.200 78.380 146.260 78.405 ;
        RECT 127.350 77.115 127.880 77.455 ;
        RECT 125.320 75.795 125.940 76.195 ;
        RECT 123.720 74.525 124.250 74.865 ;
        RECT 121.630 73.215 122.250 73.615 ;
        RECT 109.150 70.995 109.620 71.385 ;
        RECT 121.690 71.025 122.150 73.215 ;
        RECT 123.810 72.295 124.190 74.525 ;
        RECT 125.370 73.605 125.830 75.795 ;
        RECT 127.460 74.875 127.840 77.115 ;
        RECT 129.050 76.195 129.510 77.495 ;
        RECT 131.200 77.455 131.580 78.380 ;
        RECT 131.100 77.115 131.630 77.455 ;
        RECT 129.010 75.795 129.630 76.195 ;
        RECT 127.360 74.535 127.890 74.875 ;
        RECT 125.300 73.205 125.920 73.605 ;
        RECT 123.720 71.955 124.250 72.295 ;
        RECT 108.500 68.705 108.980 69.075 ;
        RECT 108.530 64.495 108.900 68.705 ;
        RECT 109.250 66.785 109.600 70.995 ;
        RECT 121.620 70.625 122.240 71.025 ;
        RECT 121.690 68.455 122.150 70.625 ;
        RECT 123.810 69.715 124.190 71.955 ;
        RECT 125.370 71.035 125.830 73.205 ;
        RECT 127.460 72.295 127.840 74.535 ;
        RECT 129.050 73.605 129.510 75.795 ;
        RECT 131.200 74.885 131.580 77.115 ;
        RECT 132.740 76.195 133.200 77.495 ;
        RECT 134.840 77.455 135.220 78.380 ;
        RECT 134.740 77.115 135.270 77.455 ;
        RECT 132.690 75.795 133.310 76.195 ;
        RECT 131.100 74.545 131.630 74.885 ;
        RECT 128.990 73.205 129.610 73.605 ;
        RECT 127.360 71.955 127.890 72.295 ;
        RECT 125.320 70.635 125.940 71.035 ;
        RECT 123.720 69.375 124.250 69.715 ;
        RECT 121.640 68.055 122.260 68.455 ;
        RECT 109.150 66.395 109.620 66.785 ;
        RECT 108.500 64.125 108.980 64.495 ;
        RECT 108.530 63.495 108.900 64.125 ;
        RECT 109.250 63.715 109.600 66.395 ;
        RECT 121.690 65.875 122.150 68.055 ;
        RECT 123.810 67.135 124.190 69.375 ;
        RECT 125.370 68.455 125.830 70.635 ;
        RECT 127.460 69.715 127.840 71.955 ;
        RECT 129.050 71.025 129.510 73.205 ;
        RECT 131.200 72.295 131.580 74.545 ;
        RECT 132.740 73.605 133.200 75.795 ;
        RECT 134.840 74.875 135.220 77.115 ;
        RECT 136.410 76.195 136.870 77.495 ;
        RECT 138.550 77.445 138.930 78.380 ;
        RECT 138.440 77.105 138.970 77.445 ;
        RECT 136.360 75.795 136.980 76.195 ;
        RECT 134.740 74.535 135.270 74.875 ;
        RECT 132.690 73.205 133.310 73.605 ;
        RECT 131.100 71.955 131.630 72.295 ;
        RECT 129.010 70.625 129.630 71.025 ;
        RECT 127.360 69.375 127.890 69.715 ;
        RECT 125.320 68.055 125.940 68.455 ;
        RECT 123.720 66.795 124.250 67.135 ;
        RECT 121.650 65.475 122.270 65.875 ;
        RECT 106.975 63.125 108.900 63.495 ;
        RECT 109.245 62.765 119.830 63.715 ;
        RECT 121.690 63.295 122.150 65.475 ;
        RECT 123.810 64.555 124.190 66.795 ;
        RECT 125.370 65.865 125.830 68.055 ;
        RECT 127.460 67.135 127.840 69.375 ;
        RECT 129.050 68.445 129.510 70.625 ;
        RECT 131.200 69.715 131.580 71.955 ;
        RECT 132.740 71.035 133.200 73.205 ;
        RECT 134.840 72.295 135.220 74.535 ;
        RECT 136.410 73.615 136.870 75.795 ;
        RECT 138.550 74.885 138.930 77.105 ;
        RECT 140.090 76.195 140.550 77.495 ;
        RECT 142.190 77.445 142.570 78.380 ;
        RECT 142.100 77.105 142.630 77.445 ;
        RECT 140.050 75.795 140.670 76.195 ;
        RECT 138.440 74.545 138.970 74.885 ;
        RECT 136.350 73.215 136.970 73.615 ;
        RECT 134.740 71.955 135.270 72.295 ;
        RECT 132.690 70.635 133.310 71.035 ;
        RECT 131.100 69.375 131.630 69.715 ;
        RECT 129.000 68.045 129.620 68.445 ;
        RECT 127.360 66.795 127.890 67.135 ;
        RECT 125.300 65.465 125.920 65.865 ;
        RECT 123.720 64.215 124.250 64.555 ;
        RECT 121.630 62.895 122.250 63.295 ;
        RECT 108.540 61.585 108.890 61.605 ;
        RECT 108.520 61.225 108.960 61.585 ;
        RECT 108.540 56.995 108.890 61.225 ;
        RECT 109.220 59.295 109.570 61.605 ;
        RECT 109.150 58.935 109.570 59.295 ;
        RECT 108.520 56.635 108.960 56.995 ;
        RECT 108.540 52.435 108.890 56.635 ;
        RECT 109.220 54.725 109.570 58.935 ;
        RECT 109.150 54.365 109.570 54.725 ;
        RECT 108.520 52.075 108.960 52.435 ;
        RECT 108.540 47.855 108.890 52.075 ;
        RECT 109.220 50.135 109.570 54.365 ;
        RECT 110.855 53.350 111.905 53.380 ;
        RECT 110.855 52.300 117.810 53.350 ;
        RECT 110.855 52.270 111.905 52.300 ;
        RECT 109.150 49.775 109.570 50.135 ;
        RECT 108.520 47.495 108.960 47.855 ;
        RECT 108.540 43.265 108.890 47.495 ;
        RECT 109.220 45.555 109.570 49.775 ;
        RECT 118.880 50.015 119.830 62.765 ;
        RECT 121.690 60.695 122.150 62.895 ;
        RECT 123.810 61.975 124.190 64.215 ;
        RECT 125.370 63.285 125.830 65.465 ;
        RECT 127.460 64.555 127.840 66.795 ;
        RECT 129.050 65.885 129.510 68.045 ;
        RECT 131.200 67.135 131.580 69.375 ;
        RECT 132.740 68.445 133.200 70.635 ;
        RECT 134.840 69.715 135.220 71.955 ;
        RECT 136.410 71.025 136.870 73.215 ;
        RECT 138.550 72.295 138.930 74.545 ;
        RECT 140.090 73.605 140.550 75.795 ;
        RECT 142.190 74.875 142.570 77.105 ;
        RECT 143.770 76.205 144.230 77.495 ;
        RECT 145.880 77.445 146.260 78.380 ;
        RECT 145.780 77.105 146.310 77.445 ;
        RECT 143.730 75.805 144.350 76.205 ;
        RECT 142.100 74.535 142.630 74.875 ;
        RECT 140.030 73.205 140.650 73.605 ;
        RECT 138.440 71.955 138.970 72.295 ;
        RECT 136.360 70.625 136.980 71.025 ;
        RECT 134.740 69.375 135.270 69.715 ;
        RECT 132.690 68.045 133.310 68.445 ;
        RECT 131.100 66.795 131.630 67.135 ;
        RECT 129.000 65.485 129.620 65.885 ;
        RECT 127.360 64.215 127.890 64.555 ;
        RECT 125.320 62.885 125.940 63.285 ;
        RECT 123.720 61.635 124.250 61.975 ;
        RECT 121.640 60.295 122.260 60.695 ;
        RECT 121.690 58.135 122.150 60.295 ;
        RECT 123.810 59.395 124.190 61.635 ;
        RECT 125.370 60.705 125.830 62.885 ;
        RECT 127.460 61.975 127.840 64.215 ;
        RECT 129.050 63.285 129.510 65.485 ;
        RECT 131.200 64.545 131.580 66.795 ;
        RECT 132.740 65.885 133.200 68.045 ;
        RECT 134.840 67.135 135.220 69.375 ;
        RECT 136.410 68.445 136.870 70.625 ;
        RECT 138.550 69.715 138.930 71.955 ;
        RECT 140.090 71.025 140.550 73.205 ;
        RECT 142.190 72.295 142.570 74.535 ;
        RECT 143.770 73.605 144.230 75.805 ;
        RECT 145.880 74.875 146.260 77.105 ;
        RECT 145.780 74.535 146.310 74.875 ;
        RECT 143.730 73.205 144.350 73.605 ;
        RECT 142.100 71.955 142.630 72.295 ;
        RECT 140.040 70.625 140.660 71.025 ;
        RECT 138.440 69.375 138.970 69.715 ;
        RECT 136.350 68.045 136.970 68.445 ;
        RECT 134.740 66.795 135.270 67.135 ;
        RECT 132.690 65.485 133.310 65.885 ;
        RECT 131.100 64.205 131.630 64.545 ;
        RECT 129.000 62.885 129.620 63.285 ;
        RECT 127.360 61.635 127.890 61.975 ;
        RECT 125.340 60.305 125.960 60.705 ;
        RECT 123.720 59.055 124.250 59.395 ;
        RECT 121.640 57.735 122.260 58.135 ;
        RECT 121.690 55.545 122.150 57.735 ;
        RECT 123.810 56.815 124.190 59.055 ;
        RECT 125.370 58.135 125.830 60.305 ;
        RECT 127.460 59.395 127.840 61.635 ;
        RECT 129.050 60.705 129.510 62.885 ;
        RECT 131.200 61.985 131.580 64.205 ;
        RECT 132.740 63.285 133.200 65.485 ;
        RECT 134.840 64.555 135.220 66.795 ;
        RECT 136.410 65.865 136.870 68.045 ;
        RECT 138.550 67.135 138.930 69.375 ;
        RECT 140.090 68.445 140.550 70.625 ;
        RECT 142.190 69.705 142.570 71.955 ;
        RECT 143.770 71.015 144.230 73.205 ;
        RECT 145.880 72.295 146.260 74.535 ;
        RECT 145.780 71.955 146.310 72.295 ;
        RECT 143.730 70.615 144.350 71.015 ;
        RECT 142.100 69.365 142.630 69.705 ;
        RECT 140.030 68.045 140.650 68.445 ;
        RECT 138.440 66.795 138.970 67.135 ;
        RECT 136.350 65.465 136.970 65.865 ;
        RECT 134.740 64.215 135.270 64.555 ;
        RECT 132.680 62.885 133.300 63.285 ;
        RECT 131.100 61.645 131.630 61.985 ;
        RECT 129.010 60.305 129.630 60.705 ;
        RECT 127.360 59.055 127.890 59.395 ;
        RECT 125.320 57.735 125.940 58.135 ;
        RECT 123.720 56.475 124.250 56.815 ;
        RECT 121.650 55.145 122.270 55.545 ;
        RECT 121.690 52.965 122.150 55.145 ;
        RECT 123.810 54.235 124.190 56.475 ;
        RECT 125.370 55.555 125.830 57.735 ;
        RECT 127.460 56.815 127.840 59.055 ;
        RECT 129.050 58.145 129.510 60.305 ;
        RECT 131.200 59.395 131.580 61.645 ;
        RECT 132.740 60.705 133.200 62.885 ;
        RECT 134.840 61.975 135.220 64.215 ;
        RECT 136.410 63.275 136.870 65.465 ;
        RECT 138.550 64.555 138.930 66.795 ;
        RECT 140.090 65.855 140.550 68.045 ;
        RECT 142.190 67.145 142.570 69.365 ;
        RECT 143.770 68.435 144.230 70.615 ;
        RECT 145.880 69.715 146.260 71.955 ;
        RECT 145.780 69.375 146.310 69.715 ;
        RECT 143.710 68.035 144.330 68.435 ;
        RECT 142.100 66.805 142.630 67.145 ;
        RECT 140.060 65.455 140.680 65.855 ;
        RECT 138.440 64.215 138.970 64.555 ;
        RECT 136.360 62.875 136.980 63.275 ;
        RECT 134.740 61.635 135.270 61.975 ;
        RECT 132.690 60.305 133.310 60.705 ;
        RECT 131.100 59.055 131.630 59.395 ;
        RECT 128.990 57.745 129.610 58.145 ;
        RECT 127.360 56.475 127.890 56.815 ;
        RECT 125.330 55.155 125.950 55.555 ;
        RECT 123.720 53.895 124.250 54.235 ;
        RECT 121.650 52.565 122.270 52.965 ;
        RECT 121.690 50.015 122.150 52.565 ;
        RECT 123.810 51.655 124.190 53.895 ;
        RECT 125.370 52.975 125.830 55.155 ;
        RECT 127.460 54.235 127.840 56.475 ;
        RECT 129.050 55.545 129.510 57.745 ;
        RECT 131.200 56.825 131.580 59.055 ;
        RECT 132.740 58.115 133.200 60.305 ;
        RECT 134.840 59.395 135.220 61.635 ;
        RECT 136.410 60.705 136.870 62.875 ;
        RECT 138.550 61.975 138.930 64.215 ;
        RECT 140.090 63.285 140.550 65.455 ;
        RECT 142.190 64.555 142.570 66.805 ;
        RECT 143.770 65.865 144.230 68.035 ;
        RECT 145.880 67.125 146.260 69.375 ;
        RECT 145.780 66.785 146.310 67.125 ;
        RECT 143.730 65.465 144.350 65.865 ;
        RECT 142.080 64.215 142.610 64.555 ;
        RECT 140.040 62.885 140.660 63.285 ;
        RECT 138.440 61.635 138.970 61.975 ;
        RECT 136.370 60.305 136.990 60.705 ;
        RECT 134.740 59.055 135.270 59.395 ;
        RECT 132.690 57.715 133.310 58.115 ;
        RECT 131.100 56.485 131.630 56.825 ;
        RECT 129.000 55.145 129.620 55.545 ;
        RECT 127.360 53.895 127.890 54.235 ;
        RECT 125.320 52.575 125.940 52.975 ;
        RECT 123.720 51.315 124.250 51.655 ;
        RECT 123.810 51.235 124.190 51.315 ;
        RECT 125.370 50.015 125.830 52.575 ;
        RECT 127.460 51.655 127.840 53.895 ;
        RECT 129.050 52.985 129.510 55.145 ;
        RECT 131.200 54.235 131.580 56.485 ;
        RECT 132.740 55.545 133.200 57.715 ;
        RECT 134.840 56.815 135.220 59.055 ;
        RECT 136.410 58.135 136.870 60.305 ;
        RECT 138.550 59.395 138.930 61.635 ;
        RECT 140.090 60.705 140.550 62.885 ;
        RECT 142.190 61.975 142.570 64.215 ;
        RECT 143.770 63.285 144.230 65.465 ;
        RECT 145.880 64.555 146.260 66.785 ;
        RECT 145.780 64.215 146.310 64.555 ;
        RECT 143.740 62.885 144.360 63.285 ;
        RECT 142.080 61.635 142.610 61.975 ;
        RECT 140.030 60.305 140.650 60.705 ;
        RECT 138.440 59.055 138.970 59.395 ;
        RECT 136.370 57.735 136.990 58.135 ;
        RECT 134.740 56.475 135.270 56.815 ;
        RECT 132.690 55.145 133.310 55.545 ;
        RECT 131.100 53.895 131.630 54.235 ;
        RECT 129.000 52.585 129.620 52.985 ;
        RECT 127.360 51.315 127.890 51.655 ;
        RECT 127.460 51.235 127.840 51.315 ;
        RECT 129.050 50.015 129.510 52.585 ;
        RECT 131.200 51.655 131.580 53.895 ;
        RECT 132.740 52.975 133.200 55.145 ;
        RECT 134.840 54.235 135.220 56.475 ;
        RECT 136.410 55.555 136.870 57.735 ;
        RECT 138.550 56.815 138.930 59.055 ;
        RECT 140.090 58.125 140.550 60.305 ;
        RECT 142.190 59.405 142.570 61.635 ;
        RECT 143.770 60.715 144.230 62.885 ;
        RECT 145.880 61.965 146.260 64.215 ;
        RECT 145.780 61.625 146.310 61.965 ;
        RECT 143.740 60.315 144.360 60.715 ;
        RECT 142.080 59.065 142.610 59.405 ;
        RECT 140.050 57.725 140.670 58.125 ;
        RECT 138.440 56.475 138.970 56.815 ;
        RECT 136.360 55.155 136.980 55.555 ;
        RECT 134.740 53.895 135.270 54.235 ;
        RECT 132.690 52.575 133.310 52.975 ;
        RECT 131.100 51.315 131.630 51.655 ;
        RECT 131.200 51.235 131.580 51.315 ;
        RECT 132.740 50.015 133.200 52.575 ;
        RECT 134.840 51.645 135.220 53.895 ;
        RECT 136.410 52.965 136.870 55.155 ;
        RECT 138.550 54.235 138.930 56.475 ;
        RECT 140.090 55.555 140.550 57.725 ;
        RECT 142.190 56.815 142.570 59.065 ;
        RECT 143.770 58.115 144.230 60.315 ;
        RECT 145.880 59.395 146.260 61.625 ;
        RECT 145.780 59.055 146.310 59.395 ;
        RECT 143.730 57.715 144.350 58.115 ;
        RECT 142.080 56.475 142.610 56.815 ;
        RECT 140.050 55.155 140.670 55.555 ;
        RECT 138.440 53.895 138.970 54.235 ;
        RECT 136.370 52.565 136.990 52.965 ;
        RECT 134.740 51.305 135.270 51.645 ;
        RECT 134.840 51.235 135.220 51.305 ;
        RECT 136.410 50.015 136.870 52.565 ;
        RECT 138.550 51.655 138.930 53.895 ;
        RECT 140.090 52.965 140.550 55.155 ;
        RECT 142.190 54.225 142.570 56.475 ;
        RECT 143.770 55.535 144.230 57.715 ;
        RECT 145.880 56.805 146.260 59.055 ;
        RECT 145.780 56.465 146.310 56.805 ;
        RECT 143.720 55.135 144.340 55.535 ;
        RECT 142.080 53.885 142.610 54.225 ;
        RECT 140.050 52.565 140.670 52.965 ;
        RECT 138.440 51.315 138.970 51.655 ;
        RECT 138.550 51.235 138.930 51.315 ;
        RECT 140.090 50.015 140.550 52.565 ;
        RECT 142.190 51.645 142.570 53.885 ;
        RECT 143.770 52.965 144.230 55.135 ;
        RECT 145.880 54.235 146.260 56.465 ;
        RECT 145.780 53.895 146.310 54.235 ;
        RECT 143.730 52.565 144.350 52.965 ;
        RECT 142.080 51.305 142.610 51.645 ;
        RECT 142.190 51.235 142.570 51.305 ;
        RECT 143.770 50.015 144.230 52.565 ;
        RECT 145.880 51.645 146.260 53.895 ;
        RECT 145.780 51.305 146.310 51.645 ;
        RECT 145.880 51.245 146.260 51.305 ;
        RECT 118.880 49.555 144.230 50.015 ;
        RECT 131.150 48.680 131.880 49.555 ;
        RECT 131.120 47.950 131.910 48.680 ;
        RECT 109.150 45.195 109.570 45.555 ;
        RECT 108.520 42.905 108.960 43.265 ;
        RECT 108.540 38.685 108.890 42.905 ;
        RECT 109.220 40.975 109.570 45.195 ;
        RECT 116.550 46.625 141.995 47.280 ;
        RECT 113.670 43.525 114.100 43.885 ;
        RECT 109.150 40.615 109.570 40.975 ;
        RECT 108.520 38.325 108.960 38.685 ;
        RECT 108.540 36.730 108.890 38.325 ;
        RECT 107.515 36.380 108.890 36.730 ;
        RECT 108.540 36.355 108.890 36.380 ;
        RECT 109.220 36.695 109.570 40.615 ;
        RECT 113.720 39.295 114.040 43.525 ;
        RECT 114.300 41.595 114.620 43.875 ;
        RECT 114.230 41.245 114.660 41.595 ;
        RECT 113.670 38.935 114.100 39.295 ;
        RECT 113.720 38.045 114.040 38.935 ;
        RECT 114.300 38.065 114.620 41.245 ;
        RECT 112.870 37.725 114.040 38.045 ;
        RECT 114.270 37.745 114.650 38.065 ;
        RECT 114.300 37.725 114.620 37.745 ;
        RECT 116.550 36.855 117.205 46.625 ;
        RECT 118.770 45.145 124.300 45.575 ;
        RECT 127.805 45.265 136.545 45.820 ;
        RECT 118.770 44.045 119.200 45.145 ;
        RECT 118.720 43.725 119.240 44.045 ;
        RECT 118.770 43.085 119.200 43.725 ;
        RECT 122.240 43.555 122.670 44.115 ;
        RECT 123.870 44.035 124.300 45.145 ;
        RECT 123.810 43.715 124.330 44.035 ;
        RECT 122.170 43.235 122.690 43.555 ;
        RECT 118.720 42.765 119.240 43.085 ;
        RECT 118.770 42.125 119.200 42.765 ;
        RECT 122.240 42.605 122.670 43.235 ;
        RECT 123.870 43.085 124.300 43.715 ;
        RECT 127.330 43.565 127.760 44.115 ;
        RECT 131.590 43.685 132.110 43.955 ;
        RECT 127.260 43.245 127.780 43.565 ;
        RECT 123.810 42.765 124.330 43.085 ;
        RECT 122.170 42.285 122.690 42.605 ;
        RECT 118.720 41.805 119.240 42.125 ;
        RECT 118.770 41.155 119.200 41.805 ;
        RECT 122.240 41.645 122.670 42.285 ;
        RECT 123.870 42.115 124.300 42.765 ;
        RECT 127.330 42.605 127.760 43.245 ;
        RECT 131.590 42.995 132.020 43.685 ;
        RECT 135.990 43.475 136.545 45.265 ;
        RECT 135.990 43.195 136.550 43.475 ;
        RECT 131.590 42.725 132.110 42.995 ;
        RECT 127.260 42.285 127.780 42.605 ;
        RECT 123.810 41.795 124.330 42.115 ;
        RECT 122.170 41.325 122.690 41.645 ;
        RECT 118.720 40.835 119.240 41.155 ;
        RECT 118.770 40.205 119.200 40.835 ;
        RECT 122.240 40.685 122.670 41.325 ;
        RECT 123.870 41.165 124.300 41.795 ;
        RECT 127.330 41.645 127.760 42.285 ;
        RECT 131.590 42.035 132.020 42.725 ;
        RECT 135.990 42.525 136.545 43.195 ;
        RECT 144.160 43.105 145.280 43.135 ;
        RECT 135.990 42.245 136.550 42.525 ;
        RECT 131.590 41.765 132.110 42.035 ;
        RECT 127.260 41.325 127.780 41.645 ;
        RECT 123.810 40.845 124.330 41.165 ;
        RECT 122.170 40.365 122.690 40.685 ;
        RECT 118.720 39.885 119.240 40.205 ;
        RECT 118.770 39.255 119.200 39.885 ;
        RECT 122.240 39.725 122.670 40.365 ;
        RECT 123.870 40.205 124.300 40.845 ;
        RECT 127.330 40.685 127.760 41.325 ;
        RECT 131.590 41.075 132.020 41.765 ;
        RECT 135.990 41.565 136.545 42.245 ;
        RECT 144.160 41.985 148.130 43.105 ;
        RECT 144.160 41.955 145.280 41.985 ;
        RECT 135.990 41.285 136.550 41.565 ;
        RECT 131.590 40.805 132.110 41.075 ;
        RECT 127.260 40.365 127.780 40.685 ;
        RECT 123.810 39.885 124.330 40.205 ;
        RECT 122.170 39.405 122.690 39.725 ;
        RECT 118.720 38.935 119.240 39.255 ;
        RECT 118.770 37.490 119.200 38.935 ;
        RECT 122.240 37.710 122.670 39.405 ;
        RECT 123.870 39.245 124.300 39.885 ;
        RECT 127.330 39.725 127.760 40.365 ;
        RECT 131.590 40.115 132.020 40.805 ;
        RECT 135.990 40.605 136.545 41.285 ;
        RECT 135.990 40.325 136.550 40.605 ;
        RECT 131.590 39.845 132.110 40.115 ;
        RECT 127.260 39.405 127.780 39.725 ;
        RECT 123.810 38.925 124.330 39.245 ;
        RECT 127.330 38.230 127.760 39.405 ;
        RECT 127.325 38.025 127.760 38.230 ;
        RECT 131.590 39.155 132.020 39.845 ;
        RECT 135.990 39.645 136.545 40.325 ;
        RECT 135.990 39.365 136.550 39.645 ;
        RECT 131.590 38.885 132.110 39.155 ;
        RECT 127.325 37.710 127.755 38.025 ;
        RECT 122.240 37.280 127.800 37.710 ;
        RECT 131.590 37.655 132.020 38.885 ;
        RECT 135.990 37.985 136.545 39.365 ;
        RECT 131.450 37.400 132.140 37.655 ;
        RECT 135.990 37.425 144.290 37.985 ;
        RECT 135.990 37.420 136.545 37.425 ;
        RECT 110.670 36.695 117.205 36.855 ;
        RECT 131.455 36.715 132.140 37.400 ;
        RECT 109.220 36.360 117.205 36.695 ;
        RECT 109.220 36.355 109.570 36.360 ;
        RECT 110.670 36.200 117.205 36.360 ;
        RECT 119.690 36.030 132.140 36.715 ;
        RECT 119.690 34.610 120.375 36.030 ;
        RECT 138.240 35.625 139.060 36.385 ;
        RECT 136.190 35.355 136.825 35.375 ;
        RECT 138.270 35.355 139.030 35.625 ;
        RECT 136.165 34.670 150.060 35.355 ;
        RECT 136.190 34.650 136.825 34.670 ;
        RECT 114.680 33.925 120.375 34.610 ;
        RECT 123.360 30.935 124.165 32.570 ;
        RECT 129.210 30.985 129.955 32.100 ;
        RECT 123.340 30.180 124.185 30.935 ;
        RECT 129.190 30.290 129.975 30.985 ;
        RECT 129.210 30.265 129.955 30.290 ;
        RECT 123.360 30.155 124.165 30.180 ;
      LAYER via2 ;
        RECT 149.375 167.185 150.825 168.635 ;
        RECT 103.175 163.595 104.625 165.045 ;
        RECT 118.190 149.070 119.030 149.910 ;
        RECT 138.755 149.050 139.560 149.855 ;
        RECT 126.370 129.255 126.650 129.535 ;
        RECT 128.425 127.500 128.725 127.800 ;
        RECT 130.515 127.500 130.815 127.800 ;
        RECT 132.615 127.500 132.915 127.800 ;
        RECT 134.705 127.500 135.005 127.800 ;
        RECT 128.430 112.185 128.730 112.485 ;
        RECT 130.530 112.185 130.830 112.485 ;
        RECT 132.590 112.185 132.890 112.485 ;
        RECT 134.680 112.185 134.980 112.485 ;
        RECT 126.340 110.360 126.625 110.645 ;
        RECT 120.425 109.180 121.175 109.930 ;
        RECT 126.490 109.155 127.290 109.955 ;
        RECT 127.325 37.280 127.755 37.710 ;
        RECT 136.190 34.695 136.825 35.330 ;
        RECT 123.385 30.180 124.140 30.935 ;
        RECT 129.235 30.290 129.930 30.985 ;
      LAYER met3 ;
        RECT 32.975 177.310 34.465 177.335 ;
        RECT 32.970 175.810 150.850 177.310 ;
        RECT 32.975 175.785 34.465 175.810 ;
        RECT 103.150 168.685 104.650 168.690 ;
        RECT 103.125 167.195 104.675 168.685 ;
        RECT 103.150 163.570 104.650 167.195 ;
        RECT 149.350 167.160 150.850 175.810 ;
        RECT 138.730 151.205 139.585 151.210 ;
        RECT 118.165 151.170 119.055 151.175 ;
        RECT 118.140 150.290 119.080 151.170 ;
        RECT 138.705 150.360 139.610 151.205 ;
        RECT 118.165 149.045 119.055 150.290 ;
        RECT 138.730 149.025 139.585 150.360 ;
        RECT 126.345 129.545 126.675 129.560 ;
        RECT 126.345 129.245 135.005 129.545 ;
        RECT 126.345 129.230 126.675 129.245 ;
        RECT 128.425 127.825 128.725 129.245 ;
        RECT 130.515 127.825 130.815 129.245 ;
        RECT 132.615 127.825 132.915 129.245 ;
        RECT 134.705 127.825 135.005 129.245 ;
        RECT 128.400 127.475 128.750 127.825 ;
        RECT 130.490 127.475 130.840 127.825 ;
        RECT 132.590 127.475 132.940 127.825 ;
        RECT 134.680 127.475 135.030 127.825 ;
        RECT 128.405 112.160 128.755 112.510 ;
        RECT 130.505 112.160 130.855 112.510 ;
        RECT 132.565 112.160 132.915 112.510 ;
        RECT 134.655 112.160 135.005 112.510 ;
        RECT 128.430 110.670 128.730 112.160 ;
        RECT 130.530 110.670 130.830 112.160 ;
        RECT 132.590 110.670 132.890 112.160 ;
        RECT 134.680 110.670 134.980 112.160 ;
        RECT 126.315 110.335 135.000 110.670 ;
        RECT 126.465 109.955 127.315 109.980 ;
        RECT 120.400 109.155 127.315 109.955 ;
        RECT 126.465 109.130 127.315 109.155 ;
        RECT 127.300 37.710 127.780 37.735 ;
        RECT 127.300 37.280 132.885 37.710 ;
        RECT 127.300 37.255 127.780 37.280 ;
        RECT 132.455 35.230 132.885 37.280 ;
        RECT 135.600 35.230 136.850 35.355 ;
        RECT 132.455 34.800 136.850 35.230 ;
        RECT 135.600 34.670 136.850 34.800 ;
        RECT 123.360 28.355 124.165 30.960 ;
        RECT 129.210 29.290 129.955 31.010 ;
        RECT 129.185 28.555 129.980 29.290 ;
        RECT 129.210 28.550 129.955 28.555 ;
        RECT 123.365 28.330 124.160 28.355 ;
      LAYER via3 ;
        RECT 32.975 175.815 34.465 177.305 ;
        RECT 103.155 167.195 104.645 168.685 ;
        RECT 118.170 150.290 119.050 151.170 ;
        RECT 138.735 150.360 139.580 151.205 ;
        RECT 123.365 28.360 124.160 29.155 ;
        RECT 129.215 28.555 129.950 29.290 ;
      LAYER met4 ;
        RECT 3.990 223.750 4.290 224.760 ;
        RECT 7.670 223.750 7.970 224.760 ;
        RECT 11.350 223.750 11.650 224.760 ;
        RECT 15.030 223.750 15.330 224.760 ;
        RECT 18.710 223.750 19.010 224.760 ;
        RECT 22.390 223.750 22.690 224.760 ;
        RECT 26.070 223.750 26.370 224.760 ;
        RECT 29.750 223.750 30.050 224.760 ;
        RECT 33.430 223.750 33.730 224.760 ;
        RECT 37.110 223.750 37.410 224.760 ;
        RECT 40.790 223.750 41.090 224.760 ;
        RECT 44.470 223.750 44.770 224.760 ;
        RECT 48.150 223.750 48.450 224.760 ;
        RECT 51.830 223.750 52.130 224.760 ;
        RECT 55.510 223.750 55.810 224.760 ;
        RECT 59.190 223.750 59.490 224.760 ;
        RECT 62.870 223.750 63.170 224.760 ;
        RECT 66.550 223.750 66.850 224.760 ;
        RECT 70.230 223.750 70.530 224.760 ;
        RECT 73.910 223.750 74.210 224.760 ;
        RECT 77.590 223.750 77.890 224.760 ;
        RECT 81.270 223.750 81.570 224.760 ;
        RECT 84.950 223.750 85.250 224.760 ;
        RECT 88.630 223.750 88.930 224.760 ;
        RECT 3.810 222.090 88.930 223.750 ;
        RECT 49.000 220.760 50.500 222.090 ;
        RECT 88.630 222.080 88.930 222.090 ;
        RECT 2.500 175.810 34.470 177.310 ;
        RECT 50.500 167.190 104.650 168.690 ;
        RECT 83.090 156.465 139.585 157.320 ;
        RECT 83.090 21.190 83.945 156.465 ;
        RECT 90.175 151.775 119.055 152.665 ;
        RECT 90.320 25.625 90.920 151.775 ;
        RECT 118.165 150.285 119.055 151.775 ;
        RECT 138.730 150.355 139.585 156.465 ;
        RECT 90.320 25.015 113.005 25.625 ;
        RECT 90.320 25.000 90.920 25.015 ;
        RECT 83.090 20.590 90.920 21.190 ;
        RECT 68.240 1.000 68.840 1.010 ;
        RECT 90.320 1.000 90.920 20.590 ;
        RECT 112.395 1.000 113.005 25.015 ;
        RECT 123.360 24.215 124.165 29.160 ;
        RECT 129.210 28.550 157.235 29.295 ;
        RECT 123.360 23.410 135.185 24.215 ;
        RECT 134.480 1.000 135.080 23.410 ;
        RECT 156.560 1.000 157.160 28.550 ;
        RECT 112.395 0.235 112.400 1.000 ;
        RECT 113.000 0.235 113.005 1.000 ;
  END
END tt_um_alfiero88_VCII
END LIBRARY

