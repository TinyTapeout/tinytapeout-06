module tt_um_MichaelBell_latch_mem (VGND,
    VPWR,
    clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input VGND;
 input VPWR;
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire \RAM[0][0] ;
 wire \RAM[0][1] ;
 wire \RAM[0][2] ;
 wire \RAM[0][3] ;
 wire \RAM[0][4] ;
 wire \RAM[0][5] ;
 wire \RAM[0][6] ;
 wire \RAM[0][7] ;
 wire \RAM[10][0] ;
 wire \RAM[10][1] ;
 wire \RAM[10][2] ;
 wire \RAM[10][3] ;
 wire \RAM[10][4] ;
 wire \RAM[10][5] ;
 wire \RAM[10][6] ;
 wire \RAM[10][7] ;
 wire \RAM[11][0] ;
 wire \RAM[11][1] ;
 wire \RAM[11][2] ;
 wire \RAM[11][3] ;
 wire \RAM[11][4] ;
 wire \RAM[11][5] ;
 wire \RAM[11][6] ;
 wire \RAM[11][7] ;
 wire \RAM[12][0] ;
 wire \RAM[12][1] ;
 wire \RAM[12][2] ;
 wire \RAM[12][3] ;
 wire \RAM[12][4] ;
 wire \RAM[12][5] ;
 wire \RAM[12][6] ;
 wire \RAM[12][7] ;
 wire \RAM[13][0] ;
 wire \RAM[13][1] ;
 wire \RAM[13][2] ;
 wire \RAM[13][3] ;
 wire \RAM[13][4] ;
 wire \RAM[13][5] ;
 wire \RAM[13][6] ;
 wire \RAM[13][7] ;
 wire \RAM[14][0] ;
 wire \RAM[14][1] ;
 wire \RAM[14][2] ;
 wire \RAM[14][3] ;
 wire \RAM[14][4] ;
 wire \RAM[14][5] ;
 wire \RAM[14][6] ;
 wire \RAM[14][7] ;
 wire \RAM[15][0] ;
 wire \RAM[15][1] ;
 wire \RAM[15][2] ;
 wire \RAM[15][3] ;
 wire \RAM[15][4] ;
 wire \RAM[15][5] ;
 wire \RAM[15][6] ;
 wire \RAM[15][7] ;
 wire \RAM[16][0] ;
 wire \RAM[16][1] ;
 wire \RAM[16][2] ;
 wire \RAM[16][3] ;
 wire \RAM[16][4] ;
 wire \RAM[16][5] ;
 wire \RAM[16][6] ;
 wire \RAM[16][7] ;
 wire \RAM[17][0] ;
 wire \RAM[17][1] ;
 wire \RAM[17][2] ;
 wire \RAM[17][3] ;
 wire \RAM[17][4] ;
 wire \RAM[17][5] ;
 wire \RAM[17][6] ;
 wire \RAM[17][7] ;
 wire \RAM[18][0] ;
 wire \RAM[18][1] ;
 wire \RAM[18][2] ;
 wire \RAM[18][3] ;
 wire \RAM[18][4] ;
 wire \RAM[18][5] ;
 wire \RAM[18][6] ;
 wire \RAM[18][7] ;
 wire \RAM[19][0] ;
 wire \RAM[19][1] ;
 wire \RAM[19][2] ;
 wire \RAM[19][3] ;
 wire \RAM[19][4] ;
 wire \RAM[19][5] ;
 wire \RAM[19][6] ;
 wire \RAM[19][7] ;
 wire \RAM[1][0] ;
 wire \RAM[1][1] ;
 wire \RAM[1][2] ;
 wire \RAM[1][3] ;
 wire \RAM[1][4] ;
 wire \RAM[1][5] ;
 wire \RAM[1][6] ;
 wire \RAM[1][7] ;
 wire \RAM[20][0] ;
 wire \RAM[20][1] ;
 wire \RAM[20][2] ;
 wire \RAM[20][3] ;
 wire \RAM[20][4] ;
 wire \RAM[20][5] ;
 wire \RAM[20][6] ;
 wire \RAM[20][7] ;
 wire \RAM[21][0] ;
 wire \RAM[21][1] ;
 wire \RAM[21][2] ;
 wire \RAM[21][3] ;
 wire \RAM[21][4] ;
 wire \RAM[21][5] ;
 wire \RAM[21][6] ;
 wire \RAM[21][7] ;
 wire \RAM[22][0] ;
 wire \RAM[22][1] ;
 wire \RAM[22][2] ;
 wire \RAM[22][3] ;
 wire \RAM[22][4] ;
 wire \RAM[22][5] ;
 wire \RAM[22][6] ;
 wire \RAM[22][7] ;
 wire \RAM[23][0] ;
 wire \RAM[23][1] ;
 wire \RAM[23][2] ;
 wire \RAM[23][3] ;
 wire \RAM[23][4] ;
 wire \RAM[23][5] ;
 wire \RAM[23][6] ;
 wire \RAM[23][7] ;
 wire \RAM[24][0] ;
 wire \RAM[24][1] ;
 wire \RAM[24][2] ;
 wire \RAM[24][3] ;
 wire \RAM[24][4] ;
 wire \RAM[24][5] ;
 wire \RAM[24][6] ;
 wire \RAM[24][7] ;
 wire \RAM[25][0] ;
 wire \RAM[25][1] ;
 wire \RAM[25][2] ;
 wire \RAM[25][3] ;
 wire \RAM[25][4] ;
 wire \RAM[25][5] ;
 wire \RAM[25][6] ;
 wire \RAM[25][7] ;
 wire \RAM[26][0] ;
 wire \RAM[26][1] ;
 wire \RAM[26][2] ;
 wire \RAM[26][3] ;
 wire \RAM[26][4] ;
 wire \RAM[26][5] ;
 wire \RAM[26][6] ;
 wire \RAM[26][7] ;
 wire \RAM[27][0] ;
 wire \RAM[27][1] ;
 wire \RAM[27][2] ;
 wire \RAM[27][3] ;
 wire \RAM[27][4] ;
 wire \RAM[27][5] ;
 wire \RAM[27][6] ;
 wire \RAM[27][7] ;
 wire \RAM[28][0] ;
 wire \RAM[28][1] ;
 wire \RAM[28][2] ;
 wire \RAM[28][3] ;
 wire \RAM[28][4] ;
 wire \RAM[28][5] ;
 wire \RAM[28][6] ;
 wire \RAM[28][7] ;
 wire \RAM[29][0] ;
 wire \RAM[29][1] ;
 wire \RAM[29][2] ;
 wire \RAM[29][3] ;
 wire \RAM[29][4] ;
 wire \RAM[29][5] ;
 wire \RAM[29][6] ;
 wire \RAM[29][7] ;
 wire \RAM[2][0] ;
 wire \RAM[2][1] ;
 wire \RAM[2][2] ;
 wire \RAM[2][3] ;
 wire \RAM[2][4] ;
 wire \RAM[2][5] ;
 wire \RAM[2][6] ;
 wire \RAM[2][7] ;
 wire \RAM[30][0] ;
 wire \RAM[30][1] ;
 wire \RAM[30][2] ;
 wire \RAM[30][3] ;
 wire \RAM[30][4] ;
 wire \RAM[30][5] ;
 wire \RAM[30][6] ;
 wire \RAM[30][7] ;
 wire \RAM[31][0] ;
 wire \RAM[31][1] ;
 wire \RAM[31][2] ;
 wire \RAM[31][3] ;
 wire \RAM[31][4] ;
 wire \RAM[31][5] ;
 wire \RAM[31][6] ;
 wire \RAM[31][7] ;
 wire \RAM[32][0] ;
 wire \RAM[32][1] ;
 wire \RAM[32][2] ;
 wire \RAM[32][3] ;
 wire \RAM[32][4] ;
 wire \RAM[32][5] ;
 wire \RAM[32][6] ;
 wire \RAM[32][7] ;
 wire \RAM[33][0] ;
 wire \RAM[33][1] ;
 wire \RAM[33][2] ;
 wire \RAM[33][3] ;
 wire \RAM[33][4] ;
 wire \RAM[33][5] ;
 wire \RAM[33][6] ;
 wire \RAM[33][7] ;
 wire \RAM[34][0] ;
 wire \RAM[34][1] ;
 wire \RAM[34][2] ;
 wire \RAM[34][3] ;
 wire \RAM[34][4] ;
 wire \RAM[34][5] ;
 wire \RAM[34][6] ;
 wire \RAM[34][7] ;
 wire \RAM[35][0] ;
 wire \RAM[35][1] ;
 wire \RAM[35][2] ;
 wire \RAM[35][3] ;
 wire \RAM[35][4] ;
 wire \RAM[35][5] ;
 wire \RAM[35][6] ;
 wire \RAM[35][7] ;
 wire \RAM[36][0] ;
 wire \RAM[36][1] ;
 wire \RAM[36][2] ;
 wire \RAM[36][3] ;
 wire \RAM[36][4] ;
 wire \RAM[36][5] ;
 wire \RAM[36][6] ;
 wire \RAM[36][7] ;
 wire \RAM[37][0] ;
 wire \RAM[37][1] ;
 wire \RAM[37][2] ;
 wire \RAM[37][3] ;
 wire \RAM[37][4] ;
 wire \RAM[37][5] ;
 wire \RAM[37][6] ;
 wire \RAM[37][7] ;
 wire \RAM[38][0] ;
 wire \RAM[38][1] ;
 wire \RAM[38][2] ;
 wire \RAM[38][3] ;
 wire \RAM[38][4] ;
 wire \RAM[38][5] ;
 wire \RAM[38][6] ;
 wire \RAM[38][7] ;
 wire \RAM[39][0] ;
 wire \RAM[39][1] ;
 wire \RAM[39][2] ;
 wire \RAM[39][3] ;
 wire \RAM[39][4] ;
 wire \RAM[39][5] ;
 wire \RAM[39][6] ;
 wire \RAM[39][7] ;
 wire \RAM[3][0] ;
 wire \RAM[3][1] ;
 wire \RAM[3][2] ;
 wire \RAM[3][3] ;
 wire \RAM[3][4] ;
 wire \RAM[3][5] ;
 wire \RAM[3][6] ;
 wire \RAM[3][7] ;
 wire \RAM[40][0] ;
 wire \RAM[40][1] ;
 wire \RAM[40][2] ;
 wire \RAM[40][3] ;
 wire \RAM[40][4] ;
 wire \RAM[40][5] ;
 wire \RAM[40][6] ;
 wire \RAM[40][7] ;
 wire \RAM[41][0] ;
 wire \RAM[41][1] ;
 wire \RAM[41][2] ;
 wire \RAM[41][3] ;
 wire \RAM[41][4] ;
 wire \RAM[41][5] ;
 wire \RAM[41][6] ;
 wire \RAM[41][7] ;
 wire \RAM[42][0] ;
 wire \RAM[42][1] ;
 wire \RAM[42][2] ;
 wire \RAM[42][3] ;
 wire \RAM[42][4] ;
 wire \RAM[42][5] ;
 wire \RAM[42][6] ;
 wire \RAM[42][7] ;
 wire \RAM[43][0] ;
 wire \RAM[43][1] ;
 wire \RAM[43][2] ;
 wire \RAM[43][3] ;
 wire \RAM[43][4] ;
 wire \RAM[43][5] ;
 wire \RAM[43][6] ;
 wire \RAM[43][7] ;
 wire \RAM[44][0] ;
 wire \RAM[44][1] ;
 wire \RAM[44][2] ;
 wire \RAM[44][3] ;
 wire \RAM[44][4] ;
 wire \RAM[44][5] ;
 wire \RAM[44][6] ;
 wire \RAM[44][7] ;
 wire \RAM[45][0] ;
 wire \RAM[45][1] ;
 wire \RAM[45][2] ;
 wire \RAM[45][3] ;
 wire \RAM[45][4] ;
 wire \RAM[45][5] ;
 wire \RAM[45][6] ;
 wire \RAM[45][7] ;
 wire \RAM[46][0] ;
 wire \RAM[46][1] ;
 wire \RAM[46][2] ;
 wire \RAM[46][3] ;
 wire \RAM[46][4] ;
 wire \RAM[46][5] ;
 wire \RAM[46][6] ;
 wire \RAM[46][7] ;
 wire \RAM[47][0] ;
 wire \RAM[47][1] ;
 wire \RAM[47][2] ;
 wire \RAM[47][3] ;
 wire \RAM[47][4] ;
 wire \RAM[47][5] ;
 wire \RAM[47][6] ;
 wire \RAM[47][7] ;
 wire \RAM[48][0] ;
 wire \RAM[48][1] ;
 wire \RAM[48][2] ;
 wire \RAM[48][3] ;
 wire \RAM[48][4] ;
 wire \RAM[48][5] ;
 wire \RAM[48][6] ;
 wire \RAM[48][7] ;
 wire \RAM[49][0] ;
 wire \RAM[49][1] ;
 wire \RAM[49][2] ;
 wire \RAM[49][3] ;
 wire \RAM[49][4] ;
 wire \RAM[49][5] ;
 wire \RAM[49][6] ;
 wire \RAM[49][7] ;
 wire \RAM[4][0] ;
 wire \RAM[4][1] ;
 wire \RAM[4][2] ;
 wire \RAM[4][3] ;
 wire \RAM[4][4] ;
 wire \RAM[4][5] ;
 wire \RAM[4][6] ;
 wire \RAM[4][7] ;
 wire \RAM[50][0] ;
 wire \RAM[50][1] ;
 wire \RAM[50][2] ;
 wire \RAM[50][3] ;
 wire \RAM[50][4] ;
 wire \RAM[50][5] ;
 wire \RAM[50][6] ;
 wire \RAM[50][7] ;
 wire \RAM[51][0] ;
 wire \RAM[51][1] ;
 wire \RAM[51][2] ;
 wire \RAM[51][3] ;
 wire \RAM[51][4] ;
 wire \RAM[51][5] ;
 wire \RAM[51][6] ;
 wire \RAM[51][7] ;
 wire \RAM[52][0] ;
 wire \RAM[52][1] ;
 wire \RAM[52][2] ;
 wire \RAM[52][3] ;
 wire \RAM[52][4] ;
 wire \RAM[52][5] ;
 wire \RAM[52][6] ;
 wire \RAM[52][7] ;
 wire \RAM[53][0] ;
 wire \RAM[53][1] ;
 wire \RAM[53][2] ;
 wire \RAM[53][3] ;
 wire \RAM[53][4] ;
 wire \RAM[53][5] ;
 wire \RAM[53][6] ;
 wire \RAM[53][7] ;
 wire \RAM[54][0] ;
 wire \RAM[54][1] ;
 wire \RAM[54][2] ;
 wire \RAM[54][3] ;
 wire \RAM[54][4] ;
 wire \RAM[54][5] ;
 wire \RAM[54][6] ;
 wire \RAM[54][7] ;
 wire \RAM[55][0] ;
 wire \RAM[55][1] ;
 wire \RAM[55][2] ;
 wire \RAM[55][3] ;
 wire \RAM[55][4] ;
 wire \RAM[55][5] ;
 wire \RAM[55][6] ;
 wire \RAM[55][7] ;
 wire \RAM[56][0] ;
 wire \RAM[56][1] ;
 wire \RAM[56][2] ;
 wire \RAM[56][3] ;
 wire \RAM[56][4] ;
 wire \RAM[56][5] ;
 wire \RAM[56][6] ;
 wire \RAM[56][7] ;
 wire \RAM[57][0] ;
 wire \RAM[57][1] ;
 wire \RAM[57][2] ;
 wire \RAM[57][3] ;
 wire \RAM[57][4] ;
 wire \RAM[57][5] ;
 wire \RAM[57][6] ;
 wire \RAM[57][7] ;
 wire \RAM[58][0] ;
 wire \RAM[58][1] ;
 wire \RAM[58][2] ;
 wire \RAM[58][3] ;
 wire \RAM[58][4] ;
 wire \RAM[58][5] ;
 wire \RAM[58][6] ;
 wire \RAM[58][7] ;
 wire \RAM[59][0] ;
 wire \RAM[59][1] ;
 wire \RAM[59][2] ;
 wire \RAM[59][3] ;
 wire \RAM[59][4] ;
 wire \RAM[59][5] ;
 wire \RAM[59][6] ;
 wire \RAM[59][7] ;
 wire \RAM[5][0] ;
 wire \RAM[5][1] ;
 wire \RAM[5][2] ;
 wire \RAM[5][3] ;
 wire \RAM[5][4] ;
 wire \RAM[5][5] ;
 wire \RAM[5][6] ;
 wire \RAM[5][7] ;
 wire \RAM[60][0] ;
 wire \RAM[60][1] ;
 wire \RAM[60][2] ;
 wire \RAM[60][3] ;
 wire \RAM[60][4] ;
 wire \RAM[60][5] ;
 wire \RAM[60][6] ;
 wire \RAM[60][7] ;
 wire \RAM[61][0] ;
 wire \RAM[61][1] ;
 wire \RAM[61][2] ;
 wire \RAM[61][3] ;
 wire \RAM[61][4] ;
 wire \RAM[61][5] ;
 wire \RAM[61][6] ;
 wire \RAM[61][7] ;
 wire \RAM[62][0] ;
 wire \RAM[62][1] ;
 wire \RAM[62][2] ;
 wire \RAM[62][3] ;
 wire \RAM[62][4] ;
 wire \RAM[62][5] ;
 wire \RAM[62][6] ;
 wire \RAM[62][7] ;
 wire \RAM[63][0] ;
 wire \RAM[63][1] ;
 wire \RAM[63][2] ;
 wire \RAM[63][3] ;
 wire \RAM[63][4] ;
 wire \RAM[63][5] ;
 wire \RAM[63][6] ;
 wire \RAM[63][7] ;
 wire \RAM[6][0] ;
 wire \RAM[6][1] ;
 wire \RAM[6][2] ;
 wire \RAM[6][3] ;
 wire \RAM[6][4] ;
 wire \RAM[6][5] ;
 wire \RAM[6][6] ;
 wire \RAM[6][7] ;
 wire \RAM[7][0] ;
 wire \RAM[7][1] ;
 wire \RAM[7][2] ;
 wire \RAM[7][3] ;
 wire \RAM[7][4] ;
 wire \RAM[7][5] ;
 wire \RAM[7][6] ;
 wire \RAM[7][7] ;
 wire \RAM[8][0] ;
 wire \RAM[8][1] ;
 wire \RAM[8][2] ;
 wire \RAM[8][3] ;
 wire \RAM[8][4] ;
 wire \RAM[8][5] ;
 wire \RAM[8][6] ;
 wire \RAM[8][7] ;
 wire \RAM[9][0] ;
 wire \RAM[9][1] ;
 wire \RAM[9][2] ;
 wire \RAM[9][3] ;
 wire \RAM[9][4] ;
 wire \RAM[9][5] ;
 wire \RAM[9][6] ;
 wire \RAM[9][7] ;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire \addr_read[0] ;
 wire \addr_read[1] ;
 wire \addr_read[2] ;
 wire \addr_read[3] ;
 wire \addr_write[0] ;
 wire \addr_write[1] ;
 wire \addr_write[2] ;
 wire \addr_write[3] ;
 wire \addr_write[4] ;
 wire \addr_write[5] ;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;
 wire \combined_out[0] ;
 wire \combined_out[1] ;
 wire \combined_out[2] ;
 wire \combined_out[3] ;
 wire \combined_out[4] ;
 wire \combined_out[5] ;
 wire \combined_out[6] ;
 wire \combined_out[7] ;
 wire \data_to_write[0] ;
 wire \data_to_write[1] ;
 wire \data_to_write[2] ;
 wire \data_to_write[3] ;
 wire \data_to_write[4] ;
 wire \data_to_write[5] ;
 wire \data_to_write[6] ;
 wire \data_to_write[7] ;
 wire \genblk1[0].sel_byte ;
 wire \genblk1[0].wr_en_this_byte ;
 wire \genblk1[10].sel_byte ;
 wire \genblk1[10].wr_en_this_byte ;
 wire \genblk1[11].sel_byte ;
 wire \genblk1[11].wr_en_this_byte ;
 wire \genblk1[12].sel_byte ;
 wire \genblk1[12].wr_en_this_byte ;
 wire \genblk1[13].sel_byte ;
 wire \genblk1[13].wr_en_this_byte ;
 wire \genblk1[14].sel_byte ;
 wire \genblk1[14].wr_en_this_byte ;
 wire \genblk1[15].sel_byte ;
 wire \genblk1[15].wr_en_this_byte ;
 wire \genblk1[16].sel_byte ;
 wire \genblk1[16].wr_en_this_byte ;
 wire \genblk1[17].sel_byte ;
 wire \genblk1[17].wr_en_this_byte ;
 wire \genblk1[18].sel_byte ;
 wire \genblk1[18].wr_en_this_byte ;
 wire \genblk1[19].sel_byte ;
 wire \genblk1[19].wr_en_this_byte ;
 wire \genblk1[1].sel_byte ;
 wire \genblk1[1].wr_en_this_byte ;
 wire \genblk1[20].sel_byte ;
 wire \genblk1[20].wr_en_this_byte ;
 wire \genblk1[21].sel_byte ;
 wire \genblk1[21].wr_en_this_byte ;
 wire \genblk1[22].sel_byte ;
 wire \genblk1[22].wr_en_this_byte ;
 wire \genblk1[23].sel_byte ;
 wire \genblk1[23].wr_en_this_byte ;
 wire \genblk1[24].sel_byte ;
 wire \genblk1[24].wr_en_this_byte ;
 wire \genblk1[25].sel_byte ;
 wire \genblk1[25].wr_en_this_byte ;
 wire \genblk1[26].sel_byte ;
 wire \genblk1[26].wr_en_this_byte ;
 wire \genblk1[27].sel_byte ;
 wire \genblk1[27].wr_en_this_byte ;
 wire \genblk1[28].sel_byte ;
 wire \genblk1[28].wr_en_this_byte ;
 wire \genblk1[29].sel_byte ;
 wire \genblk1[29].wr_en_this_byte ;
 wire \genblk1[2].sel_byte ;
 wire \genblk1[2].wr_en_this_byte ;
 wire \genblk1[30].sel_byte ;
 wire \genblk1[30].wr_en_this_byte ;
 wire \genblk1[31].sel_byte ;
 wire \genblk1[31].wr_en_this_byte ;
 wire \genblk1[32].sel_byte ;
 wire \genblk1[32].wr_en_this_byte ;
 wire \genblk1[33].sel_byte ;
 wire \genblk1[33].wr_en_this_byte ;
 wire \genblk1[34].sel_byte ;
 wire \genblk1[34].wr_en_this_byte ;
 wire \genblk1[35].sel_byte ;
 wire \genblk1[35].wr_en_this_byte ;
 wire \genblk1[36].sel_byte ;
 wire \genblk1[36].wr_en_this_byte ;
 wire \genblk1[37].sel_byte ;
 wire \genblk1[37].wr_en_this_byte ;
 wire \genblk1[38].sel_byte ;
 wire \genblk1[38].wr_en_this_byte ;
 wire \genblk1[39].sel_byte ;
 wire \genblk1[39].wr_en_this_byte ;
 wire \genblk1[3].sel_byte ;
 wire \genblk1[3].wr_en_this_byte ;
 wire \genblk1[40].sel_byte ;
 wire \genblk1[40].wr_en_this_byte ;
 wire \genblk1[41].sel_byte ;
 wire \genblk1[41].wr_en_this_byte ;
 wire \genblk1[42].sel_byte ;
 wire \genblk1[42].wr_en_this_byte ;
 wire \genblk1[43].sel_byte ;
 wire \genblk1[43].wr_en_this_byte ;
 wire \genblk1[44].sel_byte ;
 wire \genblk1[44].wr_en_this_byte ;
 wire \genblk1[45].sel_byte ;
 wire \genblk1[45].wr_en_this_byte ;
 wire \genblk1[46].sel_byte ;
 wire \genblk1[46].wr_en_this_byte ;
 wire \genblk1[47].sel_byte ;
 wire \genblk1[47].wr_en_this_byte ;
 wire \genblk1[48].sel_byte ;
 wire \genblk1[48].wr_en_this_byte ;
 wire \genblk1[49].sel_byte ;
 wire \genblk1[49].wr_en_this_byte ;
 wire \genblk1[4].sel_byte ;
 wire \genblk1[4].wr_en_this_byte ;
 wire \genblk1[50].sel_byte ;
 wire \genblk1[50].wr_en_this_byte ;
 wire \genblk1[51].sel_byte ;
 wire \genblk1[51].wr_en_this_byte ;
 wire \genblk1[52].sel_byte ;
 wire \genblk1[52].wr_en_this_byte ;
 wire \genblk1[53].sel_byte ;
 wire \genblk1[53].wr_en_this_byte ;
 wire \genblk1[54].sel_byte ;
 wire \genblk1[54].wr_en_this_byte ;
 wire \genblk1[55].sel_byte ;
 wire \genblk1[55].wr_en_this_byte ;
 wire \genblk1[56].sel_byte ;
 wire \genblk1[56].wr_en_this_byte ;
 wire \genblk1[57].sel_byte ;
 wire \genblk1[57].wr_en_this_byte ;
 wire \genblk1[58].sel_byte ;
 wire \genblk1[58].wr_en_this_byte ;
 wire \genblk1[59].sel_byte ;
 wire \genblk1[59].wr_en_this_byte ;
 wire \genblk1[5].sel_byte ;
 wire \genblk1[5].wr_en_this_byte ;
 wire \genblk1[60].sel_byte ;
 wire \genblk1[60].wr_en_this_byte ;
 wire \genblk1[61].sel_byte ;
 wire \genblk1[61].wr_en_this_byte ;
 wire \genblk1[62].sel_byte ;
 wire \genblk1[62].wr_en_this_byte ;
 wire \genblk1[63].sel_byte ;
 wire \genblk1[63].wr_en_this_byte ;
 wire \genblk1[6].sel_byte ;
 wire \genblk1[6].wr_en_this_byte ;
 wire \genblk1[7].sel_byte ;
 wire \genblk1[7].wr_en_this_byte ;
 wire \genblk1[8].sel_byte ;
 wire \genblk1[8].wr_en_this_byte ;
 wire \genblk1[9].sel_byte ;
 wire \genblk1[9].wr_en_this_byte ;
 wire \genblk2[0].partition_sel_n ;
 wire \genblk2[0].selected_out[0] ;
 wire \genblk2[0].selected_out[1] ;
 wire \genblk2[0].selected_out[2] ;
 wire \genblk2[0].selected_out[3] ;
 wire \genblk2[0].selected_out[4] ;
 wire \genblk2[0].selected_out[5] ;
 wire \genblk2[0].selected_out[6] ;
 wire \genblk2[0].selected_out[7] ;
 wire \genblk2[1].partition_sel_n ;
 wire \genblk2[1].selected_out[0] ;
 wire \genblk2[1].selected_out[1] ;
 wire \genblk2[1].selected_out[2] ;
 wire \genblk2[1].selected_out[3] ;
 wire \genblk2[1].selected_out[4] ;
 wire \genblk2[1].selected_out[5] ;
 wire \genblk2[1].selected_out[6] ;
 wire \genblk2[1].selected_out[7] ;
 wire \genblk2[2].partition_sel_n ;
 wire \genblk2[2].selected_out[0] ;
 wire \genblk2[2].selected_out[1] ;
 wire \genblk2[2].selected_out[2] ;
 wire \genblk2[2].selected_out[3] ;
 wire \genblk2[2].selected_out[4] ;
 wire \genblk2[2].selected_out[5] ;
 wire \genblk2[2].selected_out[6] ;
 wire \genblk2[2].selected_out[7] ;
 wire \genblk2[3].partition_sel_n ;
 wire \genblk2[3].selected_out[0] ;
 wire \genblk2[3].selected_out[1] ;
 wire \genblk2[3].selected_out[2] ;
 wire \genblk2[3].selected_out[3] ;
 wire \genblk2[3].selected_out[4] ;
 wire \genblk2[3].selected_out[5] ;
 wire \genblk2[3].selected_out[6] ;
 wire \genblk2[3].selected_out[7] ;
 wire net1;
 wire net10;
 wire net11;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net2;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net3;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net4;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net5;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net6;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire wr_en;
 wire wr_en_next;
 wire wr_en_ok;
 wire wr_en_valid;

 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(_0052_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(_0053_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(_0056_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(_0127_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(_0163_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(\combined_out[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(ui_in[4]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(\data_to_write[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(\data_to_write[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_0_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_0_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_0_210 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_0_214 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_0_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_241 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_0_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_0_275 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_287 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_0_303 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_0_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_320 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_332 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_0_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_10_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_149 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_10_165 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_180 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_10_189 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_216 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_10_229 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_268 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_10_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_10_305 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_10_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_68 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_10_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_11_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_11_190 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_198 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_218 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_237 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_11_277 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_11_293 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_11_315 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_11_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_123 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_174 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_18 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_233 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_12_275 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_12_290 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_294 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_12_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_92 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_13_135 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_13_165 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_181 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_13_205 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_13_220 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_13_265 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_13_332 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_13_43 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_115 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_14_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_229 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_14_249 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_14_265 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_14_280 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_14_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_14_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_14_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_92 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_15_135 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_15_156 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_160 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_205 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_263 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_15_277 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_306 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_61 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_115 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_127 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_16_144 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_174 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_16_241 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_260 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_16_305 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_108 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_143 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_186 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_17_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_17_256 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_17_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_314 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_116 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_18_131 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_18_187 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_19_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_220 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_19_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_261 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_19_274 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_19_299 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_19_44 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_19_64 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_1_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_1_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_155 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_1_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_184 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_209 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_1_286 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_1_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_1_305 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_1_329 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_1_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_1_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_124 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_131 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_20_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_145 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_20_173 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_221 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_20_236 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_20_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_73 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_80 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_21_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_119 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_21_154 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_21_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_21_177 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_21_192 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_21_207 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_214 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_231 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_241 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_21_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_21_260 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_264 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_21_278 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_297 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_21_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_80 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_100 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_132 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_155 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_22_177 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_183 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_200 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_22_214 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_221 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_22_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_22_233 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_239 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_119 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_23_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_23_18 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_23_191 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_23_222 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_23_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_23_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_23_293 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_23_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_23_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_23_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_78 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_112 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_24_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_24_162 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_24_200 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_204 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_212 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_24_218 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_24_226 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_24_237 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_24_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_24_275 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_24_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_24_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_321 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_24_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_24_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_108 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_25_149 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_155 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_175 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_191 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_25_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_25_217 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_25_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_229 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_25_236 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_25_263 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_25_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_297 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_25_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_25_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_26_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_160 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_18 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_189 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_26_203 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_211 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_215 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_26_222 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_228 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_232 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_26_244 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_26_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_36 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_58 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_71 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_27_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_27_165 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_27_188 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_27_204 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_27_212 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_27_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_229 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_27_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_239 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_27_249 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_27_300 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_27_52 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_28_18 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_28_180 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_28_187 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_28_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_28_201 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_205 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_219 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_231 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_28_246 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_28_275 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_321 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_28_42 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_94 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_135 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_29_159 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_189 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_29_202 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_210 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_29_216 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_29_231 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_293 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_306 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_52 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_120 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_2_161 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_165 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_178 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_2_18 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_2_192 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_294 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_2_299 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_2_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_2_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_48 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_2_62 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_66 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_2_79 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_99 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_132 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_165 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_178 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_30_203 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_30_218 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_238 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_290 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_306 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_321 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_42 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_150 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_31_200 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_31_211 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_291 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_295 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_6 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_89 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_32_112 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_129 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_32_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_200 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_32_215 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_221 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_269 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_98 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_33_204 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_262 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_33_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_75 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_87 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_34_121 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_135 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_34_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_168 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_191 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_34_220 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_247 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_34_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_34_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_264 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_294 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_71 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_103 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_122 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_147 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_222 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_240 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_262 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_122 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_145 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_164 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_20 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_36_234 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_36_300 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_36_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_36_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_36_90 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_104 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_37_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_157 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_160 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_312 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_182 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_222 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_306 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_3_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_3_140 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_3_156 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_3_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_3_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_3_221 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_3_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_3_276 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_287 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_297 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_3_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_34 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_48 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_4_107 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_4_164 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_4_179 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_4_288 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_292 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_4_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_4_305 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_4_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_4_332 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_4_48 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_52 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_94 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_5_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_147 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_5_209 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_5_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_30 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_123 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_6_176 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_244 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_6_265 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_6_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_313 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_98 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_7_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_18 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_199 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_7_221 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_7_261 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_7_277 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_7_288 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_7_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_7_312 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_95 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_8_100 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_148 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_168 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_18 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_8_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_201 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_219 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_8_234 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_8_249 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_289 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_8_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_8_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_8_331 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_8_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_155 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_9_175 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_9_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_42 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_49 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_50 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_52 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_56 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_58 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_40 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_59 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_60 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_61 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_62 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_63 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_64 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_66 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_67 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_68 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_70 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_71 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_72 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_73 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_74 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_75 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_76 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_42 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_43 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_44 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_45 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_46 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_47 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_48 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_78 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_79 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_80 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_81 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_82 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_83 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_84 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_85 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_86 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_87 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_88 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_138 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_139 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_140 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_141 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_142 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_143 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_144 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_145 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_146 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_147 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_148 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_149 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_150 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_151 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_152 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_153 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_154 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_155 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_156 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_157 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_158 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_159 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_160 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_161 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_162 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_163 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_164 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_165 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_166 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_167 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_168 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_169 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_170 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_171 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_172 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_173 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_174 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_175 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_176 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_177 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_178 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_179 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_180 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_181 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_182 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_183 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_184 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_185 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_186 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_187 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_188 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_189 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_190 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_191 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_192 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_89 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_90 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_91 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_92 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_93 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_193 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_194 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_195 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_196 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_197 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_198 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_199 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_200 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_201 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_202 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_203 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_204 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_205 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_206 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_207 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_208 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_209 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_210 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_211 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_212 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_213 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_214 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_215 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_216 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_217 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_218 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_219 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_220 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_221 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_222 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_223 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_224 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_225 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_226 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_227 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_228 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_229 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_230 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_231 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_232 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_233 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_234 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_235 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_236 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_237 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_238 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_239 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_240 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_241 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_242 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_243 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_244 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_245 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_246 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_247 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_94 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_95 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_96 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_97 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_98 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_99 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_248 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_249 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_250 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_251 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_252 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_253 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_254 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_255 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_256 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_257 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_258 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_259 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_260 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_261 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_262 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_263 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_264 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_265 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_266 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_267 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_268 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_269 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_270 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_271 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_272 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_273 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_274 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_275 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_276 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_277 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_278 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_279 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_280 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_281 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_282 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_283 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_284 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_285 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_286 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_287 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_288 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_289 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_290 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_291 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_292 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_293 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_294 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_295 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_296 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_297 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_298 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_299 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_300 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_301 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_302 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_100 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_101 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_102 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_103 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_104 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_105 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_106 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_107 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_108 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_109 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_110 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_111 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_112 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_113 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_114 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_115 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_116 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_117 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_118 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_119 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_120 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_121 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_122 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_123 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_124 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_125 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_126 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_127 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_128 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_129 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_130 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_131 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_132 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_133 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_134 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_135 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_136 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_137 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__or2_1 _0456_ (.A(net6),
    .B(net7),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0210_));
 sky130_fd_sc_hd__clkbuf_1 _0457_ (.A(_0210_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0000_));
 sky130_fd_sc_hd__or2b_1 _0458_ (.A(net7),
    .B_N(net6),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0211_));
 sky130_fd_sc_hd__clkbuf_1 _0459_ (.A(_0211_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0001_));
 sky130_fd_sc_hd__or2b_1 _0460_ (.A(net6),
    .B_N(net7),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0212_));
 sky130_fd_sc_hd__clkbuf_1 _0461_ (.A(_0212_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0002_));
 sky130_fd_sc_hd__nand2_1 _0462_ (.A(net6),
    .B(net7),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0003_));
 sky130_fd_sc_hd__inv_2 _0463_ (.A(wr_en_valid),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0004_));
 sky130_fd_sc_hd__or4_4 _0464_ (.A(\addr_write[0] ),
    .B(\addr_write[1] ),
    .C(\addr_write[2] ),
    .D(\addr_write[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0213_));
 sky130_fd_sc_hd__or2_1 _0465_ (.A(\addr_write[4] ),
    .B(\addr_write[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0214_));
 sky130_fd_sc_hd__clkbuf_2 _0466_ (.A(_0214_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0215_));
 sky130_fd_sc_hd__buf_2 _0467_ (.A(_0215_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0216_));
 sky130_fd_sc_hd__nor2_1 _0468_ (.A(_0213_),
    .B(_0216_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].sel_byte ));
 sky130_fd_sc_hd__clkbuf_4 _0469_ (.A(\addr_write[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0217_));
 sky130_fd_sc_hd__or4b_4 _0470_ (.A(\addr_write[1] ),
    .B(\addr_write[2] ),
    .C(\addr_write[3] ),
    .D_N(_0217_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0218_));
 sky130_fd_sc_hd__nor2_1 _0471_ (.A(_0216_),
    .B(_0218_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].sel_byte ));
 sky130_fd_sc_hd__clkbuf_4 _0472_ (.A(\addr_write[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0219_));
 sky130_fd_sc_hd__or4b_4 _0473_ (.A(\addr_write[0] ),
    .B(\addr_write[2] ),
    .C(\addr_write[3] ),
    .D_N(_0219_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0220_));
 sky130_fd_sc_hd__nor2_1 _0474_ (.A(_0216_),
    .B(_0220_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].sel_byte ));
 sky130_fd_sc_hd__buf_4 _0475_ (.A(\addr_write[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0221_));
 sky130_fd_sc_hd__buf_4 _0476_ (.A(\addr_write[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0222_));
 sky130_fd_sc_hd__nand2_1 _0477_ (.A(\addr_write[0] ),
    .B(\addr_write[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0223_));
 sky130_fd_sc_hd__or3_2 _0478_ (.A(_0221_),
    .B(_0222_),
    .C(_0223_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0224_));
 sky130_fd_sc_hd__nor2_1 _0479_ (.A(_0216_),
    .B(_0224_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].sel_byte ));
 sky130_fd_sc_hd__or4b_4 _0480_ (.A(\addr_write[0] ),
    .B(\addr_write[1] ),
    .C(\addr_write[3] ),
    .D_N(\addr_write[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0225_));
 sky130_fd_sc_hd__nor2_1 _0481_ (.A(_0216_),
    .B(_0225_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].sel_byte ));
 sky130_fd_sc_hd__or4bb_4 _0482_ (.A(_0219_),
    .B(_0222_),
    .C_N(_0221_),
    .D_N(_0217_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0226_));
 sky130_fd_sc_hd__nor2_1 _0483_ (.A(_0216_),
    .B(_0226_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].sel_byte ));
 sky130_fd_sc_hd__or4bb_4 _0484_ (.A(_0217_),
    .B(_0222_),
    .C_N(_0221_),
    .D_N(_0219_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0227_));
 sky130_fd_sc_hd__nor2_1 _0485_ (.A(_0216_),
    .B(_0227_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].sel_byte ));
 sky130_fd_sc_hd__or3b_2 _0486_ (.A(\addr_write[3] ),
    .B(_0223_),
    .C_N(\addr_write[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0228_));
 sky130_fd_sc_hd__nor2_1 _0487_ (.A(_0216_),
    .B(_0228_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].sel_byte ));
 sky130_fd_sc_hd__or4b_2 _0488_ (.A(\addr_write[0] ),
    .B(\addr_write[1] ),
    .C(\addr_write[2] ),
    .D_N(\addr_write[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0229_));
 sky130_fd_sc_hd__nor2_1 _0489_ (.A(_0216_),
    .B(_0229_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[8].sel_byte ));
 sky130_fd_sc_hd__or4bb_4 _0490_ (.A(_0219_),
    .B(_0221_),
    .C_N(_0222_),
    .D_N(_0217_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0230_));
 sky130_fd_sc_hd__nor2_1 _0491_ (.A(_0216_),
    .B(_0230_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[9].sel_byte ));
 sky130_fd_sc_hd__or4bb_4 _0492_ (.A(_0217_),
    .B(_0221_),
    .C_N(_0222_),
    .D_N(_0219_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0231_));
 sky130_fd_sc_hd__nor2_1 _0493_ (.A(_0215_),
    .B(_0231_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[10].sel_byte ));
 sky130_fd_sc_hd__or3b_2 _0494_ (.A(_0223_),
    .B(\addr_write[2] ),
    .C_N(\addr_write[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0232_));
 sky130_fd_sc_hd__nor2_1 _0495_ (.A(_0215_),
    .B(_0232_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[11].sel_byte ));
 sky130_fd_sc_hd__or4bb_4 _0496_ (.A(_0217_),
    .B(_0219_),
    .C_N(_0221_),
    .D_N(_0222_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0233_));
 sky130_fd_sc_hd__nor2_1 _0497_ (.A(_0215_),
    .B(_0233_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[12].sel_byte ));
 sky130_fd_sc_hd__nand4b_4 _0498_ (.A_N(_0219_),
    .B(_0221_),
    .C(_0222_),
    .D(_0217_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0234_));
 sky130_fd_sc_hd__nor2_1 _0499_ (.A(_0215_),
    .B(_0234_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[13].sel_byte ));
 sky130_fd_sc_hd__nand4b_4 _0500_ (.A_N(_0217_),
    .B(_0219_),
    .C(_0221_),
    .D(_0222_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0235_));
 sky130_fd_sc_hd__nor2_1 _0501_ (.A(_0215_),
    .B(_0235_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[14].sel_byte ));
 sky130_fd_sc_hd__nand4_4 _0502_ (.A(_0217_),
    .B(_0219_),
    .C(_0221_),
    .D(_0222_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0236_));
 sky130_fd_sc_hd__nor2_1 _0503_ (.A(_0215_),
    .B(_0236_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[15].sel_byte ));
 sky130_fd_sc_hd__or2b_1 _0504_ (.A(\addr_write[5] ),
    .B_N(\addr_write[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0237_));
 sky130_fd_sc_hd__clkbuf_2 _0505_ (.A(_0237_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0238_));
 sky130_fd_sc_hd__buf_2 _0506_ (.A(_0238_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0239_));
 sky130_fd_sc_hd__nor2_1 _0507_ (.A(_0213_),
    .B(_0239_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[16].sel_byte ));
 sky130_fd_sc_hd__nor2_1 _0508_ (.A(_0218_),
    .B(_0239_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[17].sel_byte ));
 sky130_fd_sc_hd__nor2_1 _0509_ (.A(_0220_),
    .B(_0239_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[18].sel_byte ));
 sky130_fd_sc_hd__nor2_1 _0510_ (.A(_0224_),
    .B(_0239_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[19].sel_byte ));
 sky130_fd_sc_hd__nor2_1 _0511_ (.A(_0225_),
    .B(_0239_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[20].sel_byte ));
 sky130_fd_sc_hd__nor2_1 _0512_ (.A(_0226_),
    .B(_0239_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[21].sel_byte ));
 sky130_fd_sc_hd__nor2_1 _0513_ (.A(_0227_),
    .B(_0239_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[22].sel_byte ));
 sky130_fd_sc_hd__nor2_1 _0514_ (.A(_0228_),
    .B(_0239_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[23].sel_byte ));
 sky130_fd_sc_hd__nor2_1 _0515_ (.A(_0229_),
    .B(_0239_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[24].sel_byte ));
 sky130_fd_sc_hd__nor2_1 _0516_ (.A(_0230_),
    .B(_0239_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[25].sel_byte ));
 sky130_fd_sc_hd__nor2_1 _0517_ (.A(_0231_),
    .B(_0238_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[26].sel_byte ));
 sky130_fd_sc_hd__nor2_1 _0518_ (.A(_0232_),
    .B(_0238_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[27].sel_byte ));
 sky130_fd_sc_hd__nor2_1 _0519_ (.A(_0233_),
    .B(_0238_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[28].sel_byte ));
 sky130_fd_sc_hd__nor2_1 _0520_ (.A(_0234_),
    .B(_0238_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[29].sel_byte ));
 sky130_fd_sc_hd__nor2_1 _0521_ (.A(_0235_),
    .B(_0238_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[30].sel_byte ));
 sky130_fd_sc_hd__nor2_1 _0522_ (.A(_0236_),
    .B(_0238_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[31].sel_byte ));
 sky130_fd_sc_hd__or2b_1 _0523_ (.A(\addr_write[4] ),
    .B_N(\addr_write[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0240_));
 sky130_fd_sc_hd__clkbuf_2 _0524_ (.A(_0240_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0241_));
 sky130_fd_sc_hd__buf_2 _0525_ (.A(_0241_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0242_));
 sky130_fd_sc_hd__nor2_1 _0526_ (.A(_0213_),
    .B(_0242_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[32].sel_byte ));
 sky130_fd_sc_hd__nor2_1 _0527_ (.A(_0218_),
    .B(_0242_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[33].sel_byte ));
 sky130_fd_sc_hd__nor2_1 _0528_ (.A(_0220_),
    .B(_0242_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[34].sel_byte ));
 sky130_fd_sc_hd__nor2_1 _0529_ (.A(_0224_),
    .B(_0242_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[35].sel_byte ));
 sky130_fd_sc_hd__nor2_1 _0530_ (.A(_0225_),
    .B(_0242_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[36].sel_byte ));
 sky130_fd_sc_hd__nor2_1 _0531_ (.A(_0226_),
    .B(_0242_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[37].sel_byte ));
 sky130_fd_sc_hd__nor2_1 _0532_ (.A(_0227_),
    .B(_0242_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[38].sel_byte ));
 sky130_fd_sc_hd__nor2_1 _0533_ (.A(_0228_),
    .B(_0242_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[39].sel_byte ));
 sky130_fd_sc_hd__nor2_1 _0534_ (.A(_0229_),
    .B(_0242_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[40].sel_byte ));
 sky130_fd_sc_hd__nor2_1 _0535_ (.A(_0230_),
    .B(_0242_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[41].sel_byte ));
 sky130_fd_sc_hd__nor2_1 _0536_ (.A(_0231_),
    .B(_0241_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[42].sel_byte ));
 sky130_fd_sc_hd__nor2_1 _0537_ (.A(_0232_),
    .B(_0241_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[43].sel_byte ));
 sky130_fd_sc_hd__nor2_1 _0538_ (.A(_0233_),
    .B(_0241_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[44].sel_byte ));
 sky130_fd_sc_hd__nor2_1 _0539_ (.A(_0234_),
    .B(_0241_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[45].sel_byte ));
 sky130_fd_sc_hd__nor2_1 _0540_ (.A(_0235_),
    .B(_0241_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[46].sel_byte ));
 sky130_fd_sc_hd__nor2_1 _0541_ (.A(_0236_),
    .B(_0241_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[47].sel_byte ));
 sky130_fd_sc_hd__nand2_2 _0542_ (.A(\addr_write[4] ),
    .B(\addr_write[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0243_));
 sky130_fd_sc_hd__buf_2 _0543_ (.A(_0243_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0244_));
 sky130_fd_sc_hd__nor2_1 _0544_ (.A(_0213_),
    .B(_0244_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[48].sel_byte ));
 sky130_fd_sc_hd__nor2_1 _0545_ (.A(_0218_),
    .B(_0244_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[49].sel_byte ));
 sky130_fd_sc_hd__nor2_1 _0546_ (.A(_0220_),
    .B(_0244_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[50].sel_byte ));
 sky130_fd_sc_hd__nor2_1 _0547_ (.A(_0224_),
    .B(_0244_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[51].sel_byte ));
 sky130_fd_sc_hd__nor2_1 _0548_ (.A(_0225_),
    .B(_0244_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[52].sel_byte ));
 sky130_fd_sc_hd__nor2_1 _0549_ (.A(_0226_),
    .B(_0244_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[53].sel_byte ));
 sky130_fd_sc_hd__nor2_1 _0550_ (.A(_0227_),
    .B(_0244_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[54].sel_byte ));
 sky130_fd_sc_hd__nor2_1 _0551_ (.A(_0228_),
    .B(_0244_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[55].sel_byte ));
 sky130_fd_sc_hd__nor2_1 _0552_ (.A(_0229_),
    .B(_0244_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[56].sel_byte ));
 sky130_fd_sc_hd__nor2_1 _0553_ (.A(_0230_),
    .B(_0244_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[57].sel_byte ));
 sky130_fd_sc_hd__nor2_1 _0554_ (.A(_0231_),
    .B(_0243_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[58].sel_byte ));
 sky130_fd_sc_hd__nor2_1 _0555_ (.A(_0232_),
    .B(_0243_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[59].sel_byte ));
 sky130_fd_sc_hd__nor2_1 _0556_ (.A(_0233_),
    .B(_0243_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[60].sel_byte ));
 sky130_fd_sc_hd__nor2_1 _0557_ (.A(_0234_),
    .B(_0243_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[61].sel_byte ));
 sky130_fd_sc_hd__nor2_1 _0558_ (.A(_0235_),
    .B(_0243_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[62].sel_byte ));
 sky130_fd_sc_hd__nor2_1 _0559_ (.A(_0236_),
    .B(_0243_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[63].sel_byte ));
 sky130_fd_sc_hd__and2_1 _0560_ (.A(wr_en_valid),
    .B(wr_en_ok),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0245_));
 sky130_fd_sc_hd__clkbuf_1 _0561_ (.A(_0245_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(wr_en));
 sky130_fd_sc_hd__and4bb_2 _0562_ (.A_N(\addr_read[3] ),
    .B_N(\addr_read[1] ),
    .C(\addr_read[0] ),
    .D(\addr_read[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0246_));
 sky130_fd_sc_hd__buf_4 _0563_ (.A(_0246_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0247_));
 sky130_fd_sc_hd__clkbuf_4 _0564_ (.A(_0247_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0248_));
 sky130_fd_sc_hd__buf_2 _0565_ (.A(\addr_read[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0249_));
 sky130_fd_sc_hd__buf_2 _0566_ (.A(\addr_read[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0250_));
 sky130_fd_sc_hd__buf_2 _0567_ (.A(\addr_read[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0251_));
 sky130_fd_sc_hd__buf_2 _0568_ (.A(\addr_read[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0252_));
 sky130_fd_sc_hd__and4bb_2 _0569_ (.A_N(_0249_),
    .B_N(_0250_),
    .C(_0251_),
    .D(_0252_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0253_));
 sky130_fd_sc_hd__buf_4 _0570_ (.A(_0253_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0254_));
 sky130_fd_sc_hd__buf_4 _0571_ (.A(_0254_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0255_));
 sky130_fd_sc_hd__and4_2 _0572_ (.A(_0249_),
    .B(\addr_read[3] ),
    .C(\addr_read[0] ),
    .D(\addr_read[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0256_));
 sky130_fd_sc_hd__buf_4 _0573_ (.A(_0256_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0257_));
 sky130_fd_sc_hd__clkbuf_4 _0574_ (.A(_0257_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0258_));
 sky130_fd_sc_hd__and4b_2 _0575_ (.A_N(\addr_read[2] ),
    .B(_0250_),
    .C(_0251_),
    .D(_0252_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0259_));
 sky130_fd_sc_hd__clkbuf_4 _0576_ (.A(_0259_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0260_));
 sky130_fd_sc_hd__buf_4 _0577_ (.A(_0260_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0261_));
 sky130_fd_sc_hd__a22o_1 _0578_ (.A1(\RAM[47][0] ),
    .A2(_0258_),
    .B1(_0261_),
    .B2(\RAM[43][0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0262_));
 sky130_fd_sc_hd__a221o_1 _0579_ (.A1(\RAM[37][0] ),
    .A2(_0248_),
    .B1(_0255_),
    .B2(\RAM[35][0] ),
    .C1(_0262_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0263_));
 sky130_fd_sc_hd__nor4b_1 _0580_ (.A(_0250_),
    .B(_0251_),
    .C(_0252_),
    .D_N(_0249_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0264_));
 sky130_fd_sc_hd__clkbuf_4 _0581_ (.A(net28),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0265_));
 sky130_fd_sc_hd__and4bb_2 _0582_ (.A_N(\addr_read[2] ),
    .B_N(\addr_read[1] ),
    .C(_0251_),
    .D(_0250_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0266_));
 sky130_fd_sc_hd__buf_4 _0583_ (.A(_0266_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0267_));
 sky130_fd_sc_hd__nor4b_2 _0584_ (.A(\addr_read[2] ),
    .B(\addr_read[3] ),
    .C(_0251_),
    .D_N(\addr_read[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0268_));
 sky130_fd_sc_hd__nor4b_4 _0585_ (.A(_0249_),
    .B(_0250_),
    .C(_0252_),
    .D_N(\addr_read[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0269_));
 sky130_fd_sc_hd__a22o_1 _0586_ (.A1(\RAM[34][0] ),
    .A2(_0268_),
    .B1(_0269_),
    .B2(\RAM[33][0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0270_));
 sky130_fd_sc_hd__a221o_1 _0587_ (.A1(\RAM[36][0] ),
    .A2(_0265_),
    .B1(_0267_),
    .B2(\RAM[41][0] ),
    .C1(_0270_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0271_));
 sky130_fd_sc_hd__and4b_2 _0588_ (.A_N(_0251_),
    .B(_0252_),
    .C(_0249_),
    .D(_0250_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0272_));
 sky130_fd_sc_hd__buf_4 _0589_ (.A(_0272_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0273_));
 sky130_fd_sc_hd__and4b_2 _0590_ (.A_N(_0252_),
    .B(_0251_),
    .C(_0250_),
    .D(_0249_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0274_));
 sky130_fd_sc_hd__buf_4 _0591_ (.A(_0274_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0275_));
 sky130_fd_sc_hd__and4bb_2 _0592_ (.A_N(\addr_read[3] ),
    .B_N(\addr_read[0] ),
    .C(\addr_read[1] ),
    .D(\addr_read[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0276_));
 sky130_fd_sc_hd__nor4_1 _0593_ (.A(_0249_),
    .B(_0250_),
    .C(_0251_),
    .D(_0252_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0277_));
 sky130_fd_sc_hd__a22o_1 _0594_ (.A1(\RAM[38][0] ),
    .A2(_0276_),
    .B1(net26),
    .B2(\RAM[32][0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0278_));
 sky130_fd_sc_hd__a221o_1 _0595_ (.A1(\RAM[46][0] ),
    .A2(_0273_),
    .B1(_0275_),
    .B2(\RAM[45][0] ),
    .C1(_0278_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0279_));
 sky130_fd_sc_hd__nor4b_1 _0596_ (.A(_0249_),
    .B(_0251_),
    .C(_0252_),
    .D_N(\addr_read[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0280_));
 sky130_fd_sc_hd__clkbuf_4 _0597_ (.A(net25),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0281_));
 sky130_fd_sc_hd__and4bb_2 _0598_ (.A_N(_0249_),
    .B_N(\addr_read[0] ),
    .C(_0252_),
    .D(_0250_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0282_));
 sky130_fd_sc_hd__buf_4 _0599_ (.A(_0282_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0283_));
 sky130_fd_sc_hd__and4b_2 _0600_ (.A_N(\addr_read[3] ),
    .B(\addr_read[0] ),
    .C(\addr_read[1] ),
    .D(\addr_read[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0284_));
 sky130_fd_sc_hd__clkbuf_4 _0601_ (.A(_0284_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0285_));
 sky130_fd_sc_hd__and4bb_2 _0602_ (.A_N(\addr_read[0] ),
    .B_N(\addr_read[1] ),
    .C(\addr_read[2] ),
    .D(\addr_read[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0286_));
 sky130_fd_sc_hd__buf_4 _0603_ (.A(_0286_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0287_));
 sky130_fd_sc_hd__a22o_1 _0604_ (.A1(\RAM[39][0] ),
    .A2(_0285_),
    .B1(_0287_),
    .B2(\RAM[44][0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0288_));
 sky130_fd_sc_hd__a221o_1 _0605_ (.A1(\RAM[40][0] ),
    .A2(_0281_),
    .B1(_0283_),
    .B2(\RAM[42][0] ),
    .C1(_0288_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0289_));
 sky130_fd_sc_hd__or3_1 _0606_ (.A(_0271_),
    .B(_0279_),
    .C(_0289_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0290_));
 sky130_fd_sc_hd__or2_1 _0607_ (.A(_0263_),
    .B(_0290_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0291_));
 sky130_fd_sc_hd__clkbuf_1 _0608_ (.A(_0291_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk2[2].selected_out[0] ));
 sky130_fd_sc_hd__a22o_1 _0609_ (.A1(\RAM[39][1] ),
    .A2(_0285_),
    .B1(_0287_),
    .B2(\RAM[44][1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0292_));
 sky130_fd_sc_hd__buf_4 _0610_ (.A(_0246_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0293_));
 sky130_fd_sc_hd__clkbuf_4 _0611_ (.A(_0276_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0294_));
 sky130_fd_sc_hd__a22o_1 _0612_ (.A1(\RAM[37][1] ),
    .A2(_0293_),
    .B1(_0294_),
    .B2(\RAM[38][1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0295_));
 sky130_fd_sc_hd__buf_4 _0613_ (.A(_0274_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0296_));
 sky130_fd_sc_hd__a22o_1 _0614_ (.A1(\RAM[47][1] ),
    .A2(_0257_),
    .B1(_0296_),
    .B2(\RAM[45][1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0297_));
 sky130_fd_sc_hd__a22o_1 _0615_ (.A1(\RAM[35][1] ),
    .A2(_0254_),
    .B1(_0281_),
    .B2(\RAM[40][1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0298_));
 sky130_fd_sc_hd__or4_1 _0616_ (.A(_0292_),
    .B(_0295_),
    .C(_0297_),
    .D(_0298_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0299_));
 sky130_fd_sc_hd__buf_4 _0617_ (.A(_0269_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0300_));
 sky130_fd_sc_hd__clkbuf_4 _0618_ (.A(_0300_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0301_));
 sky130_fd_sc_hd__buf_4 _0619_ (.A(net26),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0302_));
 sky130_fd_sc_hd__clkbuf_4 _0620_ (.A(_0302_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0303_));
 sky130_fd_sc_hd__buf_4 _0621_ (.A(_0266_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0304_));
 sky130_fd_sc_hd__clkbuf_4 _0622_ (.A(_0304_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0305_));
 sky130_fd_sc_hd__a22o_1 _0623_ (.A1(\RAM[46][1] ),
    .A2(_0273_),
    .B1(_0305_),
    .B2(\RAM[41][1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0306_));
 sky130_fd_sc_hd__a221o_1 _0624_ (.A1(\RAM[33][1] ),
    .A2(_0301_),
    .B1(_0303_),
    .B2(\RAM[32][1] ),
    .C1(_0306_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0307_));
 sky130_fd_sc_hd__buf_4 _0625_ (.A(_0268_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0308_));
 sky130_fd_sc_hd__buf_4 _0626_ (.A(_0308_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0309_));
 sky130_fd_sc_hd__clkbuf_4 _0627_ (.A(_0265_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0310_));
 sky130_fd_sc_hd__clkbuf_4 _0628_ (.A(_0283_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0311_));
 sky130_fd_sc_hd__a22o_1 _0629_ (.A1(\RAM[43][1] ),
    .A2(_0261_),
    .B1(_0311_),
    .B2(\RAM[42][1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0312_));
 sky130_fd_sc_hd__a221o_1 _0630_ (.A1(\RAM[34][1] ),
    .A2(_0309_),
    .B1(_0310_),
    .B2(\RAM[36][1] ),
    .C1(_0312_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0313_));
 sky130_fd_sc_hd__or3_1 _0631_ (.A(_0299_),
    .B(_0307_),
    .C(_0313_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0314_));
 sky130_fd_sc_hd__clkbuf_1 _0632_ (.A(_0314_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk2[2].selected_out[1] ));
 sky130_fd_sc_hd__buf_4 _0633_ (.A(_0260_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0315_));
 sky130_fd_sc_hd__buf_4 _0634_ (.A(_0286_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0316_));
 sky130_fd_sc_hd__a22o_1 _0635_ (.A1(\RAM[37][2] ),
    .A2(_0247_),
    .B1(_0316_),
    .B2(\RAM[44][2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0317_));
 sky130_fd_sc_hd__a221o_1 _0636_ (.A1(\RAM[43][2] ),
    .A2(_0315_),
    .B1(_0301_),
    .B2(\RAM[33][2] ),
    .C1(_0317_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0318_));
 sky130_fd_sc_hd__buf_4 _0637_ (.A(_0281_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0319_));
 sky130_fd_sc_hd__buf_4 _0638_ (.A(_0319_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0320_));
 sky130_fd_sc_hd__buf_4 _0639_ (.A(_0296_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0321_));
 sky130_fd_sc_hd__buf_4 _0640_ (.A(_0284_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0322_));
 sky130_fd_sc_hd__a22o_1 _0641_ (.A1(\RAM[34][2] ),
    .A2(_0308_),
    .B1(_0322_),
    .B2(\RAM[39][2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0323_));
 sky130_fd_sc_hd__a221o_1 _0642_ (.A1(\RAM[40][2] ),
    .A2(_0320_),
    .B1(_0321_),
    .B2(\RAM[45][2] ),
    .C1(_0323_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0324_));
 sky130_fd_sc_hd__a22o_1 _0643_ (.A1(\RAM[47][2] ),
    .A2(_0257_),
    .B1(_0272_),
    .B2(\RAM[46][2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0325_));
 sky130_fd_sc_hd__a22o_1 _0644_ (.A1(\RAM[41][2] ),
    .A2(_0304_),
    .B1(_0283_),
    .B2(\RAM[42][2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0326_));
 sky130_fd_sc_hd__clkbuf_4 _0645_ (.A(net26),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0327_));
 sky130_fd_sc_hd__a22o_1 _0646_ (.A1(\RAM[35][2] ),
    .A2(_0254_),
    .B1(_0327_),
    .B2(\RAM[32][2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0328_));
 sky130_fd_sc_hd__a22o_1 _0647_ (.A1(\RAM[38][2] ),
    .A2(_0294_),
    .B1(_0265_),
    .B2(\RAM[36][2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0329_));
 sky130_fd_sc_hd__or4_1 _0648_ (.A(_0325_),
    .B(_0326_),
    .C(_0328_),
    .D(_0329_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0330_));
 sky130_fd_sc_hd__or3_1 _0649_ (.A(_0318_),
    .B(_0324_),
    .C(_0330_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0331_));
 sky130_fd_sc_hd__clkbuf_1 _0650_ (.A(_0331_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk2[2].selected_out[2] ));
 sky130_fd_sc_hd__a22o_1 _0651_ (.A1(\RAM[37][3] ),
    .A2(_0247_),
    .B1(_0311_),
    .B2(\RAM[42][3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0332_));
 sky130_fd_sc_hd__a221o_1 _0652_ (.A1(\RAM[43][3] ),
    .A2(_0315_),
    .B1(_0301_),
    .B2(\RAM[33][3] ),
    .C1(_0332_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0333_));
 sky130_fd_sc_hd__buf_4 _0653_ (.A(_0276_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0334_));
 sky130_fd_sc_hd__a22o_1 _0654_ (.A1(\RAM[39][3] ),
    .A2(_0284_),
    .B1(_0266_),
    .B2(\RAM[41][3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0335_));
 sky130_fd_sc_hd__a221o_1 _0655_ (.A1(\RAM[38][3] ),
    .A2(_0334_),
    .B1(_0327_),
    .B2(\RAM[32][3] ),
    .C1(_0335_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0336_));
 sky130_fd_sc_hd__a22o_1 _0656_ (.A1(\RAM[47][3] ),
    .A2(_0256_),
    .B1(net25),
    .B2(\RAM[40][3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0337_));
 sky130_fd_sc_hd__a221o_1 _0657_ (.A1(\RAM[36][3] ),
    .A2(_0265_),
    .B1(_0316_),
    .B2(\RAM[44][3] ),
    .C1(_0337_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0338_));
 sky130_fd_sc_hd__buf_4 _0658_ (.A(_0253_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0339_));
 sky130_fd_sc_hd__buf_4 _0659_ (.A(_0268_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0340_));
 sky130_fd_sc_hd__a22o_1 _0660_ (.A1(\RAM[34][3] ),
    .A2(_0340_),
    .B1(_0274_),
    .B2(\RAM[45][3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0341_));
 sky130_fd_sc_hd__a221o_1 _0661_ (.A1(\RAM[35][3] ),
    .A2(_0339_),
    .B1(_0273_),
    .B2(\RAM[46][3] ),
    .C1(_0341_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0342_));
 sky130_fd_sc_hd__or3_1 _0662_ (.A(_0336_),
    .B(_0338_),
    .C(_0342_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0343_));
 sky130_fd_sc_hd__or2_1 _0663_ (.A(_0333_),
    .B(_0343_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0344_));
 sky130_fd_sc_hd__clkbuf_1 _0664_ (.A(_0344_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk2[2].selected_out[3] ));
 sky130_fd_sc_hd__buf_4 _0665_ (.A(_0257_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0345_));
 sky130_fd_sc_hd__clkbuf_4 _0666_ (.A(_0272_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0346_));
 sky130_fd_sc_hd__a22o_1 _0667_ (.A1(\RAM[34][4] ),
    .A2(_0308_),
    .B1(_0346_),
    .B2(\RAM[46][4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0347_));
 sky130_fd_sc_hd__a221o_1 _0668_ (.A1(\RAM[47][4] ),
    .A2(_0345_),
    .B1(_0320_),
    .B2(\RAM[40][4] ),
    .C1(_0347_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0348_));
 sky130_fd_sc_hd__a22o_1 _0669_ (.A1(\RAM[37][4] ),
    .A2(_0246_),
    .B1(_0287_),
    .B2(\RAM[44][4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0349_));
 sky130_fd_sc_hd__a221o_1 _0670_ (.A1(\RAM[38][4] ),
    .A2(_0294_),
    .B1(_0265_),
    .B2(\RAM[36][4] ),
    .C1(_0349_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0350_));
 sky130_fd_sc_hd__a22o_1 _0671_ (.A1(\RAM[39][4] ),
    .A2(_0285_),
    .B1(_0266_),
    .B2(\RAM[41][4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0351_));
 sky130_fd_sc_hd__a221o_1 _0672_ (.A1(\RAM[35][4] ),
    .A2(_0339_),
    .B1(_0296_),
    .B2(\RAM[45][4] ),
    .C1(_0351_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0352_));
 sky130_fd_sc_hd__clkbuf_4 _0673_ (.A(_0300_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0353_));
 sky130_fd_sc_hd__a22o_1 _0674_ (.A1(\RAM[43][4] ),
    .A2(_0259_),
    .B1(_0283_),
    .B2(\RAM[42][4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0354_));
 sky130_fd_sc_hd__a221o_1 _0675_ (.A1(\RAM[33][4] ),
    .A2(_0353_),
    .B1(_0302_),
    .B2(\RAM[32][4] ),
    .C1(_0354_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0355_));
 sky130_fd_sc_hd__or3_1 _0676_ (.A(_0350_),
    .B(_0352_),
    .C(_0355_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0356_));
 sky130_fd_sc_hd__or2_1 _0677_ (.A(_0348_),
    .B(_0356_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0357_));
 sky130_fd_sc_hd__clkbuf_1 _0678_ (.A(_0357_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk2[2].selected_out[4] ));
 sky130_fd_sc_hd__a22o_1 _0679_ (.A1(\RAM[35][5] ),
    .A2(_0253_),
    .B1(_0304_),
    .B2(\RAM[41][5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0358_));
 sky130_fd_sc_hd__a22o_1 _0680_ (.A1(\RAM[39][5] ),
    .A2(_0285_),
    .B1(_0260_),
    .B2(\RAM[43][5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0359_));
 sky130_fd_sc_hd__a22o_1 _0681_ (.A1(\RAM[34][5] ),
    .A2(_0340_),
    .B1(_0281_),
    .B2(\RAM[40][5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0360_));
 sky130_fd_sc_hd__a22o_1 _0682_ (.A1(\RAM[38][5] ),
    .A2(_0294_),
    .B1(_0265_),
    .B2(\RAM[36][5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0361_));
 sky130_fd_sc_hd__or4_1 _0683_ (.A(_0358_),
    .B(_0359_),
    .C(_0360_),
    .D(_0361_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0362_));
 sky130_fd_sc_hd__a22o_1 _0684_ (.A1(\RAM[46][5] ),
    .A2(_0273_),
    .B1(_0275_),
    .B2(\RAM[45][5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0363_));
 sky130_fd_sc_hd__a221o_1 _0685_ (.A1(\RAM[47][5] ),
    .A2(_0345_),
    .B1(_0301_),
    .B2(\RAM[33][5] ),
    .C1(_0363_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0364_));
 sky130_fd_sc_hd__clkbuf_4 _0686_ (.A(_0316_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0365_));
 sky130_fd_sc_hd__a22o_1 _0687_ (.A1(\RAM[32][5] ),
    .A2(_0302_),
    .B1(_0311_),
    .B2(\RAM[42][5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0366_));
 sky130_fd_sc_hd__a221o_1 _0688_ (.A1(\RAM[37][5] ),
    .A2(_0248_),
    .B1(_0365_),
    .B2(\RAM[44][5] ),
    .C1(_0366_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0367_));
 sky130_fd_sc_hd__or3_1 _0689_ (.A(_0362_),
    .B(_0364_),
    .C(_0367_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0368_));
 sky130_fd_sc_hd__clkbuf_1 _0690_ (.A(_0368_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk2[2].selected_out[5] ));
 sky130_fd_sc_hd__clkbuf_4 _0691_ (.A(_0322_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0369_));
 sky130_fd_sc_hd__buf_4 _0692_ (.A(net28),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0370_));
 sky130_fd_sc_hd__a22o_1 _0693_ (.A1(\RAM[34][6] ),
    .A2(_0308_),
    .B1(_0370_),
    .B2(\RAM[36][6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0371_));
 sky130_fd_sc_hd__a221o_1 _0694_ (.A1(\RAM[39][6] ),
    .A2(_0369_),
    .B1(_0321_),
    .B2(\RAM[45][6] ),
    .C1(_0371_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0372_));
 sky130_fd_sc_hd__a22o_1 _0695_ (.A1(\RAM[43][6] ),
    .A2(_0259_),
    .B1(_0272_),
    .B2(\RAM[46][6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0373_));
 sky130_fd_sc_hd__a221o_1 _0696_ (.A1(\RAM[35][6] ),
    .A2(_0254_),
    .B1(_0353_),
    .B2(\RAM[33][6] ),
    .C1(_0373_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0374_));
 sky130_fd_sc_hd__a22o_1 _0697_ (.A1(\RAM[37][6] ),
    .A2(_0246_),
    .B1(net25),
    .B2(\RAM[40][6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0375_));
 sky130_fd_sc_hd__a221o_1 _0698_ (.A1(\RAM[41][6] ),
    .A2(_0304_),
    .B1(_0316_),
    .B2(\RAM[44][6] ),
    .C1(_0375_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0376_));
 sky130_fd_sc_hd__a22o_1 _0699_ (.A1(\RAM[47][6] ),
    .A2(_0257_),
    .B1(_0282_),
    .B2(\RAM[42][6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0377_));
 sky130_fd_sc_hd__a221o_1 _0700_ (.A1(\RAM[38][6] ),
    .A2(_0334_),
    .B1(_0302_),
    .B2(\RAM[32][6] ),
    .C1(_0377_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0378_));
 sky130_fd_sc_hd__or3_1 _0701_ (.A(_0374_),
    .B(_0376_),
    .C(_0378_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0379_));
 sky130_fd_sc_hd__or2_1 _0702_ (.A(_0372_),
    .B(_0379_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0380_));
 sky130_fd_sc_hd__clkbuf_1 _0703_ (.A(_0380_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk2[2].selected_out[6] ));
 sky130_fd_sc_hd__a22o_1 _0704_ (.A1(\RAM[38][7] ),
    .A2(_0334_),
    .B1(_0311_),
    .B2(\RAM[42][7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0381_));
 sky130_fd_sc_hd__a221o_1 _0705_ (.A1(\RAM[43][7] ),
    .A2(_0315_),
    .B1(_0310_),
    .B2(\RAM[36][7] ),
    .C1(_0381_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0382_));
 sky130_fd_sc_hd__a22o_1 _0706_ (.A1(\RAM[37][7] ),
    .A2(_0247_),
    .B1(_0275_),
    .B2(\RAM[45][7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0383_));
 sky130_fd_sc_hd__a221o_1 _0707_ (.A1(\RAM[32][7] ),
    .A2(_0302_),
    .B1(_0365_),
    .B2(\RAM[44][7] ),
    .C1(_0383_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0384_));
 sky130_fd_sc_hd__a22o_1 _0708_ (.A1(\RAM[33][7] ),
    .A2(_0300_),
    .B1(_0304_),
    .B2(\RAM[41][7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0385_));
 sky130_fd_sc_hd__a22o_1 _0709_ (.A1(\RAM[47][7] ),
    .A2(_0257_),
    .B1(_0273_),
    .B2(\RAM[46][7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0386_));
 sky130_fd_sc_hd__a22o_1 _0710_ (.A1(\RAM[34][7] ),
    .A2(_0340_),
    .B1(_0254_),
    .B2(\RAM[35][7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0387_));
 sky130_fd_sc_hd__a22o_1 _0711_ (.A1(\RAM[39][7] ),
    .A2(_0322_),
    .B1(_0281_),
    .B2(\RAM[40][7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0388_));
 sky130_fd_sc_hd__or4_1 _0712_ (.A(_0385_),
    .B(_0386_),
    .C(_0387_),
    .D(_0388_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0389_));
 sky130_fd_sc_hd__or3_1 _0713_ (.A(_0382_),
    .B(_0384_),
    .C(_0389_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0390_));
 sky130_fd_sc_hd__clkbuf_1 _0714_ (.A(_0390_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk2[2].selected_out[7] ));
 sky130_fd_sc_hd__clkbuf_4 _0715_ (.A(_0283_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0391_));
 sky130_fd_sc_hd__a22o_1 _0716_ (.A1(\RAM[54][0] ),
    .A2(_0334_),
    .B1(_0305_),
    .B2(\RAM[57][0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0392_));
 sky130_fd_sc_hd__a221o_1 _0717_ (.A1(\RAM[56][0] ),
    .A2(_0320_),
    .B1(_0391_),
    .B2(\RAM[58][0] ),
    .C1(_0392_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0393_));
 sky130_fd_sc_hd__a22o_1 _0718_ (.A1(\RAM[49][0] ),
    .A2(_0269_),
    .B1(net115),
    .B2(\RAM[52][0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0394_));
 sky130_fd_sc_hd__a221o_1 _0719_ (.A1(\RAM[55][0] ),
    .A2(_0322_),
    .B1(_0339_),
    .B2(\RAM[51][0] ),
    .C1(_0394_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0395_));
 sky130_fd_sc_hd__a22o_1 _0720_ (.A1(\RAM[63][0] ),
    .A2(_0256_),
    .B1(_0293_),
    .B2(\RAM[53][0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0396_));
 sky130_fd_sc_hd__a221o_1 _0721_ (.A1(\RAM[48][0] ),
    .A2(_0327_),
    .B1(_0296_),
    .B2(\RAM[61][0] ),
    .C1(_0396_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0397_));
 sky130_fd_sc_hd__a22o_1 _0722_ (.A1(\RAM[62][0] ),
    .A2(_0272_),
    .B1(_0287_),
    .B2(\RAM[60][0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0398_));
 sky130_fd_sc_hd__a221o_1 _0723_ (.A1(\RAM[50][0] ),
    .A2(_0308_),
    .B1(_0261_),
    .B2(\RAM[59][0] ),
    .C1(_0398_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0399_));
 sky130_fd_sc_hd__or3_1 _0724_ (.A(_0395_),
    .B(_0397_),
    .C(_0399_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0400_));
 sky130_fd_sc_hd__or2_1 _0725_ (.A(_0393_),
    .B(_0400_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0401_));
 sky130_fd_sc_hd__clkbuf_1 _0726_ (.A(_0401_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk2[3].selected_out[0] ));
 sky130_fd_sc_hd__a22o_1 _0727_ (.A1(\RAM[62][1] ),
    .A2(_0346_),
    .B1(_0275_),
    .B2(\RAM[61][1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0402_));
 sky130_fd_sc_hd__a221o_1 _0728_ (.A1(\RAM[52][1] ),
    .A2(_0310_),
    .B1(_0391_),
    .B2(\RAM[58][1] ),
    .C1(_0402_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0403_));
 sky130_fd_sc_hd__a22o_1 _0729_ (.A1(\RAM[63][1] ),
    .A2(_0256_),
    .B1(_0253_),
    .B2(\RAM[51][1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0404_));
 sky130_fd_sc_hd__a221o_1 _0730_ (.A1(\RAM[50][1] ),
    .A2(_0308_),
    .B1(_0327_),
    .B2(\RAM[48][1] ),
    .C1(_0404_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0405_));
 sky130_fd_sc_hd__a22o_1 _0731_ (.A1(\RAM[59][1] ),
    .A2(_0259_),
    .B1(_0294_),
    .B2(\RAM[54][1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0406_));
 sky130_fd_sc_hd__a221o_1 _0732_ (.A1(\RAM[55][1] ),
    .A2(_0322_),
    .B1(_0316_),
    .B2(\RAM[60][1] ),
    .C1(_0406_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0407_));
 sky130_fd_sc_hd__a22o_1 _0733_ (.A1(\RAM[56][1] ),
    .A2(net114),
    .B1(_0304_),
    .B2(\RAM[57][1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0408_));
 sky130_fd_sc_hd__a221o_1 _0734_ (.A1(\RAM[53][1] ),
    .A2(_0247_),
    .B1(_0353_),
    .B2(\RAM[49][1] ),
    .C1(_0408_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0409_));
 sky130_fd_sc_hd__or3_1 _0735_ (.A(_0405_),
    .B(_0407_),
    .C(_0409_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0410_));
 sky130_fd_sc_hd__or2_1 _0736_ (.A(_0403_),
    .B(_0410_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0411_));
 sky130_fd_sc_hd__clkbuf_1 _0737_ (.A(_0411_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk2[3].selected_out[1] ));
 sky130_fd_sc_hd__a22o_1 _0738_ (.A1(\RAM[52][2] ),
    .A2(_0310_),
    .B1(_0302_),
    .B2(\RAM[48][2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0412_));
 sky130_fd_sc_hd__a22o_1 _0739_ (.A1(\RAM[53][2] ),
    .A2(_0248_),
    .B1(_0369_),
    .B2(\RAM[55][2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0413_));
 sky130_fd_sc_hd__a22o_1 _0740_ (.A1(\RAM[50][2] ),
    .A2(_0308_),
    .B1(_0283_),
    .B2(\RAM[58][2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0414_));
 sky130_fd_sc_hd__a221o_1 _0741_ (.A1(\RAM[59][2] ),
    .A2(_0315_),
    .B1(_0321_),
    .B2(\RAM[61][2] ),
    .C1(_0414_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0415_));
 sky130_fd_sc_hd__a2111o_1 _0742_ (.A1(\RAM[51][2] ),
    .A2(_0255_),
    .B1(_0412_),
    .C1(_0413_),
    .D1(_0415_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0416_));
 sky130_fd_sc_hd__buf_4 _0743_ (.A(_0334_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0417_));
 sky130_fd_sc_hd__a22o_1 _0744_ (.A1(\RAM[49][2] ),
    .A2(_0353_),
    .B1(_0346_),
    .B2(\RAM[62][2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0418_));
 sky130_fd_sc_hd__a221o_1 _0745_ (.A1(\RAM[54][2] ),
    .A2(_0417_),
    .B1(_0365_),
    .B2(\RAM[60][2] ),
    .C1(_0418_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0419_));
 sky130_fd_sc_hd__a221o_1 _0746_ (.A1(\RAM[63][2] ),
    .A2(_0345_),
    .B1(_0305_),
    .B2(\RAM[57][2] ),
    .C1(_0419_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0420_));
 sky130_fd_sc_hd__a211o_1 _0747_ (.A1(\RAM[56][2] ),
    .A2(_0320_),
    .B1(_0416_),
    .C1(_0420_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk2[3].selected_out[2] ));
 sky130_fd_sc_hd__buf_4 _0748_ (.A(_0273_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0421_));
 sky130_fd_sc_hd__a22o_1 _0749_ (.A1(\RAM[51][3] ),
    .A2(_0339_),
    .B1(_0319_),
    .B2(\RAM[56][3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0422_));
 sky130_fd_sc_hd__a221o_1 _0750_ (.A1(\RAM[54][3] ),
    .A2(_0417_),
    .B1(_0421_),
    .B2(\RAM[62][3] ),
    .C1(_0422_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0423_));
 sky130_fd_sc_hd__a22o_1 _0751_ (.A1(\RAM[63][3] ),
    .A2(_0258_),
    .B1(_0305_),
    .B2(\RAM[57][3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0424_));
 sky130_fd_sc_hd__a221o_1 _0752_ (.A1(\RAM[59][3] ),
    .A2(_0315_),
    .B1(_0391_),
    .B2(\RAM[58][3] ),
    .C1(_0424_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0425_));
 sky130_fd_sc_hd__a22o_1 _0753_ (.A1(\RAM[61][3] ),
    .A2(_0274_),
    .B1(_0287_),
    .B2(\RAM[60][3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0426_));
 sky130_fd_sc_hd__a22o_1 _0754_ (.A1(\RAM[50][3] ),
    .A2(_0340_),
    .B1(_0265_),
    .B2(\RAM[52][3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0427_));
 sky130_fd_sc_hd__a22o_1 _0755_ (.A1(\RAM[49][3] ),
    .A2(_0300_),
    .B1(_0327_),
    .B2(\RAM[48][3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0428_));
 sky130_fd_sc_hd__a22o_1 _0756_ (.A1(\RAM[53][3] ),
    .A2(_0293_),
    .B1(_0322_),
    .B2(\RAM[55][3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0429_));
 sky130_fd_sc_hd__or4_1 _0757_ (.A(_0426_),
    .B(_0427_),
    .C(_0428_),
    .D(_0429_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0430_));
 sky130_fd_sc_hd__or3_1 _0758_ (.A(_0423_),
    .B(_0425_),
    .C(_0430_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0431_));
 sky130_fd_sc_hd__clkbuf_1 _0759_ (.A(_0431_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk2[3].selected_out[3] ));
 sky130_fd_sc_hd__a22o_1 _0760_ (.A1(\RAM[63][4] ),
    .A2(_0258_),
    .B1(_0346_),
    .B2(\RAM[62][4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0432_));
 sky130_fd_sc_hd__a221o_1 _0761_ (.A1(\RAM[57][4] ),
    .A2(_0305_),
    .B1(_0365_),
    .B2(\RAM[60][4] ),
    .C1(_0432_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0433_));
 sky130_fd_sc_hd__a22o_1 _0762_ (.A1(\RAM[54][4] ),
    .A2(_0334_),
    .B1(_0339_),
    .B2(\RAM[51][4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0434_));
 sky130_fd_sc_hd__a221o_1 _0763_ (.A1(\RAM[53][4] ),
    .A2(_0248_),
    .B1(_0391_),
    .B2(\RAM[58][4] ),
    .C1(_0434_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0435_));
 sky130_fd_sc_hd__a22o_1 _0764_ (.A1(\RAM[50][4] ),
    .A2(_0340_),
    .B1(_0327_),
    .B2(\RAM[48][4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0436_));
 sky130_fd_sc_hd__a22o_1 _0765_ (.A1(\RAM[55][4] ),
    .A2(_0285_),
    .B1(_0281_),
    .B2(\RAM[56][4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0437_));
 sky130_fd_sc_hd__a22o_1 _0766_ (.A1(\RAM[52][4] ),
    .A2(_0265_),
    .B1(_0296_),
    .B2(\RAM[61][4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0438_));
 sky130_fd_sc_hd__a22o_1 _0767_ (.A1(\RAM[59][4] ),
    .A2(_0260_),
    .B1(_0300_),
    .B2(\RAM[49][4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0439_));
 sky130_fd_sc_hd__or4_1 _0768_ (.A(_0436_),
    .B(_0437_),
    .C(_0438_),
    .D(_0439_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0440_));
 sky130_fd_sc_hd__or3_1 _0769_ (.A(_0433_),
    .B(_0435_),
    .C(_0440_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0441_));
 sky130_fd_sc_hd__clkbuf_1 _0770_ (.A(_0441_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk2[3].selected_out[4] ));
 sky130_fd_sc_hd__a22o_1 _0771_ (.A1(\RAM[54][5] ),
    .A2(_0334_),
    .B1(_0346_),
    .B2(\RAM[62][5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0442_));
 sky130_fd_sc_hd__a221o_1 _0772_ (.A1(\RAM[59][5] ),
    .A2(_0315_),
    .B1(_0310_),
    .B2(\RAM[52][5] ),
    .C1(_0442_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0443_));
 sky130_fd_sc_hd__a22o_1 _0773_ (.A1(\RAM[55][5] ),
    .A2(_0284_),
    .B1(_0282_),
    .B2(\RAM[58][5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0444_));
 sky130_fd_sc_hd__a221o_1 _0774_ (.A1(\RAM[51][5] ),
    .A2(_0254_),
    .B1(_0296_),
    .B2(\RAM[61][5] ),
    .C1(_0444_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0445_));
 sky130_fd_sc_hd__a22o_1 _0775_ (.A1(\RAM[49][5] ),
    .A2(_0269_),
    .B1(_0287_),
    .B2(\RAM[60][5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0446_));
 sky130_fd_sc_hd__a221o_1 _0776_ (.A1(\RAM[53][5] ),
    .A2(_0293_),
    .B1(_0319_),
    .B2(\RAM[56][5] ),
    .C1(_0446_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0447_));
 sky130_fd_sc_hd__a22o_1 _0777_ (.A1(\RAM[63][5] ),
    .A2(_0257_),
    .B1(_0277_),
    .B2(\RAM[48][5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0448_));
 sky130_fd_sc_hd__a221o_1 _0778_ (.A1(\RAM[50][5] ),
    .A2(_0308_),
    .B1(_0267_),
    .B2(\RAM[57][5] ),
    .C1(_0448_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0449_));
 sky130_fd_sc_hd__or3_1 _0779_ (.A(_0445_),
    .B(_0447_),
    .C(_0449_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0450_));
 sky130_fd_sc_hd__or2_1 _0780_ (.A(_0443_),
    .B(_0450_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0451_));
 sky130_fd_sc_hd__clkbuf_1 _0781_ (.A(_0451_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk2[3].selected_out[5] ));
 sky130_fd_sc_hd__a22o_1 _0782_ (.A1(\RAM[59][6] ),
    .A2(_0261_),
    .B1(_0319_),
    .B2(\RAM[56][6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0452_));
 sky130_fd_sc_hd__a221o_1 _0783_ (.A1(\RAM[48][6] ),
    .A2(_0302_),
    .B1(_0321_),
    .B2(\RAM[61][6] ),
    .C1(_0452_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0453_));
 sky130_fd_sc_hd__a22o_1 _0784_ (.A1(\RAM[55][6] ),
    .A2(_0322_),
    .B1(_0267_),
    .B2(\RAM[57][6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0454_));
 sky130_fd_sc_hd__a221o_1 _0785_ (.A1(\RAM[50][6] ),
    .A2(_0309_),
    .B1(_0391_),
    .B2(\RAM[58][6] ),
    .C1(_0454_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0455_));
 sky130_fd_sc_hd__a22o_1 _0786_ (.A1(\RAM[51][6] ),
    .A2(_0254_),
    .B1(_0287_),
    .B2(\RAM[60][6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0022_));
 sky130_fd_sc_hd__a22o_1 _0787_ (.A1(\RAM[63][6] ),
    .A2(_0257_),
    .B1(_0293_),
    .B2(\RAM[53][6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0023_));
 sky130_fd_sc_hd__a22o_1 _0788_ (.A1(\RAM[54][6] ),
    .A2(_0294_),
    .B1(_0273_),
    .B2(\RAM[62][6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0024_));
 sky130_fd_sc_hd__a22o_1 _0789_ (.A1(\RAM[49][6] ),
    .A2(_0300_),
    .B1(_0265_),
    .B2(\RAM[52][6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0025_));
 sky130_fd_sc_hd__or4_1 _0790_ (.A(_0022_),
    .B(_0023_),
    .C(_0024_),
    .D(_0025_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0026_));
 sky130_fd_sc_hd__or3_1 _0791_ (.A(_0453_),
    .B(_0455_),
    .C(_0026_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0027_));
 sky130_fd_sc_hd__clkbuf_1 _0792_ (.A(_0027_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk2[3].selected_out[6] ));
 sky130_fd_sc_hd__a22o_1 _0793_ (.A1(\RAM[63][7] ),
    .A2(_0258_),
    .B1(_0370_),
    .B2(\RAM[52][7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0028_));
 sky130_fd_sc_hd__a221o_1 _0794_ (.A1(\RAM[51][7] ),
    .A2(_0255_),
    .B1(_0320_),
    .B2(\RAM[56][7] ),
    .C1(_0028_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0029_));
 sky130_fd_sc_hd__a22o_1 _0795_ (.A1(\RAM[59][7] ),
    .A2(_0259_),
    .B1(_0269_),
    .B2(\RAM[49][7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0030_));
 sky130_fd_sc_hd__a221o_1 _0796_ (.A1(\RAM[62][7] ),
    .A2(_0273_),
    .B1(_0296_),
    .B2(\RAM[61][7] ),
    .C1(_0030_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0031_));
 sky130_fd_sc_hd__a22o_1 _0797_ (.A1(\RAM[55][7] ),
    .A2(_0284_),
    .B1(_0287_),
    .B2(\RAM[60][7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0032_));
 sky130_fd_sc_hd__a221o_1 _0798_ (.A1(\RAM[54][7] ),
    .A2(_0334_),
    .B1(_0267_),
    .B2(\RAM[57][7] ),
    .C1(_0032_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0033_));
 sky130_fd_sc_hd__a22o_1 _0799_ (.A1(\RAM[53][7] ),
    .A2(_0246_),
    .B1(_0282_),
    .B2(\RAM[58][7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0034_));
 sky130_fd_sc_hd__a221o_1 _0800_ (.A1(\RAM[50][7] ),
    .A2(_0308_),
    .B1(_0327_),
    .B2(\RAM[48][7] ),
    .C1(_0034_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0035_));
 sky130_fd_sc_hd__or3_1 _0801_ (.A(_0031_),
    .B(_0033_),
    .C(_0035_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0036_));
 sky130_fd_sc_hd__or2_1 _0802_ (.A(_0029_),
    .B(_0036_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0037_));
 sky130_fd_sc_hd__clkbuf_1 _0803_ (.A(_0037_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk2[3].selected_out[7] ));
 sky130_fd_sc_hd__a22o_1 _0804_ (.A1(\RAM[31][0] ),
    .A2(_0258_),
    .B1(_0339_),
    .B2(\RAM[19][0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0038_));
 sky130_fd_sc_hd__a221o_1 _0805_ (.A1(\RAM[25][0] ),
    .A2(_0305_),
    .B1(_0391_),
    .B2(\RAM[26][0] ),
    .C1(_0038_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0039_));
 sky130_fd_sc_hd__a22o_1 _0806_ (.A1(\RAM[17][0] ),
    .A2(_0353_),
    .B1(_0370_),
    .B2(\RAM[20][0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0040_));
 sky130_fd_sc_hd__a221o_1 _0807_ (.A1(\RAM[27][0] ),
    .A2(_0315_),
    .B1(_0321_),
    .B2(\RAM[29][0] ),
    .C1(_0040_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0041_));
 sky130_fd_sc_hd__a22o_1 _0808_ (.A1(\RAM[22][0] ),
    .A2(_0294_),
    .B1(net26),
    .B2(\RAM[16][0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0042_));
 sky130_fd_sc_hd__a22o_1 _0809_ (.A1(\RAM[18][0] ),
    .A2(_0340_),
    .B1(_0293_),
    .B2(\RAM[21][0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0043_));
 sky130_fd_sc_hd__a22o_1 _0810_ (.A1(\RAM[23][0] ),
    .A2(_0285_),
    .B1(_0281_),
    .B2(\RAM[24][0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0044_));
 sky130_fd_sc_hd__a22o_1 _0811_ (.A1(\RAM[30][0] ),
    .A2(_0273_),
    .B1(_0316_),
    .B2(\RAM[28][0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0045_));
 sky130_fd_sc_hd__or4_1 _0812_ (.A(_0042_),
    .B(_0043_),
    .C(_0044_),
    .D(_0045_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0046_));
 sky130_fd_sc_hd__or3_1 _0813_ (.A(_0039_),
    .B(_0041_),
    .C(_0046_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0047_));
 sky130_fd_sc_hd__clkbuf_1 _0814_ (.A(_0047_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk2[1].selected_out[0] ));
 sky130_fd_sc_hd__a22o_1 _0815_ (.A1(\RAM[17][1] ),
    .A2(_0353_),
    .B1(_0370_),
    .B2(\RAM[20][1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0048_));
 sky130_fd_sc_hd__a221o_1 _0816_ (.A1(\RAM[27][1] ),
    .A2(_0315_),
    .B1(_0421_),
    .B2(\RAM[30][1] ),
    .C1(_0048_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0049_));
 sky130_fd_sc_hd__a22o_1 _0817_ (.A1(\RAM[31][1] ),
    .A2(_0258_),
    .B1(_0311_),
    .B2(\RAM[26][1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0050_));
 sky130_fd_sc_hd__a221o_1 _0818_ (.A1(\RAM[24][1] ),
    .A2(_0320_),
    .B1(_0365_),
    .B2(\RAM[28][1] ),
    .C1(_0050_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0051_));
 sky130_fd_sc_hd__a22o_1 _0819_ (.A1(\RAM[18][1] ),
    .A2(_0340_),
    .B1(_0293_),
    .B2(\RAM[21][1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0052_));
 sky130_fd_sc_hd__a22o_1 _0820_ (.A1(\RAM[25][1] ),
    .A2(_0304_),
    .B1(_0296_),
    .B2(\RAM[29][1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0053_));
 sky130_fd_sc_hd__a22o_1 _0821_ (.A1(\RAM[23][1] ),
    .A2(_0285_),
    .B1(_0254_),
    .B2(\RAM[19][1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0054_));
 sky130_fd_sc_hd__a22o_1 _0822_ (.A1(\RAM[22][1] ),
    .A2(_0294_),
    .B1(_0327_),
    .B2(\RAM[16][1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0055_));
 sky130_fd_sc_hd__or4_2 _0823_ (.A(_0052_),
    .B(_0053_),
    .C(_0054_),
    .D(_0055_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0056_));
 sky130_fd_sc_hd__or3_1 _0824_ (.A(_0049_),
    .B(_0051_),
    .C(_0056_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0057_));
 sky130_fd_sc_hd__clkbuf_1 _0825_ (.A(_0057_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk2[1].selected_out[1] ));
 sky130_fd_sc_hd__a22o_1 _0826_ (.A1(\RAM[17][2] ),
    .A2(_0301_),
    .B1(_0370_),
    .B2(\RAM[20][2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0058_));
 sky130_fd_sc_hd__a221o_1 _0827_ (.A1(\RAM[21][2] ),
    .A2(_0248_),
    .B1(_0320_),
    .B2(\RAM[24][2] ),
    .C1(_0058_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0059_));
 sky130_fd_sc_hd__a22o_1 _0828_ (.A1(\RAM[28][2] ),
    .A2(_0286_),
    .B1(_0282_),
    .B2(\RAM[26][2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0060_));
 sky130_fd_sc_hd__a221o_1 _0829_ (.A1(\RAM[30][2] ),
    .A2(_0273_),
    .B1(_0267_),
    .B2(\RAM[25][2] ),
    .C1(_0060_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0061_));
 sky130_fd_sc_hd__a22o_1 _0830_ (.A1(\RAM[18][2] ),
    .A2(_0340_),
    .B1(_0294_),
    .B2(\RAM[22][2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0062_));
 sky130_fd_sc_hd__a221o_1 _0831_ (.A1(\RAM[27][2] ),
    .A2(_0260_),
    .B1(_0296_),
    .B2(\RAM[29][2] ),
    .C1(_0062_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0063_));
 sky130_fd_sc_hd__a22o_1 _0832_ (.A1(\RAM[23][2] ),
    .A2(_0285_),
    .B1(_0253_),
    .B2(\RAM[19][2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0064_));
 sky130_fd_sc_hd__a221o_1 _0833_ (.A1(\RAM[31][2] ),
    .A2(_0257_),
    .B1(_0327_),
    .B2(\RAM[16][2] ),
    .C1(_0064_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0065_));
 sky130_fd_sc_hd__or3_1 _0834_ (.A(_0061_),
    .B(_0063_),
    .C(_0065_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0066_));
 sky130_fd_sc_hd__or2_1 _0835_ (.A(_0059_),
    .B(_0066_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0067_));
 sky130_fd_sc_hd__clkbuf_1 _0836_ (.A(_0067_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk2[1].selected_out[2] ));
 sky130_fd_sc_hd__a22o_1 _0837_ (.A1(\RAM[30][3] ),
    .A2(_0346_),
    .B1(_0275_),
    .B2(\RAM[29][3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0068_));
 sky130_fd_sc_hd__a221o_1 _0838_ (.A1(\RAM[21][3] ),
    .A2(_0248_),
    .B1(_0303_),
    .B2(\RAM[16][3] ),
    .C1(_0068_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0069_));
 sky130_fd_sc_hd__a22o_1 _0839_ (.A1(\RAM[25][3] ),
    .A2(_0266_),
    .B1(_0286_),
    .B2(\RAM[28][3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0070_));
 sky130_fd_sc_hd__a221o_1 _0840_ (.A1(\RAM[24][3] ),
    .A2(_0281_),
    .B1(_0283_),
    .B2(\RAM[26][3] ),
    .C1(_0070_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0071_));
 sky130_fd_sc_hd__a22o_1 _0841_ (.A1(\RAM[18][3] ),
    .A2(net27),
    .B1(_0276_),
    .B2(\RAM[22][3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0072_));
 sky130_fd_sc_hd__a221o_1 _0842_ (.A1(\RAM[27][3] ),
    .A2(_0260_),
    .B1(_0353_),
    .B2(\RAM[17][3] ),
    .C1(_0072_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0073_));
 sky130_fd_sc_hd__a22o_1 _0843_ (.A1(\RAM[31][3] ),
    .A2(_0256_),
    .B1(_0285_),
    .B2(\RAM[23][3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0074_));
 sky130_fd_sc_hd__a221o_1 _0844_ (.A1(\RAM[19][3] ),
    .A2(_0339_),
    .B1(_0370_),
    .B2(\RAM[20][3] ),
    .C1(_0074_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0075_));
 sky130_fd_sc_hd__or3_1 _0845_ (.A(_0071_),
    .B(_0073_),
    .C(_0075_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0076_));
 sky130_fd_sc_hd__or2_1 _0846_ (.A(_0069_),
    .B(_0076_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0077_));
 sky130_fd_sc_hd__clkbuf_1 _0847_ (.A(_0077_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk2[1].selected_out[3] ));
 sky130_fd_sc_hd__a22o_1 _0848_ (.A1(\RAM[19][4] ),
    .A2(_0339_),
    .B1(_0275_),
    .B2(\RAM[29][4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0078_));
 sky130_fd_sc_hd__a221o_1 _0849_ (.A1(\RAM[30][4] ),
    .A2(_0421_),
    .B1(_0302_),
    .B2(\RAM[16][4] ),
    .C1(_0078_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0079_));
 sky130_fd_sc_hd__a22o_1 _0850_ (.A1(\RAM[31][4] ),
    .A2(_0258_),
    .B1(_0353_),
    .B2(\RAM[17][4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0080_));
 sky130_fd_sc_hd__a221o_1 _0851_ (.A1(\RAM[22][4] ),
    .A2(_0417_),
    .B1(_0320_),
    .B2(\RAM[24][4] ),
    .C1(_0080_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0081_));
 sky130_fd_sc_hd__a22o_1 _0852_ (.A1(\RAM[27][4] ),
    .A2(_0260_),
    .B1(_0304_),
    .B2(\RAM[25][4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0082_));
 sky130_fd_sc_hd__a22o_1 _0853_ (.A1(\RAM[18][4] ),
    .A2(_0340_),
    .B1(_0293_),
    .B2(\RAM[21][4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0083_));
 sky130_fd_sc_hd__a22o_1 _0854_ (.A1(\RAM[23][4] ),
    .A2(_0285_),
    .B1(_0265_),
    .B2(\RAM[20][4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0084_));
 sky130_fd_sc_hd__a22o_1 _0855_ (.A1(\RAM[28][4] ),
    .A2(_0287_),
    .B1(_0283_),
    .B2(\RAM[26][4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0085_));
 sky130_fd_sc_hd__or4_1 _0856_ (.A(_0082_),
    .B(_0083_),
    .C(_0084_),
    .D(_0085_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0086_));
 sky130_fd_sc_hd__or3_1 _0857_ (.A(_0079_),
    .B(_0081_),
    .C(_0086_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0087_));
 sky130_fd_sc_hd__clkbuf_1 _0858_ (.A(_0087_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk2[1].selected_out[4] ));
 sky130_fd_sc_hd__a22o_1 _0859_ (.A1(\RAM[31][5] ),
    .A2(_0258_),
    .B1(_0339_),
    .B2(\RAM[19][5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0088_));
 sky130_fd_sc_hd__a221o_1 _0860_ (.A1(\RAM[30][5] ),
    .A2(_0421_),
    .B1(_0391_),
    .B2(\RAM[26][5] ),
    .C1(_0088_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0089_));
 sky130_fd_sc_hd__a22o_1 _0861_ (.A1(\RAM[24][5] ),
    .A2(net25),
    .B1(_0286_),
    .B2(\RAM[28][5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0090_));
 sky130_fd_sc_hd__a221o_1 _0862_ (.A1(\RAM[23][5] ),
    .A2(_0322_),
    .B1(_0353_),
    .B2(\RAM[17][5] ),
    .C1(_0090_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0091_));
 sky130_fd_sc_hd__a22o_1 _0863_ (.A1(\RAM[18][5] ),
    .A2(net27),
    .B1(_0293_),
    .B2(\RAM[21][5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0092_));
 sky130_fd_sc_hd__a221o_1 _0864_ (.A1(\RAM[16][5] ),
    .A2(_0327_),
    .B1(_0267_),
    .B2(\RAM[25][5] ),
    .C1(_0092_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0093_));
 sky130_fd_sc_hd__a22o_1 _0865_ (.A1(\RAM[22][5] ),
    .A2(_0276_),
    .B1(_0274_),
    .B2(\RAM[29][5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0094_));
 sky130_fd_sc_hd__a221o_1 _0866_ (.A1(\RAM[27][5] ),
    .A2(_0260_),
    .B1(_0370_),
    .B2(\RAM[20][5] ),
    .C1(_0094_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0095_));
 sky130_fd_sc_hd__or3_1 _0867_ (.A(_0091_),
    .B(_0093_),
    .C(_0095_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0096_));
 sky130_fd_sc_hd__or2_1 _0868_ (.A(_0089_),
    .B(_0096_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0097_));
 sky130_fd_sc_hd__clkbuf_1 _0869_ (.A(_0097_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk2[1].selected_out[5] ));
 sky130_fd_sc_hd__a22o_1 _0870_ (.A1(\RAM[27][6] ),
    .A2(_0261_),
    .B1(_0346_),
    .B2(\RAM[30][6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0098_));
 sky130_fd_sc_hd__a221o_1 _0871_ (.A1(\RAM[31][6] ),
    .A2(_0345_),
    .B1(_0369_),
    .B2(\RAM[23][6] ),
    .C1(_0098_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0099_));
 sky130_fd_sc_hd__a22o_1 _0872_ (.A1(\RAM[17][6] ),
    .A2(_0353_),
    .B1(_0267_),
    .B2(\RAM[25][6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0100_));
 sky130_fd_sc_hd__a221o_1 _0873_ (.A1(\RAM[16][6] ),
    .A2(_0302_),
    .B1(_0391_),
    .B2(\RAM[26][6] ),
    .C1(_0100_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0101_));
 sky130_fd_sc_hd__a22o_1 _0874_ (.A1(\RAM[22][6] ),
    .A2(_0294_),
    .B1(_0296_),
    .B2(\RAM[29][6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0102_));
 sky130_fd_sc_hd__a22o_1 _0875_ (.A1(\RAM[20][6] ),
    .A2(net28),
    .B1(_0281_),
    .B2(\RAM[24][6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0103_));
 sky130_fd_sc_hd__a22o_1 _0876_ (.A1(\RAM[21][6] ),
    .A2(_0293_),
    .B1(_0287_),
    .B2(\RAM[28][6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0104_));
 sky130_fd_sc_hd__a22o_1 _0877_ (.A1(\RAM[18][6] ),
    .A2(_0340_),
    .B1(_0254_),
    .B2(\RAM[19][6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0105_));
 sky130_fd_sc_hd__or4_1 _0878_ (.A(_0102_),
    .B(_0103_),
    .C(_0104_),
    .D(_0105_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0106_));
 sky130_fd_sc_hd__or3_1 _0879_ (.A(_0099_),
    .B(_0101_),
    .C(_0106_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0107_));
 sky130_fd_sc_hd__clkbuf_1 _0880_ (.A(_0107_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk2[1].selected_out[6] ));
 sky130_fd_sc_hd__a22o_1 _0881_ (.A1(\RAM[31][7] ),
    .A2(_0258_),
    .B1(_0247_),
    .B2(\RAM[21][7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0108_));
 sky130_fd_sc_hd__a221o_1 _0882_ (.A1(\RAM[23][7] ),
    .A2(_0369_),
    .B1(_0421_),
    .B2(\RAM[30][7] ),
    .C1(_0108_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0109_));
 sky130_fd_sc_hd__a22o_1 _0883_ (.A1(\RAM[22][7] ),
    .A2(_0334_),
    .B1(_0275_),
    .B2(\RAM[29][7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0110_));
 sky130_fd_sc_hd__a221o_1 _0884_ (.A1(\RAM[18][7] ),
    .A2(_0309_),
    .B1(_0302_),
    .B2(\RAM[16][7] ),
    .C1(_0110_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0111_));
 sky130_fd_sc_hd__a22o_1 _0885_ (.A1(\RAM[19][7] ),
    .A2(_0254_),
    .B1(_0304_),
    .B2(\RAM[25][7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0112_));
 sky130_fd_sc_hd__a22o_1 _0886_ (.A1(\RAM[20][7] ),
    .A2(net28),
    .B1(_0283_),
    .B2(\RAM[26][7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0113_));
 sky130_fd_sc_hd__a22o_1 _0887_ (.A1(\RAM[27][7] ),
    .A2(_0260_),
    .B1(_0281_),
    .B2(\RAM[24][7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0114_));
 sky130_fd_sc_hd__a22o_1 _0888_ (.A1(\RAM[17][7] ),
    .A2(_0300_),
    .B1(_0316_),
    .B2(\RAM[28][7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0115_));
 sky130_fd_sc_hd__or4_1 _0889_ (.A(_0112_),
    .B(_0113_),
    .C(_0114_),
    .D(_0115_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0116_));
 sky130_fd_sc_hd__or3_1 _0890_ (.A(_0109_),
    .B(_0111_),
    .C(_0116_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0117_));
 sky130_fd_sc_hd__clkbuf_1 _0891_ (.A(_0117_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk2[1].selected_out[7] ));
 sky130_fd_sc_hd__or4_2 _0892_ (.A(_0249_),
    .B(_0250_),
    .C(_0251_),
    .D(_0252_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0118_));
 sky130_fd_sc_hd__buf_2 _0893_ (.A(_0118_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0119_));
 sky130_fd_sc_hd__a22o_1 _0894_ (.A1(\RAM[1][0] ),
    .A2(_0300_),
    .B1(_0267_),
    .B2(\RAM[9][0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0120_));
 sky130_fd_sc_hd__a221o_1 _0895_ (.A1(\RAM[11][0] ),
    .A2(_0315_),
    .B1(_0365_),
    .B2(\RAM[12][0] ),
    .C1(_0120_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0121_));
 sky130_fd_sc_hd__a22o_1 _0896_ (.A1(\RAM[7][0] ),
    .A2(_0369_),
    .B1(_0310_),
    .B2(\RAM[4][0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0122_));
 sky130_fd_sc_hd__a2111o_1 _0897_ (.A1(\RAM[13][0] ),
    .A2(_0321_),
    .B1(_0121_),
    .C1(_0122_),
    .D1(_0303_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0123_));
 sky130_fd_sc_hd__a22o_1 _0898_ (.A1(\RAM[5][0] ),
    .A2(_0247_),
    .B1(_0311_),
    .B2(\RAM[10][0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0124_));
 sky130_fd_sc_hd__a22o_1 _0899_ (.A1(\RAM[2][0] ),
    .A2(_0309_),
    .B1(_0255_),
    .B2(\RAM[3][0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0125_));
 sky130_fd_sc_hd__a22o_1 _0900_ (.A1(\RAM[14][0] ),
    .A2(_0421_),
    .B1(_0319_),
    .B2(\RAM[8][0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0126_));
 sky130_fd_sc_hd__a22o_1 _0901_ (.A1(\RAM[15][0] ),
    .A2(_0345_),
    .B1(_0417_),
    .B2(\RAM[6][0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0127_));
 sky130_fd_sc_hd__or4_1 _0902_ (.A(_0124_),
    .B(_0125_),
    .C(_0126_),
    .D(_0127_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0128_));
 sky130_fd_sc_hd__o22a_1 _0903_ (.A1(\RAM[0][0] ),
    .A2(_0119_),
    .B1(_0123_),
    .B2(_0128_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk2[0].selected_out[0] ));
 sky130_fd_sc_hd__a22o_1 _0904_ (.A1(\RAM[6][1] ),
    .A2(_0417_),
    .B1(_0421_),
    .B2(\RAM[14][1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0129_));
 sky130_fd_sc_hd__a22o_1 _0905_ (.A1(\RAM[11][1] ),
    .A2(_0261_),
    .B1(_0311_),
    .B2(\RAM[10][1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0130_));
 sky130_fd_sc_hd__a221o_1 _0906_ (.A1(\RAM[5][1] ),
    .A2(_0248_),
    .B1(_0320_),
    .B2(\RAM[8][1] ),
    .C1(_0130_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0131_));
 sky130_fd_sc_hd__a2111o_1 _0907_ (.A1(\RAM[15][1] ),
    .A2(_0345_),
    .B1(_0303_),
    .C1(_0129_),
    .D1(_0131_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0132_));
 sky130_fd_sc_hd__a22o_1 _0908_ (.A1(\RAM[4][1] ),
    .A2(_0370_),
    .B1(_0305_),
    .B2(\RAM[9][1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0133_));
 sky130_fd_sc_hd__a22o_1 _0909_ (.A1(\RAM[3][1] ),
    .A2(_0255_),
    .B1(_0301_),
    .B2(\RAM[1][1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0134_));
 sky130_fd_sc_hd__a22o_1 _0910_ (.A1(\RAM[13][1] ),
    .A2(_0321_),
    .B1(_0365_),
    .B2(\RAM[12][1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0135_));
 sky130_fd_sc_hd__a22o_1 _0911_ (.A1(\RAM[2][1] ),
    .A2(_0309_),
    .B1(_0369_),
    .B2(\RAM[7][1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0136_));
 sky130_fd_sc_hd__or4_1 _0912_ (.A(_0133_),
    .B(_0134_),
    .C(_0135_),
    .D(_0136_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0137_));
 sky130_fd_sc_hd__o22a_1 _0913_ (.A1(\RAM[0][1] ),
    .A2(_0119_),
    .B1(_0132_),
    .B2(_0137_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk2[0].selected_out[1] ));
 sky130_fd_sc_hd__a22o_1 _0914_ (.A1(\RAM[15][2] ),
    .A2(_0257_),
    .B1(_0334_),
    .B2(\RAM[6][2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0138_));
 sky130_fd_sc_hd__a221o_1 _0915_ (.A1(\RAM[5][2] ),
    .A2(_0248_),
    .B1(_0301_),
    .B2(\RAM[1][2] ),
    .C1(_0138_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0139_));
 sky130_fd_sc_hd__a22o_1 _0916_ (.A1(\RAM[3][2] ),
    .A2(_0255_),
    .B1(_0320_),
    .B2(\RAM[8][2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0140_));
 sky130_fd_sc_hd__a2111o_1 _0917_ (.A1(\RAM[14][2] ),
    .A2(_0421_),
    .B1(_0303_),
    .C1(_0139_),
    .D1(_0140_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0141_));
 sky130_fd_sc_hd__a22o_1 _0918_ (.A1(\RAM[13][2] ),
    .A2(_0275_),
    .B1(_0316_),
    .B2(\RAM[12][2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0142_));
 sky130_fd_sc_hd__a22o_1 _0919_ (.A1(\RAM[2][2] ),
    .A2(_0309_),
    .B1(_0322_),
    .B2(\RAM[7][2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0143_));
 sky130_fd_sc_hd__a22o_1 _0920_ (.A1(\RAM[4][2] ),
    .A2(_0370_),
    .B1(_0305_),
    .B2(\RAM[9][2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0144_));
 sky130_fd_sc_hd__a22o_1 _0921_ (.A1(\RAM[11][2] ),
    .A2(_0315_),
    .B1(_0391_),
    .B2(\RAM[10][2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0145_));
 sky130_fd_sc_hd__or4_1 _0922_ (.A(_0142_),
    .B(_0143_),
    .C(_0144_),
    .D(_0145_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0146_));
 sky130_fd_sc_hd__o22a_1 _0923_ (.A1(\RAM[0][2] ),
    .A2(_0119_),
    .B1(_0141_),
    .B2(_0146_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk2[0].selected_out[2] ));
 sky130_fd_sc_hd__a22o_1 _0924_ (.A1(\RAM[1][3] ),
    .A2(_0300_),
    .B1(_0267_),
    .B2(\RAM[9][3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0147_));
 sky130_fd_sc_hd__a221o_1 _0925_ (.A1(\RAM[12][3] ),
    .A2(_0365_),
    .B1(_0391_),
    .B2(\RAM[10][3] ),
    .C1(_0147_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0148_));
 sky130_fd_sc_hd__a22o_1 _0926_ (.A1(\RAM[7][3] ),
    .A2(_0369_),
    .B1(_0310_),
    .B2(\RAM[4][3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0149_));
 sky130_fd_sc_hd__a2111o_1 _0927_ (.A1(\RAM[13][3] ),
    .A2(_0321_),
    .B1(_0148_),
    .C1(_0149_),
    .D1(_0303_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0150_));
 sky130_fd_sc_hd__a22o_1 _0928_ (.A1(\RAM[5][3] ),
    .A2(_0247_),
    .B1(_0261_),
    .B2(\RAM[11][3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0151_));
 sky130_fd_sc_hd__a22o_1 _0929_ (.A1(\RAM[2][3] ),
    .A2(_0309_),
    .B1(_0255_),
    .B2(\RAM[3][3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0152_));
 sky130_fd_sc_hd__a22o_1 _0930_ (.A1(\RAM[14][3] ),
    .A2(_0346_),
    .B1(_0319_),
    .B2(\RAM[8][3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0153_));
 sky130_fd_sc_hd__a22o_1 _0931_ (.A1(\RAM[15][3] ),
    .A2(_0345_),
    .B1(_0417_),
    .B2(\RAM[6][3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0154_));
 sky130_fd_sc_hd__or4_1 _0932_ (.A(_0151_),
    .B(_0152_),
    .C(_0153_),
    .D(_0154_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0155_));
 sky130_fd_sc_hd__o22a_1 _0933_ (.A1(\RAM[0][3] ),
    .A2(_0119_),
    .B1(_0150_),
    .B2(_0155_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk2[0].selected_out[3] ));
 sky130_fd_sc_hd__a22o_1 _0934_ (.A1(\RAM[1][4] ),
    .A2(_0300_),
    .B1(_0267_),
    .B2(\RAM[9][4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0156_));
 sky130_fd_sc_hd__a221o_1 _0935_ (.A1(\RAM[11][4] ),
    .A2(_0261_),
    .B1(_0365_),
    .B2(\RAM[12][4] ),
    .C1(_0156_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0157_));
 sky130_fd_sc_hd__a22o_1 _0936_ (.A1(\RAM[7][4] ),
    .A2(_0369_),
    .B1(_0310_),
    .B2(\RAM[4][4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0158_));
 sky130_fd_sc_hd__a2111o_1 _0937_ (.A1(\RAM[13][4] ),
    .A2(_0321_),
    .B1(_0157_),
    .C1(_0158_),
    .D1(_0303_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0159_));
 sky130_fd_sc_hd__a22o_1 _0938_ (.A1(\RAM[5][4] ),
    .A2(_0247_),
    .B1(_0311_),
    .B2(\RAM[10][4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0160_));
 sky130_fd_sc_hd__a22o_1 _0939_ (.A1(\RAM[2][4] ),
    .A2(_0309_),
    .B1(_0255_),
    .B2(\RAM[3][4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0161_));
 sky130_fd_sc_hd__a22o_1 _0940_ (.A1(\RAM[14][4] ),
    .A2(_0346_),
    .B1(_0319_),
    .B2(\RAM[8][4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0162_));
 sky130_fd_sc_hd__a22o_1 _0941_ (.A1(\RAM[15][4] ),
    .A2(_0345_),
    .B1(_0417_),
    .B2(\RAM[6][4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0163_));
 sky130_fd_sc_hd__or4_1 _0942_ (.A(_0160_),
    .B(_0161_),
    .C(_0162_),
    .D(_0163_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0164_));
 sky130_fd_sc_hd__o22a_1 _0943_ (.A1(\RAM[0][4] ),
    .A2(_0119_),
    .B1(_0159_),
    .B2(_0164_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk2[0].selected_out[4] ));
 sky130_fd_sc_hd__a22o_1 _0944_ (.A1(\RAM[6][5] ),
    .A2(_0417_),
    .B1(_0421_),
    .B2(\RAM[14][5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0165_));
 sky130_fd_sc_hd__a22o_1 _0945_ (.A1(\RAM[11][5] ),
    .A2(_0261_),
    .B1(_0311_),
    .B2(\RAM[10][5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0166_));
 sky130_fd_sc_hd__a221o_1 _0946_ (.A1(\RAM[5][5] ),
    .A2(_0248_),
    .B1(_0319_),
    .B2(\RAM[8][5] ),
    .C1(_0166_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0167_));
 sky130_fd_sc_hd__a2111o_1 _0947_ (.A1(\RAM[15][5] ),
    .A2(_0345_),
    .B1(_0303_),
    .C1(_0165_),
    .D1(_0167_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0168_));
 sky130_fd_sc_hd__a22o_1 _0948_ (.A1(\RAM[4][5] ),
    .A2(_0370_),
    .B1(_0305_),
    .B2(\RAM[9][5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0169_));
 sky130_fd_sc_hd__a22o_1 _0949_ (.A1(\RAM[3][5] ),
    .A2(_0339_),
    .B1(_0301_),
    .B2(\RAM[1][5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0170_));
 sky130_fd_sc_hd__a22o_1 _0950_ (.A1(\RAM[13][5] ),
    .A2(_0275_),
    .B1(_0365_),
    .B2(\RAM[12][5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0171_));
 sky130_fd_sc_hd__a22o_1 _0951_ (.A1(\RAM[2][5] ),
    .A2(_0309_),
    .B1(_0369_),
    .B2(\RAM[7][5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0172_));
 sky130_fd_sc_hd__or4_1 _0952_ (.A(_0169_),
    .B(_0170_),
    .C(_0171_),
    .D(_0172_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0173_));
 sky130_fd_sc_hd__o22a_1 _0953_ (.A1(\RAM[0][5] ),
    .A2(_0119_),
    .B1(_0168_),
    .B2(_0173_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk2[0].selected_out[5] ));
 sky130_fd_sc_hd__a22o_1 _0954_ (.A1(\RAM[9][6] ),
    .A2(_0304_),
    .B1(_0316_),
    .B2(\RAM[12][6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0174_));
 sky130_fd_sc_hd__a221o_1 _0955_ (.A1(\RAM[11][6] ),
    .A2(_0261_),
    .B1(_0301_),
    .B2(\RAM[1][6] ),
    .C1(_0174_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0175_));
 sky130_fd_sc_hd__a22o_1 _0956_ (.A1(\RAM[7][6] ),
    .A2(_0369_),
    .B1(_0310_),
    .B2(\RAM[4][6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0176_));
 sky130_fd_sc_hd__a2111o_1 _0957_ (.A1(\RAM[13][6] ),
    .A2(_0321_),
    .B1(_0175_),
    .C1(_0176_),
    .D1(_0303_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0177_));
 sky130_fd_sc_hd__a22o_1 _0958_ (.A1(\RAM[5][6] ),
    .A2(_0247_),
    .B1(_0311_),
    .B2(\RAM[10][6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0178_));
 sky130_fd_sc_hd__a22o_1 _0959_ (.A1(\RAM[2][6] ),
    .A2(_0309_),
    .B1(_0255_),
    .B2(\RAM[3][6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0179_));
 sky130_fd_sc_hd__a22o_1 _0960_ (.A1(\RAM[14][6] ),
    .A2(_0346_),
    .B1(_0319_),
    .B2(\RAM[8][6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0180_));
 sky130_fd_sc_hd__a22o_1 _0961_ (.A1(\RAM[15][6] ),
    .A2(_0258_),
    .B1(_0417_),
    .B2(\RAM[6][6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0181_));
 sky130_fd_sc_hd__or4_1 _0962_ (.A(_0178_),
    .B(_0179_),
    .C(_0180_),
    .D(_0181_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0182_));
 sky130_fd_sc_hd__o22a_1 _0963_ (.A1(\RAM[0][6] ),
    .A2(_0119_),
    .B1(_0177_),
    .B2(_0182_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk2[0].selected_out[6] ));
 sky130_fd_sc_hd__a22o_1 _0964_ (.A1(\RAM[6][7] ),
    .A2(_0417_),
    .B1(_0421_),
    .B2(\RAM[14][7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0183_));
 sky130_fd_sc_hd__a22o_1 _0965_ (.A1(\RAM[11][7] ),
    .A2(_0260_),
    .B1(_0283_),
    .B2(\RAM[10][7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0184_));
 sky130_fd_sc_hd__a221o_1 _0966_ (.A1(\RAM[5][7] ),
    .A2(_0248_),
    .B1(_0319_),
    .B2(\RAM[8][7] ),
    .C1(_0184_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0185_));
 sky130_fd_sc_hd__a2111o_1 _0967_ (.A1(\RAM[15][7] ),
    .A2(_0345_),
    .B1(_0303_),
    .C1(_0183_),
    .D1(_0185_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0186_));
 sky130_fd_sc_hd__a22o_1 _0968_ (.A1(\RAM[13][7] ),
    .A2(_0275_),
    .B1(_0316_),
    .B2(\RAM[12][7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0187_));
 sky130_fd_sc_hd__a221o_1 _0969_ (.A1(\RAM[3][7] ),
    .A2(_0255_),
    .B1(_0301_),
    .B2(\RAM[1][7] ),
    .C1(_0187_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0188_));
 sky130_fd_sc_hd__a22o_1 _0970_ (.A1(\RAM[2][7] ),
    .A2(_0308_),
    .B1(_0322_),
    .B2(\RAM[7][7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0189_));
 sky130_fd_sc_hd__a221o_1 _0971_ (.A1(\RAM[4][7] ),
    .A2(_0310_),
    .B1(_0305_),
    .B2(\RAM[9][7] ),
    .C1(_0189_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0190_));
 sky130_fd_sc_hd__or2_1 _0972_ (.A(_0188_),
    .B(_0190_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0191_));
 sky130_fd_sc_hd__o22a_1 _0973_ (.A1(\RAM[0][7] ),
    .A2(_0119_),
    .B1(_0186_),
    .B2(_0191_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk2[0].selected_out[7] ));
 sky130_fd_sc_hd__nor2b_2 _0974_ (.A(wr_en_next),
    .B_N(net8),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0192_));
 sky130_fd_sc_hd__clkbuf_4 _0975_ (.A(_0192_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0193_));
 sky130_fd_sc_hd__mux2_1 _0976_ (.A0(net95),
    .A1(net9),
    .S(_0193_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0194_));
 sky130_fd_sc_hd__clkbuf_1 _0977_ (.A(_0194_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0006_));
 sky130_fd_sc_hd__mux2_1 _0978_ (.A0(net87),
    .A1(net10),
    .S(_0193_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0195_));
 sky130_fd_sc_hd__clkbuf_1 _0979_ (.A(_0195_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0007_));
 sky130_fd_sc_hd__mux2_1 _0980_ (.A0(net78),
    .A1(net11),
    .S(_0193_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0196_));
 sky130_fd_sc_hd__clkbuf_1 _0981_ (.A(_0196_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0008_));
 sky130_fd_sc_hd__mux2_1 _0982_ (.A0(net69),
    .A1(net12),
    .S(_0193_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0197_));
 sky130_fd_sc_hd__clkbuf_1 _0983_ (.A(_0197_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0009_));
 sky130_fd_sc_hd__mux2_1 _0984_ (.A0(net62),
    .A1(net13),
    .S(_0193_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0198_));
 sky130_fd_sc_hd__clkbuf_1 _0985_ (.A(_0198_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0010_));
 sky130_fd_sc_hd__mux2_1 _0986_ (.A0(net54),
    .A1(net14),
    .S(_0193_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0199_));
 sky130_fd_sc_hd__clkbuf_1 _0987_ (.A(_0199_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0011_));
 sky130_fd_sc_hd__mux2_1 _0988_ (.A0(net46),
    .A1(net15),
    .S(_0193_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0200_));
 sky130_fd_sc_hd__clkbuf_1 _0989_ (.A(_0200_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0012_));
 sky130_fd_sc_hd__mux2_1 _0990_ (.A0(net36),
    .A1(net16),
    .S(_0193_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0201_));
 sky130_fd_sc_hd__clkbuf_1 _0991_ (.A(_0201_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0013_));
 sky130_fd_sc_hd__inv_2 _0992__1 (.A(clknet_1_1__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net112));
 sky130_fd_sc_hd__mux2_1 _0993_ (.A0(_0217_),
    .A1(net2),
    .S(_0193_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0202_));
 sky130_fd_sc_hd__clkbuf_1 _0994_ (.A(_0202_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0014_));
 sky130_fd_sc_hd__mux2_1 _0995_ (.A0(_0219_),
    .A1(net3),
    .S(_0192_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0203_));
 sky130_fd_sc_hd__clkbuf_1 _0996_ (.A(_0203_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0015_));
 sky130_fd_sc_hd__mux2_1 _0997_ (.A0(_0221_),
    .A1(net4),
    .S(_0192_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0204_));
 sky130_fd_sc_hd__clkbuf_1 _0998_ (.A(_0204_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0016_));
 sky130_fd_sc_hd__mux2_1 _0999_ (.A0(_0222_),
    .A1(net5),
    .S(_0192_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0205_));
 sky130_fd_sc_hd__clkbuf_1 _1000_ (.A(_0205_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0017_));
 sky130_fd_sc_hd__mux2_1 _1001_ (.A0(\addr_write[4] ),
    .A1(net6),
    .S(_0192_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0206_));
 sky130_fd_sc_hd__clkbuf_1 _1002_ (.A(_0206_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0018_));
 sky130_fd_sc_hd__mux2_1 _1003_ (.A0(\addr_write[5] ),
    .A1(net7),
    .S(_0192_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0207_));
 sky130_fd_sc_hd__clkbuf_1 _1004_ (.A(_0207_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0019_));
 sky130_fd_sc_hd__and2_1 _1005_ (.A(net1),
    .B(_0193_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0208_));
 sky130_fd_sc_hd__clkbuf_1 _1006_ (.A(_0208_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0020_));
 sky130_fd_sc_hd__and2_1 _1007_ (.A(net113),
    .B(net1),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0209_));
 sky130_fd_sc_hd__clkbuf_1 _1008_ (.A(_0209_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0021_));
 sky130_fd_sc_hd__dfxtp_1 _1009_ (.CLK(clknet_1_1__leaf_clk),
    .D(_0006_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\data_to_write[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1010_ (.CLK(clknet_1_0__leaf_clk),
    .D(_0007_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\data_to_write[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1011_ (.CLK(clknet_1_1__leaf_clk),
    .D(_0008_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\data_to_write[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1012_ (.CLK(clknet_1_0__leaf_clk),
    .D(_0009_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\data_to_write[3] ));
 sky130_fd_sc_hd__dfxtp_2 _1013_ (.CLK(clknet_1_0__leaf_clk),
    .D(_0010_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\data_to_write[4] ));
 sky130_fd_sc_hd__dfxtp_1 _1014_ (.CLK(clknet_1_0__leaf_clk),
    .D(_0011_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\data_to_write[5] ));
 sky130_fd_sc_hd__dfxtp_1 _1015_ (.CLK(clknet_1_0__leaf_clk),
    .D(_0012_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\data_to_write[6] ));
 sky130_fd_sc_hd__dfxtp_1 _1016_ (.CLK(clknet_1_0__leaf_clk),
    .D(_0013_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\data_to_write[7] ));
 sky130_fd_sc_hd__dlxtp_1 _1017_ (.D(net93),
    .GATE(\genblk1[63].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[63][0] ));
 sky130_fd_sc_hd__dlxtp_1 _1018_ (.D(net85),
    .GATE(\genblk1[63].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[63][1] ));
 sky130_fd_sc_hd__dlxtp_1 _1019_ (.D(net77),
    .GATE(\genblk1[63].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[63][2] ));
 sky130_fd_sc_hd__dlxtp_1 _1020_ (.D(net69),
    .GATE(\genblk1[63].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[63][3] ));
 sky130_fd_sc_hd__dlxtp_1 _1021_ (.D(net62),
    .GATE(\genblk1[63].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[63][4] ));
 sky130_fd_sc_hd__dlxtp_1 _1022_ (.D(net52),
    .GATE(\genblk1[63].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[63][5] ));
 sky130_fd_sc_hd__dlxtp_1 _1023_ (.D(net44),
    .GATE(\genblk1[63].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[63][6] ));
 sky130_fd_sc_hd__dlxtp_1 _1024_ (.D(net36),
    .GATE(\genblk1[63].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[63][7] ));
 sky130_fd_sc_hd__dlxtp_1 _1025_ (.D(net93),
    .GATE(\genblk1[62].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[62][0] ));
 sky130_fd_sc_hd__dlxtp_1 _1026_ (.D(net87),
    .GATE(\genblk1[62].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[62][1] ));
 sky130_fd_sc_hd__dlxtp_1 _1027_ (.D(net78),
    .GATE(\genblk1[62].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[62][2] ));
 sky130_fd_sc_hd__dlxtp_1 _1028_ (.D(net69),
    .GATE(\genblk1[62].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[62][3] ));
 sky130_fd_sc_hd__dlxtp_1 _1029_ (.D(net62),
    .GATE(\genblk1[62].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[62][4] ));
 sky130_fd_sc_hd__dlxtp_1 _1030_ (.D(net54),
    .GATE(\genblk1[62].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[62][5] ));
 sky130_fd_sc_hd__dlxtp_1 _1031_ (.D(net44),
    .GATE(\genblk1[62].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[62][6] ));
 sky130_fd_sc_hd__dlxtp_1 _1032_ (.D(net34),
    .GATE(\genblk1[62].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[62][7] ));
 sky130_fd_sc_hd__dlxtp_1 _1033_ (.D(net93),
    .GATE(\genblk1[61].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[61][0] ));
 sky130_fd_sc_hd__dlxtp_1 _1034_ (.D(net87),
    .GATE(\genblk1[61].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[61][1] ));
 sky130_fd_sc_hd__dlxtp_1 _1035_ (.D(net77),
    .GATE(\genblk1[61].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[61][2] ));
 sky130_fd_sc_hd__dlxtp_1 _1036_ (.D(net68),
    .GATE(\genblk1[61].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[61][3] ));
 sky130_fd_sc_hd__dlxtp_1 _1037_ (.D(net60),
    .GATE(\genblk1[61].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[61][4] ));
 sky130_fd_sc_hd__dlxtp_1 _1038_ (.D(net52),
    .GATE(\genblk1[61].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[61][5] ));
 sky130_fd_sc_hd__dlxtp_1 _1039_ (.D(net45),
    .GATE(\genblk1[61].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[61][6] ));
 sky130_fd_sc_hd__dlxtp_1 _1040_ (.D(net34),
    .GATE(\genblk1[61].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[61][7] ));
 sky130_fd_sc_hd__dlxtp_1 _1041_ (.D(net93),
    .GATE(\genblk1[60].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[60][0] ));
 sky130_fd_sc_hd__dlxtp_1 _1042_ (.D(net85),
    .GATE(\genblk1[60].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[60][1] ));
 sky130_fd_sc_hd__dlxtp_1 _1043_ (.D(net78),
    .GATE(\genblk1[60].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[60][2] ));
 sky130_fd_sc_hd__dlxtp_1 _1044_ (.D(net68),
    .GATE(\genblk1[60].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[60][3] ));
 sky130_fd_sc_hd__dlxtp_1 _1045_ (.D(net62),
    .GATE(\genblk1[60].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[60][4] ));
 sky130_fd_sc_hd__dlxtp_1 _1046_ (.D(net52),
    .GATE(\genblk1[60].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[60][5] ));
 sky130_fd_sc_hd__dlxtp_1 _1047_ (.D(net44),
    .GATE(\genblk1[60].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[60][6] ));
 sky130_fd_sc_hd__dlxtp_1 _1048_ (.D(net34),
    .GATE(\genblk1[60].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[60][7] ));
 sky130_fd_sc_hd__dlxtp_1 _1049_ (.D(net94),
    .GATE(\genblk1[59].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[59][0] ));
 sky130_fd_sc_hd__dlxtp_1 _1050_ (.D(net85),
    .GATE(\genblk1[59].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[59][1] ));
 sky130_fd_sc_hd__dlxtp_1 _1051_ (.D(net77),
    .GATE(\genblk1[59].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[59][2] ));
 sky130_fd_sc_hd__dlxtp_1 _1052_ (.D(net69),
    .GATE(\genblk1[59].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[59][3] ));
 sky130_fd_sc_hd__dlxtp_1 _1053_ (.D(net60),
    .GATE(\genblk1[59].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[59][4] ));
 sky130_fd_sc_hd__dlxtp_1 _1054_ (.D(net54),
    .GATE(\genblk1[59].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[59][5] ));
 sky130_fd_sc_hd__dlxtp_1 _1055_ (.D(net45),
    .GATE(\genblk1[59].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[59][6] ));
 sky130_fd_sc_hd__dlxtp_1 _1056_ (.D(net34),
    .GATE(\genblk1[59].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[59][7] ));
 sky130_fd_sc_hd__dlxtp_1 _1057_ (.D(net95),
    .GATE(\genblk1[58].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[58][0] ));
 sky130_fd_sc_hd__dlxtp_1 _1058_ (.D(net87),
    .GATE(\genblk1[58].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[58][1] ));
 sky130_fd_sc_hd__dlxtp_1 _1059_ (.D(net77),
    .GATE(\genblk1[58].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[58][2] ));
 sky130_fd_sc_hd__dlxtp_1 _1060_ (.D(net69),
    .GATE(\genblk1[58].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[58][3] ));
 sky130_fd_sc_hd__dlxtp_1 _1061_ (.D(net62),
    .GATE(\genblk1[58].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[58][4] ));
 sky130_fd_sc_hd__dlxtp_1 _1062_ (.D(net52),
    .GATE(\genblk1[58].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[58][5] ));
 sky130_fd_sc_hd__dlxtp_1 _1063_ (.D(net45),
    .GATE(\genblk1[58].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[58][6] ));
 sky130_fd_sc_hd__dlxtp_1 _1064_ (.D(net34),
    .GATE(\genblk1[58].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[58][7] ));
 sky130_fd_sc_hd__dlxtp_1 _1065_ (.D(net95),
    .GATE(\genblk1[57].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[57][0] ));
 sky130_fd_sc_hd__dlxtp_1 _1066_ (.D(net85),
    .GATE(\genblk1[57].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[57][1] ));
 sky130_fd_sc_hd__dlxtp_1 _1067_ (.D(net77),
    .GATE(\genblk1[57].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[57][2] ));
 sky130_fd_sc_hd__dlxtp_1 _1068_ (.D(net69),
    .GATE(\genblk1[57].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[57][3] ));
 sky130_fd_sc_hd__dlxtp_1 _1069_ (.D(net62),
    .GATE(\genblk1[57].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[57][4] ));
 sky130_fd_sc_hd__dlxtp_1 _1070_ (.D(net52),
    .GATE(\genblk1[57].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[57][5] ));
 sky130_fd_sc_hd__dlxtp_1 _1071_ (.D(net44),
    .GATE(\genblk1[57].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[57][6] ));
 sky130_fd_sc_hd__dlxtp_1 _1072_ (.D(net34),
    .GATE(\genblk1[57].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[57][7] ));
 sky130_fd_sc_hd__dlxtp_1 _1073_ (.D(net95),
    .GATE(\genblk1[56].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[56][0] ));
 sky130_fd_sc_hd__dlxtp_1 _1074_ (.D(net85),
    .GATE(\genblk1[56].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[56][1] ));
 sky130_fd_sc_hd__dlxtp_1 _1075_ (.D(net77),
    .GATE(\genblk1[56].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[56][2] ));
 sky130_fd_sc_hd__dlxtp_1 _1076_ (.D(net69),
    .GATE(\genblk1[56].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[56][3] ));
 sky130_fd_sc_hd__dlxtp_1 _1077_ (.D(net59),
    .GATE(\genblk1[56].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[56][4] ));
 sky130_fd_sc_hd__dlxtp_1 _1078_ (.D(net53),
    .GATE(\genblk1[56].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[56][5] ));
 sky130_fd_sc_hd__dlxtp_1 _1079_ (.D(net45),
    .GATE(\genblk1[56].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[56][6] ));
 sky130_fd_sc_hd__dlxtp_1 _1080_ (.D(net36),
    .GATE(\genblk1[56].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[56][7] ));
 sky130_fd_sc_hd__dlxtp_1 _1081_ (.D(net93),
    .GATE(\genblk1[55].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[55][0] ));
 sky130_fd_sc_hd__dlxtp_1 _1082_ (.D(net85),
    .GATE(\genblk1[55].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[55][1] ));
 sky130_fd_sc_hd__dlxtp_1 _1083_ (.D(net78),
    .GATE(\genblk1[55].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[55][2] ));
 sky130_fd_sc_hd__dlxtp_1 _1084_ (.D(net69),
    .GATE(\genblk1[55].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[55][3] ));
 sky130_fd_sc_hd__dlxtp_1 _1085_ (.D(net59),
    .GATE(\genblk1[55].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[55][4] ));
 sky130_fd_sc_hd__dlxtp_1 _1086_ (.D(net52),
    .GATE(\genblk1[55].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[55][5] ));
 sky130_fd_sc_hd__dlxtp_1 _1087_ (.D(net45),
    .GATE(\genblk1[55].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[55][6] ));
 sky130_fd_sc_hd__dlxtp_1 _1088_ (.D(net34),
    .GATE(\genblk1[55].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[55][7] ));
 sky130_fd_sc_hd__dlxtp_1 _1089_ (.D(net95),
    .GATE(\genblk1[54].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[54][0] ));
 sky130_fd_sc_hd__dlxtp_1 _1090_ (.D(net86),
    .GATE(\genblk1[54].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[54][1] ));
 sky130_fd_sc_hd__dlxtp_1 _1091_ (.D(net78),
    .GATE(\genblk1[54].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[54][2] ));
 sky130_fd_sc_hd__dlxtp_1 _1092_ (.D(net70),
    .GATE(\genblk1[54].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[54][3] ));
 sky130_fd_sc_hd__dlxtp_1 _1093_ (.D(net62),
    .GATE(\genblk1[54].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[54][4] ));
 sky130_fd_sc_hd__dlxtp_1 _1094_ (.D(net54),
    .GATE(\genblk1[54].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[54][5] ));
 sky130_fd_sc_hd__dlxtp_1 _1095_ (.D(net44),
    .GATE(\genblk1[54].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[54][6] ));
 sky130_fd_sc_hd__dlxtp_1 _1096_ (.D(net35),
    .GATE(\genblk1[54].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[54][7] ));
 sky130_fd_sc_hd__dlxtp_1 _1097_ (.D(net93),
    .GATE(\genblk1[53].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[53][0] ));
 sky130_fd_sc_hd__dlxtp_1 _1098_ (.D(net86),
    .GATE(\genblk1[53].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[53][1] ));
 sky130_fd_sc_hd__dlxtp_1 _1099_ (.D(net78),
    .GATE(\genblk1[53].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[53][2] ));
 sky130_fd_sc_hd__dlxtp_1 _1100_ (.D(net69),
    .GATE(\genblk1[53].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[53][3] ));
 sky130_fd_sc_hd__dlxtp_1 _1101_ (.D(\data_to_write[4] ),
    .GATE(\genblk1[53].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[53][4] ));
 sky130_fd_sc_hd__dlxtp_1 _1102_ (.D(net53),
    .GATE(\genblk1[53].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[53][5] ));
 sky130_fd_sc_hd__dlxtp_1 _1103_ (.D(net44),
    .GATE(\genblk1[53].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[53][6] ));
 sky130_fd_sc_hd__dlxtp_1 _1104_ (.D(net34),
    .GATE(\genblk1[53].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[53][7] ));
 sky130_fd_sc_hd__dlxtp_1 _1105_ (.D(net93),
    .GATE(\genblk1[52].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[52][0] ));
 sky130_fd_sc_hd__dlxtp_1 _1106_ (.D(net87),
    .GATE(\genblk1[52].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[52][1] ));
 sky130_fd_sc_hd__dlxtp_1 _1107_ (.D(net77),
    .GATE(\genblk1[52].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[52][2] ));
 sky130_fd_sc_hd__dlxtp_1 _1108_ (.D(net68),
    .GATE(\genblk1[52].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[52][3] ));
 sky130_fd_sc_hd__dlxtp_1 _1109_ (.D(net60),
    .GATE(\genblk1[52].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[52][4] ));
 sky130_fd_sc_hd__dlxtp_1 _1110_ (.D(net54),
    .GATE(\genblk1[52].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[52][5] ));
 sky130_fd_sc_hd__dlxtp_1 _1111_ (.D(net44),
    .GATE(\genblk1[52].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[52][6] ));
 sky130_fd_sc_hd__dlxtp_1 _1112_ (.D(net37),
    .GATE(\genblk1[52].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[52][7] ));
 sky130_fd_sc_hd__dlxtp_1 _1113_ (.D(net93),
    .GATE(\genblk1[51].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[51][0] ));
 sky130_fd_sc_hd__dlxtp_1 _1114_ (.D(net85),
    .GATE(\genblk1[51].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[51][1] ));
 sky130_fd_sc_hd__dlxtp_1 _1115_ (.D(net77),
    .GATE(\genblk1[51].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[51][2] ));
 sky130_fd_sc_hd__dlxtp_1 _1116_ (.D(net70),
    .GATE(\genblk1[51].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[51][3] ));
 sky130_fd_sc_hd__dlxtp_1 _1117_ (.D(net62),
    .GATE(\genblk1[51].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[51][4] ));
 sky130_fd_sc_hd__dlxtp_1 _1118_ (.D(net52),
    .GATE(\genblk1[51].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[51][5] ));
 sky130_fd_sc_hd__dlxtp_1 _1119_ (.D(net44),
    .GATE(\genblk1[51].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[51][6] ));
 sky130_fd_sc_hd__dlxtp_1 _1120_ (.D(net37),
    .GATE(\genblk1[51].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[51][7] ));
 sky130_fd_sc_hd__dlxtp_1 _1121_ (.D(net94),
    .GATE(\genblk1[50].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[50][0] ));
 sky130_fd_sc_hd__dlxtp_1 _1122_ (.D(net85),
    .GATE(\genblk1[50].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[50][1] ));
 sky130_fd_sc_hd__dlxtp_1 _1123_ (.D(net77),
    .GATE(\genblk1[50].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[50][2] ));
 sky130_fd_sc_hd__dlxtp_1 _1124_ (.D(net68),
    .GATE(\genblk1[50].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[50][3] ));
 sky130_fd_sc_hd__dlxtp_1 _1125_ (.D(net60),
    .GATE(\genblk1[50].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[50][4] ));
 sky130_fd_sc_hd__dlxtp_1 _1126_ (.D(net52),
    .GATE(\genblk1[50].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[50][5] ));
 sky130_fd_sc_hd__dlxtp_1 _1127_ (.D(net44),
    .GATE(\genblk1[50].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[50][6] ));
 sky130_fd_sc_hd__dlxtp_1 _1128_ (.D(net35),
    .GATE(\genblk1[50].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[50][7] ));
 sky130_fd_sc_hd__dlxtp_1 _1129_ (.D(net93),
    .GATE(\genblk1[49].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[49][0] ));
 sky130_fd_sc_hd__dlxtp_1 _1130_ (.D(net85),
    .GATE(\genblk1[49].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[49][1] ));
 sky130_fd_sc_hd__dlxtp_1 _1131_ (.D(net78),
    .GATE(\genblk1[49].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[49][2] ));
 sky130_fd_sc_hd__dlxtp_1 _1132_ (.D(net68),
    .GATE(\genblk1[49].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[49][3] ));
 sky130_fd_sc_hd__dlxtp_1 _1133_ (.D(net60),
    .GATE(\genblk1[49].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[49][4] ));
 sky130_fd_sc_hd__dlxtp_1 _1134_ (.D(net52),
    .GATE(\genblk1[49].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[49][5] ));
 sky130_fd_sc_hd__dlxtp_1 _1135_ (.D(net44),
    .GATE(\genblk1[49].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[49][6] ));
 sky130_fd_sc_hd__dlxtp_1 _1136_ (.D(net34),
    .GATE(\genblk1[49].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[49][7] ));
 sky130_fd_sc_hd__dlxtp_1 _1137_ (.D(net93),
    .GATE(\genblk1[48].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[48][0] ));
 sky130_fd_sc_hd__dlxtp_1 _1138_ (.D(net85),
    .GATE(\genblk1[48].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[48][1] ));
 sky130_fd_sc_hd__dlxtp_1 _1139_ (.D(net77),
    .GATE(\genblk1[48].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[48][2] ));
 sky130_fd_sc_hd__dlxtp_1 _1140_ (.D(net68),
    .GATE(\genblk1[48].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[48][3] ));
 sky130_fd_sc_hd__dlxtp_1 _1141_ (.D(net59),
    .GATE(\genblk1[48].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[48][4] ));
 sky130_fd_sc_hd__dlxtp_1 _1142_ (.D(net52),
    .GATE(\genblk1[48].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[48][5] ));
 sky130_fd_sc_hd__dlxtp_1 _1143_ (.D(net45),
    .GATE(\genblk1[48].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[48][6] ));
 sky130_fd_sc_hd__dlxtp_1 _1144_ (.D(net34),
    .GATE(\genblk1[48].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[48][7] ));
 sky130_fd_sc_hd__dlxtp_1 _1145_ (.D(net95),
    .GATE(\genblk1[47].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[47][0] ));
 sky130_fd_sc_hd__dlxtp_1 _1146_ (.D(net84),
    .GATE(\genblk1[47].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[47][1] ));
 sky130_fd_sc_hd__dlxtp_1 _1147_ (.D(net72),
    .GATE(\genblk1[47].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[47][2] ));
 sky130_fd_sc_hd__dlxtp_1 _1148_ (.D(net63),
    .GATE(\genblk1[47].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[47][3] ));
 sky130_fd_sc_hd__dlxtp_1 _1149_ (.D(net61),
    .GATE(\genblk1[47].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[47][4] ));
 sky130_fd_sc_hd__dlxtp_1 _1150_ (.D(net54),
    .GATE(\genblk1[47].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[47][5] ));
 sky130_fd_sc_hd__dlxtp_1 _1151_ (.D(net42),
    .GATE(\genblk1[47].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[47][6] ));
 sky130_fd_sc_hd__dlxtp_1 _1152_ (.D(net33),
    .GATE(\genblk1[47].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[47][7] ));
 sky130_fd_sc_hd__dlxtp_1 _1153_ (.D(net92),
    .GATE(\genblk1[46].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[46][0] ));
 sky130_fd_sc_hd__dlxtp_1 _1154_ (.D(net84),
    .GATE(\genblk1[46].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[46][1] ));
 sky130_fd_sc_hd__dlxtp_1 _1155_ (.D(net72),
    .GATE(\genblk1[46].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[46][2] ));
 sky130_fd_sc_hd__dlxtp_1 _1156_ (.D(net63),
    .GATE(\genblk1[46].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[46][3] ));
 sky130_fd_sc_hd__dlxtp_1 _1157_ (.D(net61),
    .GATE(\genblk1[46].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[46][4] ));
 sky130_fd_sc_hd__dlxtp_1 _1158_ (.D(net53),
    .GATE(\genblk1[46].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[46][5] ));
 sky130_fd_sc_hd__dlxtp_1 _1159_ (.D(net42),
    .GATE(\genblk1[46].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[46][6] ));
 sky130_fd_sc_hd__dlxtp_1 _1160_ (.D(net33),
    .GATE(\genblk1[46].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[46][7] ));
 sky130_fd_sc_hd__dlxtp_1 _1161_ (.D(net92),
    .GATE(\genblk1[45].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[45][0] ));
 sky130_fd_sc_hd__dlxtp_1 _1162_ (.D(net84),
    .GATE(\genblk1[45].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[45][1] ));
 sky130_fd_sc_hd__dlxtp_1 _1163_ (.D(net73),
    .GATE(\genblk1[45].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[45][2] ));
 sky130_fd_sc_hd__dlxtp_1 _1164_ (.D(net63),
    .GATE(\genblk1[45].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[45][3] ));
 sky130_fd_sc_hd__dlxtp_1 _1165_ (.D(net59),
    .GATE(\genblk1[45].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[45][4] ));
 sky130_fd_sc_hd__dlxtp_1 _1166_ (.D(net53),
    .GATE(\genblk1[45].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[45][5] ));
 sky130_fd_sc_hd__dlxtp_1 _1167_ (.D(net43),
    .GATE(\genblk1[45].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[45][6] ));
 sky130_fd_sc_hd__dlxtp_1 _1168_ (.D(net33),
    .GATE(\genblk1[45].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[45][7] ));
 sky130_fd_sc_hd__dlxtp_1 _1169_ (.D(net92),
    .GATE(\genblk1[44].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[44][0] ));
 sky130_fd_sc_hd__dlxtp_1 _1170_ (.D(net84),
    .GATE(\genblk1[44].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[44][1] ));
 sky130_fd_sc_hd__dlxtp_1 _1171_ (.D(net74),
    .GATE(\genblk1[44].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[44][2] ));
 sky130_fd_sc_hd__dlxtp_1 _1172_ (.D(net63),
    .GATE(\genblk1[44].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[44][3] ));
 sky130_fd_sc_hd__dlxtp_1 _1173_ (.D(net61),
    .GATE(\genblk1[44].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[44][4] ));
 sky130_fd_sc_hd__dlxtp_1 _1174_ (.D(net50),
    .GATE(\genblk1[44].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[44][5] ));
 sky130_fd_sc_hd__dlxtp_1 _1175_ (.D(net42),
    .GATE(\genblk1[44].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[44][6] ));
 sky130_fd_sc_hd__dlxtp_1 _1176_ (.D(net35),
    .GATE(\genblk1[44].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[44][7] ));
 sky130_fd_sc_hd__dlxtp_1 _1177_ (.D(net95),
    .GATE(\genblk1[43].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[43][0] ));
 sky130_fd_sc_hd__dlxtp_1 _1178_ (.D(net86),
    .GATE(\genblk1[43].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[43][1] ));
 sky130_fd_sc_hd__dlxtp_1 _1179_ (.D(net74),
    .GATE(\genblk1[43].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[43][2] ));
 sky130_fd_sc_hd__dlxtp_1 _1180_ (.D(net70),
    .GATE(\genblk1[43].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[43][3] ));
 sky130_fd_sc_hd__dlxtp_1 _1181_ (.D(net61),
    .GATE(\genblk1[43].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[43][4] ));
 sky130_fd_sc_hd__dlxtp_1 _1182_ (.D(net48),
    .GATE(\genblk1[43].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[43][5] ));
 sky130_fd_sc_hd__dlxtp_1 _1183_ (.D(net43),
    .GATE(\genblk1[43].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[43][6] ));
 sky130_fd_sc_hd__dlxtp_1 _1184_ (.D(net30),
    .GATE(\genblk1[43].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[43][7] ));
 sky130_fd_sc_hd__dlxtp_1 _1185_ (.D(net92),
    .GATE(\genblk1[42].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[42][0] ));
 sky130_fd_sc_hd__dlxtp_1 _1186_ (.D(net86),
    .GATE(\genblk1[42].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[42][1] ));
 sky130_fd_sc_hd__dlxtp_1 _1187_ (.D(net72),
    .GATE(\genblk1[42].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[42][2] ));
 sky130_fd_sc_hd__dlxtp_1 _1188_ (.D(net67),
    .GATE(\genblk1[42].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[42][3] ));
 sky130_fd_sc_hd__dlxtp_1 _1189_ (.D(net61),
    .GATE(\genblk1[42].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[42][4] ));
 sky130_fd_sc_hd__dlxtp_1 _1190_ (.D(net50),
    .GATE(\genblk1[42].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[42][5] ));
 sky130_fd_sc_hd__dlxtp_1 _1191_ (.D(net42),
    .GATE(\genblk1[42].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[42][6] ));
 sky130_fd_sc_hd__dlxtp_1 _1192_ (.D(net30),
    .GATE(\genblk1[42].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[42][7] ));
 sky130_fd_sc_hd__dlxtp_1 _1193_ (.D(net92),
    .GATE(\genblk1[41].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[41][0] ));
 sky130_fd_sc_hd__dlxtp_1 _1194_ (.D(net84),
    .GATE(\genblk1[41].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[41][1] ));
 sky130_fd_sc_hd__dlxtp_1 _1195_ (.D(net72),
    .GATE(\genblk1[41].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[41][2] ));
 sky130_fd_sc_hd__dlxtp_1 _1196_ (.D(net68),
    .GATE(\genblk1[41].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[41][3] ));
 sky130_fd_sc_hd__dlxtp_1 _1197_ (.D(net59),
    .GATE(\genblk1[41].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[41][4] ));
 sky130_fd_sc_hd__dlxtp_1 _1198_ (.D(net48),
    .GATE(\genblk1[41].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[41][5] ));
 sky130_fd_sc_hd__dlxtp_1 _1199_ (.D(net42),
    .GATE(\genblk1[41].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[41][6] ));
 sky130_fd_sc_hd__dlxtp_1 _1200_ (.D(net33),
    .GATE(\genblk1[41].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[41][7] ));
 sky130_fd_sc_hd__dlxtp_1 _1201_ (.D(net92),
    .GATE(\genblk1[40].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[40][0] ));
 sky130_fd_sc_hd__dlxtp_1 _1202_ (.D(net83),
    .GATE(\genblk1[40].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[40][1] ));
 sky130_fd_sc_hd__dlxtp_1 _1203_ (.D(net73),
    .GATE(\genblk1[40].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[40][2] ));
 sky130_fd_sc_hd__dlxtp_1 _1204_ (.D(net63),
    .GATE(\genblk1[40].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[40][3] ));
 sky130_fd_sc_hd__dlxtp_1 _1205_ (.D(net61),
    .GATE(\genblk1[40].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[40][4] ));
 sky130_fd_sc_hd__dlxtp_1 _1206_ (.D(net48),
    .GATE(\genblk1[40].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[40][5] ));
 sky130_fd_sc_hd__dlxtp_1 _1207_ (.D(net42),
    .GATE(\genblk1[40].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[40][6] ));
 sky130_fd_sc_hd__dlxtp_1 _1208_ (.D(net33),
    .GATE(\genblk1[40].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[40][7] ));
 sky130_fd_sc_hd__dlxtp_1 _1209_ (.D(net92),
    .GATE(\genblk1[39].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[39][0] ));
 sky130_fd_sc_hd__dlxtp_1 _1210_ (.D(net84),
    .GATE(\genblk1[39].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[39][1] ));
 sky130_fd_sc_hd__dlxtp_1 _1211_ (.D(net73),
    .GATE(\genblk1[39].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[39][2] ));
 sky130_fd_sc_hd__dlxtp_1 _1212_ (.D(net68),
    .GATE(\genblk1[39].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[39][3] ));
 sky130_fd_sc_hd__dlxtp_1 _1213_ (.D(net59),
    .GATE(\genblk1[39].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[39][4] ));
 sky130_fd_sc_hd__dlxtp_1 _1214_ (.D(net48),
    .GATE(\genblk1[39].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[39][5] ));
 sky130_fd_sc_hd__dlxtp_1 _1215_ (.D(net43),
    .GATE(\genblk1[39].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[39][6] ));
 sky130_fd_sc_hd__dlxtp_1 _1216_ (.D(net33),
    .GATE(\genblk1[39].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[39][7] ));
 sky130_fd_sc_hd__dlxtp_1 _1217_ (.D(net92),
    .GATE(\genblk1[38].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[38][0] ));
 sky130_fd_sc_hd__dlxtp_1 _1218_ (.D(net86),
    .GATE(\genblk1[38].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[38][1] ));
 sky130_fd_sc_hd__dlxtp_1 _1219_ (.D(net72),
    .GATE(\genblk1[38].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[38][2] ));
 sky130_fd_sc_hd__dlxtp_1 _1220_ (.D(net68),
    .GATE(\genblk1[38].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[38][3] ));
 sky130_fd_sc_hd__dlxtp_1 _1221_ (.D(net59),
    .GATE(\genblk1[38].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[38][4] ));
 sky130_fd_sc_hd__dlxtp_1 _1222_ (.D(net48),
    .GATE(\genblk1[38].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[38][5] ));
 sky130_fd_sc_hd__dlxtp_1 _1223_ (.D(net42),
    .GATE(\genblk1[38].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[38][6] ));
 sky130_fd_sc_hd__dlxtp_1 _1224_ (.D(net30),
    .GATE(\genblk1[38].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[38][7] ));
 sky130_fd_sc_hd__dlxtp_1 _1225_ (.D(net95),
    .GATE(\genblk1[37].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[37][0] ));
 sky130_fd_sc_hd__dlxtp_1 _1226_ (.D(net84),
    .GATE(\genblk1[37].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[37][1] ));
 sky130_fd_sc_hd__dlxtp_1 _1227_ (.D(net74),
    .GATE(\genblk1[37].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[37][2] ));
 sky130_fd_sc_hd__dlxtp_1 _1228_ (.D(net67),
    .GATE(\genblk1[37].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[37][3] ));
 sky130_fd_sc_hd__dlxtp_1 _1229_ (.D(net59),
    .GATE(\genblk1[37].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[37][4] ));
 sky130_fd_sc_hd__dlxtp_1 _1230_ (.D(net50),
    .GATE(\genblk1[37].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[37][5] ));
 sky130_fd_sc_hd__dlxtp_1 _1231_ (.D(net42),
    .GATE(\genblk1[37].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[37][6] ));
 sky130_fd_sc_hd__dlxtp_1 _1232_ (.D(net35),
    .GATE(\genblk1[37].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[37][7] ));
 sky130_fd_sc_hd__dlxtp_1 _1233_ (.D(net92),
    .GATE(\genblk1[36].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[36][0] ));
 sky130_fd_sc_hd__dlxtp_1 _1234_ (.D(net84),
    .GATE(\genblk1[36].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[36][1] ));
 sky130_fd_sc_hd__dlxtp_1 _1235_ (.D(net72),
    .GATE(\genblk1[36].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[36][2] ));
 sky130_fd_sc_hd__dlxtp_1 _1236_ (.D(net63),
    .GATE(\genblk1[36].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[36][3] ));
 sky130_fd_sc_hd__dlxtp_1 _1237_ (.D(net59),
    .GATE(\genblk1[36].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[36][4] ));
 sky130_fd_sc_hd__dlxtp_1 _1238_ (.D(net48),
    .GATE(\genblk1[36].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[36][5] ));
 sky130_fd_sc_hd__dlxtp_1 _1239_ (.D(net43),
    .GATE(\genblk1[36].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[36][6] ));
 sky130_fd_sc_hd__dlxtp_1 _1240_ (.D(net30),
    .GATE(\genblk1[36].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[36][7] ));
 sky130_fd_sc_hd__dlxtp_1 _1241_ (.D(net95),
    .GATE(\genblk1[35].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[35][0] ));
 sky130_fd_sc_hd__dlxtp_1 _1242_ (.D(net83),
    .GATE(\genblk1[35].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[35][1] ));
 sky130_fd_sc_hd__dlxtp_1 _1243_ (.D(net73),
    .GATE(\genblk1[35].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[35][2] ));
 sky130_fd_sc_hd__dlxtp_1 _1244_ (.D(net63),
    .GATE(\genblk1[35].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[35][3] ));
 sky130_fd_sc_hd__dlxtp_1 _1245_ (.D(net59),
    .GATE(\genblk1[35].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[35][4] ));
 sky130_fd_sc_hd__dlxtp_1 _1246_ (.D(net48),
    .GATE(\genblk1[35].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[35][5] ));
 sky130_fd_sc_hd__dlxtp_1 _1247_ (.D(net42),
    .GATE(\genblk1[35].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[35][6] ));
 sky130_fd_sc_hd__dlxtp_1 _1248_ (.D(net33),
    .GATE(\genblk1[35].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[35][7] ));
 sky130_fd_sc_hd__dlxtp_1 _1249_ (.D(net94),
    .GATE(\genblk1[34].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[34][0] ));
 sky130_fd_sc_hd__dlxtp_1 _1250_ (.D(net84),
    .GATE(\genblk1[34].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[34][1] ));
 sky130_fd_sc_hd__dlxtp_1 _1251_ (.D(net73),
    .GATE(\genblk1[34].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[34][2] ));
 sky130_fd_sc_hd__dlxtp_1 _1252_ (.D(net63),
    .GATE(\genblk1[34].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[34][3] ));
 sky130_fd_sc_hd__dlxtp_1 _1253_ (.D(net61),
    .GATE(\genblk1[34].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[34][4] ));
 sky130_fd_sc_hd__dlxtp_1 _1254_ (.D(net49),
    .GATE(\genblk1[34].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[34][5] ));
 sky130_fd_sc_hd__dlxtp_1 _1255_ (.D(net43),
    .GATE(\genblk1[34].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[34][6] ));
 sky130_fd_sc_hd__dlxtp_1 _1256_ (.D(net33),
    .GATE(\genblk1[34].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[34][7] ));
 sky130_fd_sc_hd__dlxtp_1 _1257_ (.D(net94),
    .GATE(\genblk1[33].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[33][0] ));
 sky130_fd_sc_hd__dlxtp_1 _1258_ (.D(net86),
    .GATE(\genblk1[33].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[33][1] ));
 sky130_fd_sc_hd__dlxtp_1 _1259_ (.D(net74),
    .GATE(\genblk1[33].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[33][2] ));
 sky130_fd_sc_hd__dlxtp_1 _1260_ (.D(net67),
    .GATE(\genblk1[33].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[33][3] ));
 sky130_fd_sc_hd__dlxtp_1 _1261_ (.D(net61),
    .GATE(\genblk1[33].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[33][4] ));
 sky130_fd_sc_hd__dlxtp_1 _1262_ (.D(net54),
    .GATE(\genblk1[33].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[33][5] ));
 sky130_fd_sc_hd__dlxtp_1 _1263_ (.D(net43),
    .GATE(\genblk1[33].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[33][6] ));
 sky130_fd_sc_hd__dlxtp_1 _1264_ (.D(net33),
    .GATE(\genblk1[33].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[33][7] ));
 sky130_fd_sc_hd__dlxtp_1 _1265_ (.D(net92),
    .GATE(\genblk1[32].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[32][0] ));
 sky130_fd_sc_hd__dlxtp_1 _1266_ (.D(net84),
    .GATE(\genblk1[32].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[32][1] ));
 sky130_fd_sc_hd__dlxtp_1 _1267_ (.D(net72),
    .GATE(\genblk1[32].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[32][2] ));
 sky130_fd_sc_hd__dlxtp_1 _1268_ (.D(net68),
    .GATE(\genblk1[32].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[32][3] ));
 sky130_fd_sc_hd__dlxtp_1 _1269_ (.D(net61),
    .GATE(\genblk1[32].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[32][4] ));
 sky130_fd_sc_hd__dlxtp_1 _1270_ (.D(net50),
    .GATE(\genblk1[32].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[32][5] ));
 sky130_fd_sc_hd__dlxtp_1 _1271_ (.D(net42),
    .GATE(\genblk1[32].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[32][6] ));
 sky130_fd_sc_hd__dlxtp_1 _1272_ (.D(net33),
    .GATE(\genblk1[32].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[32][7] ));
 sky130_fd_sc_hd__dlxtp_1 _1273_ (.D(net90),
    .GATE(\genblk1[31].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[31][0] ));
 sky130_fd_sc_hd__dlxtp_1 _1274_ (.D(net80),
    .GATE(\genblk1[31].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[31][1] ));
 sky130_fd_sc_hd__dlxtp_1 _1275_ (.D(net71),
    .GATE(\genblk1[31].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[31][2] ));
 sky130_fd_sc_hd__dlxtp_1 _1276_ (.D(net63),
    .GATE(\genblk1[31].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[31][3] ));
 sky130_fd_sc_hd__dlxtp_1 _1277_ (.D(net56),
    .GATE(\genblk1[31].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[31][4] ));
 sky130_fd_sc_hd__dlxtp_1 _1278_ (.D(net47),
    .GATE(\genblk1[31].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[31][5] ));
 sky130_fd_sc_hd__dlxtp_1 _1279_ (.D(net38),
    .GATE(\genblk1[31].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[31][6] ));
 sky130_fd_sc_hd__dlxtp_1 _1280_ (.D(net31),
    .GATE(\genblk1[31].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[31][7] ));
 sky130_fd_sc_hd__dlxtp_1 _1281_ (.D(net88),
    .GATE(\genblk1[30].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[30][0] ));
 sky130_fd_sc_hd__dlxtp_1 _1282_ (.D(net79),
    .GATE(\genblk1[30].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[30][1] ));
 sky130_fd_sc_hd__dlxtp_1 _1283_ (.D(net72),
    .GATE(\genblk1[30].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[30][2] ));
 sky130_fd_sc_hd__dlxtp_1 _1284_ (.D(net65),
    .GATE(\genblk1[30].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[30][3] ));
 sky130_fd_sc_hd__dlxtp_1 _1285_ (.D(net55),
    .GATE(\genblk1[30].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[30][4] ));
 sky130_fd_sc_hd__dlxtp_1 _1286_ (.D(net49),
    .GATE(\genblk1[30].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[30][5] ));
 sky130_fd_sc_hd__dlxtp_1 _1287_ (.D(net40),
    .GATE(\genblk1[30].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[30][6] ));
 sky130_fd_sc_hd__dlxtp_1 _1288_ (.D(net31),
    .GATE(\genblk1[30].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[30][7] ));
 sky130_fd_sc_hd__dlxtp_1 _1289_ (.D(net88),
    .GATE(\genblk1[29].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[29][0] ));
 sky130_fd_sc_hd__dlxtp_1 _1290_ (.D(net79),
    .GATE(\genblk1[29].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[29][1] ));
 sky130_fd_sc_hd__dlxtp_1 _1291_ (.D(net71),
    .GATE(\genblk1[29].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[29][2] ));
 sky130_fd_sc_hd__dlxtp_1 _1292_ (.D(net65),
    .GATE(\genblk1[29].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[29][3] ));
 sky130_fd_sc_hd__dlxtp_1 _1293_ (.D(net56),
    .GATE(\genblk1[29].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[29][4] ));
 sky130_fd_sc_hd__dlxtp_1 _1294_ (.D(net48),
    .GATE(\genblk1[29].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[29][5] ));
 sky130_fd_sc_hd__dlxtp_1 _1295_ (.D(net38),
    .GATE(\genblk1[29].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[29][6] ));
 sky130_fd_sc_hd__dlxtp_1 _1296_ (.D(net29),
    .GATE(\genblk1[29].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[29][7] ));
 sky130_fd_sc_hd__dlxtp_1 _1297_ (.D(net88),
    .GATE(\genblk1[28].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[28][0] ));
 sky130_fd_sc_hd__dlxtp_1 _1298_ (.D(net80),
    .GATE(\genblk1[28].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[28][1] ));
 sky130_fd_sc_hd__dlxtp_1 _1299_ (.D(net71),
    .GATE(\genblk1[28].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[28][2] ));
 sky130_fd_sc_hd__dlxtp_1 _1300_ (.D(net64),
    .GATE(\genblk1[28].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[28][3] ));
 sky130_fd_sc_hd__dlxtp_1 _1301_ (.D(net55),
    .GATE(\genblk1[28].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[28][4] ));
 sky130_fd_sc_hd__dlxtp_1 _1302_ (.D(net47),
    .GATE(\genblk1[28].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[28][5] ));
 sky130_fd_sc_hd__dlxtp_1 _1303_ (.D(net38),
    .GATE(\genblk1[28].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[28][6] ));
 sky130_fd_sc_hd__dlxtp_1 _1304_ (.D(net29),
    .GATE(\genblk1[28].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[28][7] ));
 sky130_fd_sc_hd__dlxtp_1 _1305_ (.D(net91),
    .GATE(\genblk1[27].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[27][0] ));
 sky130_fd_sc_hd__dlxtp_1 _1306_ (.D(net80),
    .GATE(\genblk1[27].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[27][1] ));
 sky130_fd_sc_hd__dlxtp_1 _1307_ (.D(net71),
    .GATE(\genblk1[27].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[27][2] ));
 sky130_fd_sc_hd__dlxtp_1 _1308_ (.D(net64),
    .GATE(\genblk1[27].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[27][3] ));
 sky130_fd_sc_hd__dlxtp_1 _1309_ (.D(net56),
    .GATE(\genblk1[27].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[27][4] ));
 sky130_fd_sc_hd__dlxtp_1 _1310_ (.D(net47),
    .GATE(\genblk1[27].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[27][5] ));
 sky130_fd_sc_hd__dlxtp_1 _1311_ (.D(net40),
    .GATE(\genblk1[27].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[27][6] ));
 sky130_fd_sc_hd__dlxtp_1 _1312_ (.D(net29),
    .GATE(\genblk1[27].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[27][7] ));
 sky130_fd_sc_hd__dlxtp_1 _1313_ (.D(net90),
    .GATE(\genblk1[26].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[26][0] ));
 sky130_fd_sc_hd__dlxtp_1 _1314_ (.D(net80),
    .GATE(\genblk1[26].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[26][1] ));
 sky130_fd_sc_hd__dlxtp_1 _1315_ (.D(net71),
    .GATE(\genblk1[26].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[26][2] ));
 sky130_fd_sc_hd__dlxtp_1 _1316_ (.D(net64),
    .GATE(\genblk1[26].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[26][3] ));
 sky130_fd_sc_hd__dlxtp_1 _1317_ (.D(net55),
    .GATE(\genblk1[26].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[26][4] ));
 sky130_fd_sc_hd__dlxtp_1 _1318_ (.D(net49),
    .GATE(\genblk1[26].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[26][5] ));
 sky130_fd_sc_hd__dlxtp_1 _1319_ (.D(net39),
    .GATE(\genblk1[26].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[26][6] ));
 sky130_fd_sc_hd__dlxtp_1 _1320_ (.D(net29),
    .GATE(\genblk1[26].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[26][7] ));
 sky130_fd_sc_hd__dlxtp_1 _1321_ (.D(net90),
    .GATE(\genblk1[25].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[25][0] ));
 sky130_fd_sc_hd__dlxtp_1 _1322_ (.D(net79),
    .GATE(\genblk1[25].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[25][1] ));
 sky130_fd_sc_hd__dlxtp_1 _1323_ (.D(net72),
    .GATE(\genblk1[25].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[25][2] ));
 sky130_fd_sc_hd__dlxtp_1 _1324_ (.D(net64),
    .GATE(\genblk1[25].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[25][3] ));
 sky130_fd_sc_hd__dlxtp_1 _1325_ (.D(net56),
    .GATE(\genblk1[25].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[25][4] ));
 sky130_fd_sc_hd__dlxtp_1 _1326_ (.D(net47),
    .GATE(\genblk1[25].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[25][5] ));
 sky130_fd_sc_hd__dlxtp_1 _1327_ (.D(net39),
    .GATE(\genblk1[25].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[25][6] ));
 sky130_fd_sc_hd__dlxtp_1 _1328_ (.D(net29),
    .GATE(\genblk1[25].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[25][7] ));
 sky130_fd_sc_hd__dlxtp_1 _1329_ (.D(net88),
    .GATE(\genblk1[24].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[24][0] ));
 sky130_fd_sc_hd__dlxtp_1 _1330_ (.D(net80),
    .GATE(\genblk1[24].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[24][1] ));
 sky130_fd_sc_hd__dlxtp_1 _1331_ (.D(net73),
    .GATE(\genblk1[24].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[24][2] ));
 sky130_fd_sc_hd__dlxtp_1 _1332_ (.D(net64),
    .GATE(\genblk1[24].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[24][3] ));
 sky130_fd_sc_hd__dlxtp_1 _1333_ (.D(net55),
    .GATE(\genblk1[24].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[24][4] ));
 sky130_fd_sc_hd__dlxtp_1 _1334_ (.D(net47),
    .GATE(\genblk1[24].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[24][5] ));
 sky130_fd_sc_hd__dlxtp_1 _1335_ (.D(net38),
    .GATE(\genblk1[24].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[24][6] ));
 sky130_fd_sc_hd__dlxtp_1 _1336_ (.D(net29),
    .GATE(\genblk1[24].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[24][7] ));
 sky130_fd_sc_hd__dlxtp_1 _1337_ (.D(net88),
    .GATE(\genblk1[23].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[23][0] ));
 sky130_fd_sc_hd__dlxtp_1 _1338_ (.D(net79),
    .GATE(\genblk1[23].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[23][1] ));
 sky130_fd_sc_hd__dlxtp_1 _1339_ (.D(net71),
    .GATE(\genblk1[23].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[23][2] ));
 sky130_fd_sc_hd__dlxtp_1 _1340_ (.D(net63),
    .GATE(\genblk1[23].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[23][3] ));
 sky130_fd_sc_hd__dlxtp_1 _1341_ (.D(net55),
    .GATE(\genblk1[23].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[23][4] ));
 sky130_fd_sc_hd__dlxtp_1 _1342_ (.D(net48),
    .GATE(\genblk1[23].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[23][5] ));
 sky130_fd_sc_hd__dlxtp_1 _1343_ (.D(net39),
    .GATE(\genblk1[23].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[23][6] ));
 sky130_fd_sc_hd__dlxtp_1 _1344_ (.D(net31),
    .GATE(\genblk1[23].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[23][7] ));
 sky130_fd_sc_hd__dlxtp_1 _1345_ (.D(net88),
    .GATE(\genblk1[22].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[22][0] ));
 sky130_fd_sc_hd__dlxtp_1 _1346_ (.D(net79),
    .GATE(\genblk1[22].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[22][1] ));
 sky130_fd_sc_hd__dlxtp_1 _1347_ (.D(net71),
    .GATE(\genblk1[22].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[22][2] ));
 sky130_fd_sc_hd__dlxtp_1 _1348_ (.D(net64),
    .GATE(\genblk1[22].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[22][3] ));
 sky130_fd_sc_hd__dlxtp_1 _1349_ (.D(net55),
    .GATE(\genblk1[22].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[22][4] ));
 sky130_fd_sc_hd__dlxtp_1 _1350_ (.D(net48),
    .GATE(\genblk1[22].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[22][5] ));
 sky130_fd_sc_hd__dlxtp_1 _1351_ (.D(net38),
    .GATE(\genblk1[22].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[22][6] ));
 sky130_fd_sc_hd__dlxtp_1 _1352_ (.D(net30),
    .GATE(\genblk1[22].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[22][7] ));
 sky130_fd_sc_hd__dlxtp_1 _1353_ (.D(net88),
    .GATE(\genblk1[21].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[21][0] ));
 sky130_fd_sc_hd__dlxtp_1 _1354_ (.D(net79),
    .GATE(\genblk1[21].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[21][1] ));
 sky130_fd_sc_hd__dlxtp_1 _1355_ (.D(net73),
    .GATE(\genblk1[21].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[21][2] ));
 sky130_fd_sc_hd__dlxtp_1 _1356_ (.D(net65),
    .GATE(\genblk1[21].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[21][3] ));
 sky130_fd_sc_hd__dlxtp_1 _1357_ (.D(net55),
    .GATE(\genblk1[21].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[21][4] ));
 sky130_fd_sc_hd__dlxtp_1 _1358_ (.D(net47),
    .GATE(\genblk1[21].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[21][5] ));
 sky130_fd_sc_hd__dlxtp_1 _1359_ (.D(net38),
    .GATE(\genblk1[21].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[21][6] ));
 sky130_fd_sc_hd__dlxtp_1 _1360_ (.D(net31),
    .GATE(\genblk1[21].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[21][7] ));
 sky130_fd_sc_hd__dlxtp_1 _1361_ (.D(net88),
    .GATE(\genblk1[20].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[20][0] ));
 sky130_fd_sc_hd__dlxtp_1 _1362_ (.D(net79),
    .GATE(\genblk1[20].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[20][1] ));
 sky130_fd_sc_hd__dlxtp_1 _1363_ (.D(net73),
    .GATE(\genblk1[20].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[20][2] ));
 sky130_fd_sc_hd__dlxtp_1 _1364_ (.D(net70),
    .GATE(\genblk1[20].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[20][3] ));
 sky130_fd_sc_hd__dlxtp_1 _1365_ (.D(net56),
    .GATE(\genblk1[20].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[20][4] ));
 sky130_fd_sc_hd__dlxtp_1 _1366_ (.D(net47),
    .GATE(\genblk1[20].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[20][5] ));
 sky130_fd_sc_hd__dlxtp_1 _1367_ (.D(net38),
    .GATE(\genblk1[20].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[20][6] ));
 sky130_fd_sc_hd__dlxtp_1 _1368_ (.D(net29),
    .GATE(\genblk1[20].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[20][7] ));
 sky130_fd_sc_hd__dlxtp_1 _1369_ (.D(net90),
    .GATE(\genblk1[19].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[19][0] ));
 sky130_fd_sc_hd__dlxtp_1 _1370_ (.D(net79),
    .GATE(\genblk1[19].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[19][1] ));
 sky130_fd_sc_hd__dlxtp_1 _1371_ (.D(net71),
    .GATE(\genblk1[19].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[19][2] ));
 sky130_fd_sc_hd__dlxtp_1 _1372_ (.D(net64),
    .GATE(\genblk1[19].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[19][3] ));
 sky130_fd_sc_hd__dlxtp_1 _1373_ (.D(net55),
    .GATE(\genblk1[19].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[19][4] ));
 sky130_fd_sc_hd__dlxtp_1 _1374_ (.D(net49),
    .GATE(\genblk1[19].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[19][5] ));
 sky130_fd_sc_hd__dlxtp_1 _1375_ (.D(net38),
    .GATE(\genblk1[19].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[19][6] ));
 sky130_fd_sc_hd__dlxtp_1 _1376_ (.D(net29),
    .GATE(\genblk1[19].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[19][7] ));
 sky130_fd_sc_hd__dlxtp_1 _1377_ (.D(net88),
    .GATE(\genblk1[18].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[18][0] ));
 sky130_fd_sc_hd__dlxtp_1 _1378_ (.D(net79),
    .GATE(\genblk1[18].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[18][1] ));
 sky130_fd_sc_hd__dlxtp_1 _1379_ (.D(net71),
    .GATE(\genblk1[18].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[18][2] ));
 sky130_fd_sc_hd__dlxtp_1 _1380_ (.D(net64),
    .GATE(\genblk1[18].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[18][3] ));
 sky130_fd_sc_hd__dlxtp_1 _1381_ (.D(net55),
    .GATE(\genblk1[18].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[18][4] ));
 sky130_fd_sc_hd__dlxtp_1 _1382_ (.D(net47),
    .GATE(\genblk1[18].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[18][5] ));
 sky130_fd_sc_hd__dlxtp_1 _1383_ (.D(net38),
    .GATE(\genblk1[18].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[18][6] ));
 sky130_fd_sc_hd__dlxtp_1 _1384_ (.D(net29),
    .GATE(\genblk1[18].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[18][7] ));
 sky130_fd_sc_hd__dlxtp_1 _1385_ (.D(net91),
    .GATE(\genblk1[17].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[17][0] ));
 sky130_fd_sc_hd__dlxtp_1 _1386_ (.D(net80),
    .GATE(\genblk1[17].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[17][1] ));
 sky130_fd_sc_hd__dlxtp_1 _1387_ (.D(net73),
    .GATE(\genblk1[17].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[17][2] ));
 sky130_fd_sc_hd__dlxtp_1 _1388_ (.D(net64),
    .GATE(\genblk1[17].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[17][3] ));
 sky130_fd_sc_hd__dlxtp_1 _1389_ (.D(net56),
    .GATE(\genblk1[17].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[17][4] ));
 sky130_fd_sc_hd__dlxtp_1 _1390_ (.D(net47),
    .GATE(\genblk1[17].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[17][5] ));
 sky130_fd_sc_hd__dlxtp_1 _1391_ (.D(net39),
    .GATE(\genblk1[17].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[17][6] ));
 sky130_fd_sc_hd__dlxtp_1 _1392_ (.D(net29),
    .GATE(\genblk1[17].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[17][7] ));
 sky130_fd_sc_hd__dlxtp_1 _1393_ (.D(net88),
    .GATE(\genblk1[16].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[16][0] ));
 sky130_fd_sc_hd__dlxtp_1 _1394_ (.D(net79),
    .GATE(\genblk1[16].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[16][1] ));
 sky130_fd_sc_hd__dlxtp_1 _1395_ (.D(net71),
    .GATE(\genblk1[16].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[16][2] ));
 sky130_fd_sc_hd__dlxtp_1 _1396_ (.D(net65),
    .GATE(\genblk1[16].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[16][3] ));
 sky130_fd_sc_hd__dlxtp_1 _1397_ (.D(net55),
    .GATE(\genblk1[16].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[16][4] ));
 sky130_fd_sc_hd__dlxtp_1 _1398_ (.D(net47),
    .GATE(\genblk1[16].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[16][5] ));
 sky130_fd_sc_hd__dlxtp_1 _1399_ (.D(net38),
    .GATE(\genblk1[16].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[16][6] ));
 sky130_fd_sc_hd__dlxtp_1 _1400_ (.D(net30),
    .GATE(\genblk1[16].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[16][7] ));
 sky130_fd_sc_hd__dlxtp_1 _1401_ (.D(net89),
    .GATE(\genblk1[15].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[15][0] ));
 sky130_fd_sc_hd__dlxtp_1 _1402_ (.D(net82),
    .GATE(\genblk1[15].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[15][1] ));
 sky130_fd_sc_hd__dlxtp_1 _1403_ (.D(net76),
    .GATE(\genblk1[15].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[15][2] ));
 sky130_fd_sc_hd__dlxtp_1 _1404_ (.D(net66),
    .GATE(\genblk1[15].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[15][3] ));
 sky130_fd_sc_hd__dlxtp_1 _1405_ (.D(net57),
    .GATE(\genblk1[15].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[15][4] ));
 sky130_fd_sc_hd__dlxtp_1 _1406_ (.D(net50),
    .GATE(\genblk1[15].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[15][5] ));
 sky130_fd_sc_hd__dlxtp_1 _1407_ (.D(net40),
    .GATE(\genblk1[15].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[15][6] ));
 sky130_fd_sc_hd__dlxtp_1 _1408_ (.D(net36),
    .GATE(\genblk1[15].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[15][7] ));
 sky130_fd_sc_hd__dlxtp_1 _1409_ (.D(net89),
    .GATE(\genblk1[14].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[14][0] ));
 sky130_fd_sc_hd__dlxtp_1 _1410_ (.D(net82),
    .GATE(\genblk1[14].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[14][1] ));
 sky130_fd_sc_hd__dlxtp_1 _1411_ (.D(net76),
    .GATE(\genblk1[14].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[14][2] ));
 sky130_fd_sc_hd__dlxtp_1 _1412_ (.D(net66),
    .GATE(\genblk1[14].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[14][3] ));
 sky130_fd_sc_hd__dlxtp_1 _1413_ (.D(net57),
    .GATE(\genblk1[14].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[14][4] ));
 sky130_fd_sc_hd__dlxtp_1 _1414_ (.D(net50),
    .GATE(\genblk1[14].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[14][5] ));
 sky130_fd_sc_hd__dlxtp_1 _1415_ (.D(net40),
    .GATE(\genblk1[14].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[14][6] ));
 sky130_fd_sc_hd__dlxtp_1 _1416_ (.D(net36),
    .GATE(\genblk1[14].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[14][7] ));
 sky130_fd_sc_hd__dlxtp_1 _1417_ (.D(net90),
    .GATE(\genblk1[13].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[13][0] ));
 sky130_fd_sc_hd__dlxtp_1 _1418_ (.D(net81),
    .GATE(\genblk1[13].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[13][1] ));
 sky130_fd_sc_hd__dlxtp_1 _1419_ (.D(net76),
    .GATE(\genblk1[13].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[13][2] ));
 sky130_fd_sc_hd__dlxtp_1 _1420_ (.D(net66),
    .GATE(\genblk1[13].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[13][3] ));
 sky130_fd_sc_hd__dlxtp_1 _1421_ (.D(net58),
    .GATE(\genblk1[13].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[13][4] ));
 sky130_fd_sc_hd__dlxtp_1 _1422_ (.D(net51),
    .GATE(\genblk1[13].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[13][5] ));
 sky130_fd_sc_hd__dlxtp_1 _1423_ (.D(net41),
    .GATE(\genblk1[13].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[13][6] ));
 sky130_fd_sc_hd__dlxtp_1 _1424_ (.D(net36),
    .GATE(\genblk1[13].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[13][7] ));
 sky130_fd_sc_hd__dlxtp_1 _1425_ (.D(net90),
    .GATE(\genblk1[12].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[12][0] ));
 sky130_fd_sc_hd__dlxtp_1 _1426_ (.D(net81),
    .GATE(\genblk1[12].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[12][1] ));
 sky130_fd_sc_hd__dlxtp_1 _1427_ (.D(net76),
    .GATE(\genblk1[12].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[12][2] ));
 sky130_fd_sc_hd__dlxtp_1 _1428_ (.D(net65),
    .GATE(\genblk1[12].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[12][3] ));
 sky130_fd_sc_hd__dlxtp_1 _1429_ (.D(net57),
    .GATE(\genblk1[12].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[12][4] ));
 sky130_fd_sc_hd__dlxtp_1 _1430_ (.D(net51),
    .GATE(\genblk1[12].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[12][5] ));
 sky130_fd_sc_hd__dlxtp_1 _1431_ (.D(net40),
    .GATE(\genblk1[12].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[12][6] ));
 sky130_fd_sc_hd__dlxtp_1 _1432_ (.D(net31),
    .GATE(\genblk1[12].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[12][7] ));
 sky130_fd_sc_hd__dlxtp_1 _1433_ (.D(net90),
    .GATE(\genblk1[11].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[11][0] ));
 sky130_fd_sc_hd__dlxtp_1 _1434_ (.D(net82),
    .GATE(\genblk1[11].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[11][1] ));
 sky130_fd_sc_hd__dlxtp_1 _1435_ (.D(net75),
    .GATE(\genblk1[11].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[11][2] ));
 sky130_fd_sc_hd__dlxtp_1 _1436_ (.D(net66),
    .GATE(\genblk1[11].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[11][3] ));
 sky130_fd_sc_hd__dlxtp_1 _1437_ (.D(net58),
    .GATE(\genblk1[11].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[11][4] ));
 sky130_fd_sc_hd__dlxtp_1 _1438_ (.D(net50),
    .GATE(\genblk1[11].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[11][5] ));
 sky130_fd_sc_hd__dlxtp_1 _1439_ (.D(net41),
    .GATE(\genblk1[11].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[11][6] ));
 sky130_fd_sc_hd__dlxtp_1 _1440_ (.D(net31),
    .GATE(\genblk1[11].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[11][7] ));
 sky130_fd_sc_hd__dlxtp_1 _1441_ (.D(net91),
    .GATE(\genblk1[10].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[10][0] ));
 sky130_fd_sc_hd__dlxtp_1 _1442_ (.D(net82),
    .GATE(\genblk1[10].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[10][1] ));
 sky130_fd_sc_hd__dlxtp_1 _1443_ (.D(net75),
    .GATE(\genblk1[10].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[10][2] ));
 sky130_fd_sc_hd__dlxtp_1 _1444_ (.D(net65),
    .GATE(\genblk1[10].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[10][3] ));
 sky130_fd_sc_hd__dlxtp_1 _1445_ (.D(net57),
    .GATE(\genblk1[10].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[10][4] ));
 sky130_fd_sc_hd__dlxtp_1 _1446_ (.D(net50),
    .GATE(\genblk1[10].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[10][5] ));
 sky130_fd_sc_hd__dlxtp_1 _1447_ (.D(net40),
    .GATE(\genblk1[10].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[10][6] ));
 sky130_fd_sc_hd__dlxtp_1 _1448_ (.D(net31),
    .GATE(\genblk1[10].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[10][7] ));
 sky130_fd_sc_hd__dlxtp_1 _1449_ (.D(net90),
    .GATE(\genblk1[9].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[9][0] ));
 sky130_fd_sc_hd__dlxtp_1 _1450_ (.D(net81),
    .GATE(\genblk1[9].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[9][1] ));
 sky130_fd_sc_hd__dlxtp_1 _1451_ (.D(net75),
    .GATE(\genblk1[9].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[9][2] ));
 sky130_fd_sc_hd__dlxtp_1 _1452_ (.D(net65),
    .GATE(\genblk1[9].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[9][3] ));
 sky130_fd_sc_hd__dlxtp_1 _1453_ (.D(net57),
    .GATE(\genblk1[9].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[9][4] ));
 sky130_fd_sc_hd__dlxtp_1 _1454_ (.D(net51),
    .GATE(\genblk1[9].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[9][5] ));
 sky130_fd_sc_hd__dlxtp_1 _1455_ (.D(net41),
    .GATE(\genblk1[9].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[9][6] ));
 sky130_fd_sc_hd__dlxtp_1 _1456_ (.D(net32),
    .GATE(\genblk1[9].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[9][7] ));
 sky130_fd_sc_hd__dlxtp_1 _1457_ (.D(net89),
    .GATE(\genblk1[8].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[8][0] ));
 sky130_fd_sc_hd__dlxtp_1 _1458_ (.D(net81),
    .GATE(\genblk1[8].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[8][1] ));
 sky130_fd_sc_hd__dlxtp_1 _1459_ (.D(net75),
    .GATE(\genblk1[8].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[8][2] ));
 sky130_fd_sc_hd__dlxtp_1 _1460_ (.D(net66),
    .GATE(\genblk1[8].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[8][3] ));
 sky130_fd_sc_hd__dlxtp_1 _1461_ (.D(net57),
    .GATE(\genblk1[8].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[8][4] ));
 sky130_fd_sc_hd__dlxtp_1 _1462_ (.D(net51),
    .GATE(\genblk1[8].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[8][5] ));
 sky130_fd_sc_hd__dlxtp_1 _1463_ (.D(net40),
    .GATE(\genblk1[8].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[8][6] ));
 sky130_fd_sc_hd__dlxtp_1 _1464_ (.D(net31),
    .GATE(\genblk1[8].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[8][7] ));
 sky130_fd_sc_hd__dlxtp_1 _1465_ (.D(net89),
    .GATE(\genblk1[7].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[7][0] ));
 sky130_fd_sc_hd__dlxtp_1 _1466_ (.D(net81),
    .GATE(\genblk1[7].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[7][1] ));
 sky130_fd_sc_hd__dlxtp_1 _1467_ (.D(net75),
    .GATE(\genblk1[7].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[7][2] ));
 sky130_fd_sc_hd__dlxtp_1 _1468_ (.D(net65),
    .GATE(\genblk1[7].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[7][3] ));
 sky130_fd_sc_hd__dlxtp_1 _1469_ (.D(net58),
    .GATE(\genblk1[7].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[7][4] ));
 sky130_fd_sc_hd__dlxtp_1 _1470_ (.D(net51),
    .GATE(\genblk1[7].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[7][5] ));
 sky130_fd_sc_hd__dlxtp_1 _1471_ (.D(net41),
    .GATE(\genblk1[7].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[7][6] ));
 sky130_fd_sc_hd__dlxtp_1 _1472_ (.D(net31),
    .GATE(\genblk1[7].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[7][7] ));
 sky130_fd_sc_hd__dlxtp_1 _1473_ (.D(net89),
    .GATE(\genblk1[6].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[6][0] ));
 sky130_fd_sc_hd__dlxtp_1 _1474_ (.D(net82),
    .GATE(\genblk1[6].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[6][1] ));
 sky130_fd_sc_hd__dlxtp_1 _1475_ (.D(net76),
    .GATE(\genblk1[6].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[6][2] ));
 sky130_fd_sc_hd__dlxtp_1 _1476_ (.D(net66),
    .GATE(\genblk1[6].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[6][3] ));
 sky130_fd_sc_hd__dlxtp_1 _1477_ (.D(net58),
    .GATE(\genblk1[6].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[6][4] ));
 sky130_fd_sc_hd__dlxtp_1 _1478_ (.D(net50),
    .GATE(\genblk1[6].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[6][5] ));
 sky130_fd_sc_hd__dlxtp_1 _1479_ (.D(net41),
    .GATE(\genblk1[6].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[6][6] ));
 sky130_fd_sc_hd__dlxtp_1 _1480_ (.D(net36),
    .GATE(\genblk1[6].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[6][7] ));
 sky130_fd_sc_hd__dlxtp_1 _1481_ (.D(net89),
    .GATE(\genblk1[5].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[5][0] ));
 sky130_fd_sc_hd__dlxtp_1 _1482_ (.D(net81),
    .GATE(\genblk1[5].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[5][1] ));
 sky130_fd_sc_hd__dlxtp_1 _1483_ (.D(net76),
    .GATE(\genblk1[5].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[5][2] ));
 sky130_fd_sc_hd__dlxtp_1 _1484_ (.D(net66),
    .GATE(\genblk1[5].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[5][3] ));
 sky130_fd_sc_hd__dlxtp_1 _1485_ (.D(net57),
    .GATE(\genblk1[5].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[5][4] ));
 sky130_fd_sc_hd__dlxtp_1 _1486_ (.D(net50),
    .GATE(\genblk1[5].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[5][5] ));
 sky130_fd_sc_hd__dlxtp_1 _1487_ (.D(net40),
    .GATE(\genblk1[5].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[5][6] ));
 sky130_fd_sc_hd__dlxtp_1 _1488_ (.D(net31),
    .GATE(\genblk1[5].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[5][7] ));
 sky130_fd_sc_hd__dlxtp_1 _1489_ (.D(net89),
    .GATE(\genblk1[4].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[4][0] ));
 sky130_fd_sc_hd__dlxtp_1 _1490_ (.D(net81),
    .GATE(\genblk1[4].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[4][1] ));
 sky130_fd_sc_hd__dlxtp_1 _1491_ (.D(net75),
    .GATE(\genblk1[4].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[4][2] ));
 sky130_fd_sc_hd__dlxtp_1 _1492_ (.D(net65),
    .GATE(\genblk1[4].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[4][3] ));
 sky130_fd_sc_hd__dlxtp_1 _1493_ (.D(net58),
    .GATE(\genblk1[4].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[4][4] ));
 sky130_fd_sc_hd__dlxtp_1 _1494_ (.D(net51),
    .GATE(\genblk1[4].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[4][5] ));
 sky130_fd_sc_hd__dlxtp_1 _1495_ (.D(net41),
    .GATE(\genblk1[4].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[4][6] ));
 sky130_fd_sc_hd__dlxtp_1 _1496_ (.D(net32),
    .GATE(\genblk1[4].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[4][7] ));
 sky130_fd_sc_hd__dlxtp_1 _1497_ (.D(net89),
    .GATE(\genblk1[3].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[3][0] ));
 sky130_fd_sc_hd__dlxtp_1 _1498_ (.D(net81),
    .GATE(\genblk1[3].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[3][1] ));
 sky130_fd_sc_hd__dlxtp_1 _1499_ (.D(net75),
    .GATE(\genblk1[3].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[3][2] ));
 sky130_fd_sc_hd__dlxtp_1 _1500_ (.D(net66),
    .GATE(\genblk1[3].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[3][3] ));
 sky130_fd_sc_hd__dlxtp_1 _1501_ (.D(net57),
    .GATE(\genblk1[3].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[3][4] ));
 sky130_fd_sc_hd__dlxtp_1 _1502_ (.D(net51),
    .GATE(\genblk1[3].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[3][5] ));
 sky130_fd_sc_hd__dlxtp_1 _1503_ (.D(net40),
    .GATE(\genblk1[3].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[3][6] ));
 sky130_fd_sc_hd__dlxtp_1 _1504_ (.D(net36),
    .GATE(\genblk1[3].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[3][7] ));
 sky130_fd_sc_hd__dlxtp_1 _1505_ (.D(net89),
    .GATE(\genblk1[2].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[2][0] ));
 sky130_fd_sc_hd__dlxtp_1 _1506_ (.D(net81),
    .GATE(\genblk1[2].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[2][1] ));
 sky130_fd_sc_hd__dlxtp_1 _1507_ (.D(net75),
    .GATE(\genblk1[2].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[2][2] ));
 sky130_fd_sc_hd__dlxtp_1 _1508_ (.D(net66),
    .GATE(\genblk1[2].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[2][3] ));
 sky130_fd_sc_hd__dlxtp_1 _1509_ (.D(net57),
    .GATE(\genblk1[2].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[2][4] ));
 sky130_fd_sc_hd__dlxtp_1 _1510_ (.D(net51),
    .GATE(\genblk1[2].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[2][5] ));
 sky130_fd_sc_hd__dlxtp_1 _1511_ (.D(net40),
    .GATE(\genblk1[2].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[2][6] ));
 sky130_fd_sc_hd__dlxtp_1 _1512_ (.D(net32),
    .GATE(\genblk1[2].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[2][7] ));
 sky130_fd_sc_hd__dlxtp_1 _1513_ (.D(net90),
    .GATE(\genblk1[1].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[1][0] ));
 sky130_fd_sc_hd__dlxtp_1 _1514_ (.D(net81),
    .GATE(\genblk1[1].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[1][1] ));
 sky130_fd_sc_hd__dlxtp_1 _1515_ (.D(net75),
    .GATE(\genblk1[1].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[1][2] ));
 sky130_fd_sc_hd__dlxtp_1 _1516_ (.D(net65),
    .GATE(\genblk1[1].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[1][3] ));
 sky130_fd_sc_hd__dlxtp_1 _1517_ (.D(net57),
    .GATE(\genblk1[1].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[1][4] ));
 sky130_fd_sc_hd__dlxtp_1 _1518_ (.D(net51),
    .GATE(\genblk1[1].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[1][5] ));
 sky130_fd_sc_hd__dlxtp_1 _1519_ (.D(net41),
    .GATE(\genblk1[1].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[1][6] ));
 sky130_fd_sc_hd__dlxtp_1 _1520_ (.D(net36),
    .GATE(\genblk1[1].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[1][7] ));
 sky130_fd_sc_hd__dlxtp_1 _1521_ (.D(net89),
    .GATE(\genblk1[0].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[0][0] ));
 sky130_fd_sc_hd__dlxtp_1 _1522_ (.D(net82),
    .GATE(\genblk1[0].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[0][1] ));
 sky130_fd_sc_hd__dlxtp_1 _1523_ (.D(net75),
    .GATE(\genblk1[0].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[0][2] ));
 sky130_fd_sc_hd__dlxtp_1 _1524_ (.D(net67),
    .GATE(\genblk1[0].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[0][3] ));
 sky130_fd_sc_hd__dlxtp_1 _1525_ (.D(net58),
    .GATE(\genblk1[0].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[0][4] ));
 sky130_fd_sc_hd__dlxtp_1 _1526_ (.D(\data_to_write[5] ),
    .GATE(\genblk1[0].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[0][5] ));
 sky130_fd_sc_hd__dlxtp_1 _1527_ (.D(net41),
    .GATE(\genblk1[0].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[0][6] ));
 sky130_fd_sc_hd__dlxtp_1 _1528_ (.D(net36),
    .GATE(\genblk1[0].wr_en_this_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RAM[0][7] ));
 sky130_fd_sc_hd__dfxtp_4 _1529_ (.CLK(clknet_1_1__leaf_clk),
    .D(_0003_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk2[3].partition_sel_n ));
 sky130_fd_sc_hd__dfxtp_4 _1530_ (.CLK(clknet_1_0__leaf_clk),
    .D(_0002_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk2[2].partition_sel_n ));
 sky130_fd_sc_hd__dfxtp_4 _1531_ (.CLK(clknet_1_0__leaf_clk),
    .D(_0001_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk2[1].partition_sel_n ));
 sky130_fd_sc_hd__dfxtp_4 _1532_ (.CLK(clknet_1_0__leaf_clk),
    .D(_0000_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk2[0].partition_sel_n ));
 sky130_fd_sc_hd__dfxtp_1 _1533_ (.CLK(net112),
    .D(_0004_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(wr_en_ok));
 sky130_fd_sc_hd__dfxtp_2 _1534_ (.CLK(clknet_1_1__leaf_clk),
    .D(net2),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\addr_read[0] ));
 sky130_fd_sc_hd__dfxtp_2 _1535_ (.CLK(clknet_1_1__leaf_clk),
    .D(net3),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\addr_read[1] ));
 sky130_fd_sc_hd__dfxtp_2 _1536_ (.CLK(clknet_1_1__leaf_clk),
    .D(net4),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\addr_read[2] ));
 sky130_fd_sc_hd__dfxtp_2 _1537_ (.CLK(clknet_1_1__leaf_clk),
    .D(net5),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\addr_read[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1538_ (.CLK(clknet_1_1__leaf_clk),
    .D(_0014_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\addr_write[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1539_ (.CLK(clknet_1_1__leaf_clk),
    .D(_0015_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\addr_write[1] ));
 sky130_fd_sc_hd__dfxtp_2 _1540_ (.CLK(clknet_1_1__leaf_clk),
    .D(_0016_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\addr_write[2] ));
 sky130_fd_sc_hd__dfxtp_2 _1541_ (.CLK(clknet_1_1__leaf_clk),
    .D(_0017_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\addr_write[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1542_ (.CLK(clknet_1_1__leaf_clk),
    .D(_0018_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\addr_write[4] ));
 sky130_fd_sc_hd__dfxtp_1 _1543_ (.CLK(clknet_1_0__leaf_clk),
    .D(_0019_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\addr_write[5] ));
 sky130_fd_sc_hd__dfxtp_1 _1544_ (.CLK(clknet_1_1__leaf_clk),
    .D(_0020_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(wr_en_next));
 sky130_fd_sc_hd__dfxtp_1 _1545_ (.CLK(clknet_1_1__leaf_clk),
    .D(_0021_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(wr_en_valid));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_2 fanout17 (.A(net18),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_2 fanout18 (.A(net19),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_2 fanout19 (.A(net24),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_2 fanout20 (.A(net21),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net20));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout21 (.A(net24),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_2 fanout22 (.A(net23),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net22));
 sky130_fd_sc_hd__buf_2 fanout23 (.A(net24),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_2 fanout24 (.A(wr_en),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_2 fanout29 (.A(net30),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_2 fanout30 (.A(net32),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net30));
 sky130_fd_sc_hd__buf_2 fanout31 (.A(net32),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_2 fanout32 (.A(net37),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net32));
 sky130_fd_sc_hd__buf_2 fanout33 (.A(net35),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_2 fanout34 (.A(net35),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_2 fanout35 (.A(net37),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net35));
 sky130_fd_sc_hd__buf_2 fanout36 (.A(net37),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_2 fanout37 (.A(\data_to_write[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net37));
 sky130_fd_sc_hd__buf_2 fanout38 (.A(net39),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net38));
 sky130_fd_sc_hd__buf_1 fanout39 (.A(\data_to_write[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net39));
 sky130_fd_sc_hd__buf_2 fanout40 (.A(net41),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_2 fanout41 (.A(\data_to_write[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_2 fanout42 (.A(net46),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net42));
 sky130_fd_sc_hd__buf_1 fanout43 (.A(net46),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_2 fanout44 (.A(net46),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net44));
 sky130_fd_sc_hd__buf_1 fanout45 (.A(net46),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_2 fanout46 (.A(\data_to_write[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net46));
 sky130_fd_sc_hd__buf_2 fanout47 (.A(net49),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net47));
 sky130_fd_sc_hd__buf_2 fanout48 (.A(net49),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_2 fanout49 (.A(\data_to_write[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net49));
 sky130_fd_sc_hd__buf_2 fanout50 (.A(net51),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net50));
 sky130_fd_sc_hd__buf_2 fanout51 (.A(\data_to_write[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_2 fanout52 (.A(net53),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_2 fanout53 (.A(net54),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net53));
 sky130_fd_sc_hd__buf_2 fanout54 (.A(\data_to_write[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net54));
 sky130_fd_sc_hd__buf_2 fanout55 (.A(net56),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net55));
 sky130_fd_sc_hd__clkbuf_2 fanout56 (.A(\data_to_write[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net56));
 sky130_fd_sc_hd__buf_2 fanout57 (.A(net58),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net57));
 sky130_fd_sc_hd__clkbuf_2 fanout58 (.A(\data_to_write[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net58));
 sky130_fd_sc_hd__clkbuf_2 fanout59 (.A(net61),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net59));
 sky130_fd_sc_hd__buf_1 fanout60 (.A(net62),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net60));
 sky130_fd_sc_hd__buf_2 fanout61 (.A(net62),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net61));
 sky130_fd_sc_hd__buf_2 fanout62 (.A(\data_to_write[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net62));
 sky130_fd_sc_hd__buf_2 fanout63 (.A(net64),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net63));
 sky130_fd_sc_hd__buf_2 fanout64 (.A(net70),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net64));
 sky130_fd_sc_hd__clkbuf_2 fanout65 (.A(net66),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net65));
 sky130_fd_sc_hd__buf_2 fanout66 (.A(net67),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net66));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout67 (.A(net70),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net67));
 sky130_fd_sc_hd__buf_2 fanout68 (.A(net69),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net68));
 sky130_fd_sc_hd__buf_2 fanout69 (.A(net70),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net69));
 sky130_fd_sc_hd__buf_2 fanout70 (.A(\data_to_write[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net70));
 sky130_fd_sc_hd__clkbuf_2 fanout71 (.A(net72),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net71));
 sky130_fd_sc_hd__buf_2 fanout72 (.A(net73),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net72));
 sky130_fd_sc_hd__buf_2 fanout73 (.A(net74),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net73));
 sky130_fd_sc_hd__buf_1 fanout74 (.A(\data_to_write[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net74));
 sky130_fd_sc_hd__clkbuf_2 fanout75 (.A(\data_to_write[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net75));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout76 (.A(\data_to_write[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net76));
 sky130_fd_sc_hd__clkbuf_2 fanout77 (.A(net78),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net77));
 sky130_fd_sc_hd__clkbuf_2 fanout78 (.A(\data_to_write[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net78));
 sky130_fd_sc_hd__buf_2 fanout79 (.A(net83),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net79));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout80 (.A(net83),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net80));
 sky130_fd_sc_hd__buf_2 fanout81 (.A(net83),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net81));
 sky130_fd_sc_hd__clkbuf_2 fanout82 (.A(net83),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net82));
 sky130_fd_sc_hd__buf_2 fanout83 (.A(\data_to_write[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net83));
 sky130_fd_sc_hd__clkbuf_2 fanout84 (.A(net86),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net84));
 sky130_fd_sc_hd__buf_2 fanout85 (.A(net86),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net85));
 sky130_fd_sc_hd__buf_2 fanout86 (.A(net87),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net86));
 sky130_fd_sc_hd__clkbuf_2 fanout87 (.A(\data_to_write[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net87));
 sky130_fd_sc_hd__buf_2 fanout88 (.A(net91),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net88));
 sky130_fd_sc_hd__buf_2 fanout89 (.A(net90),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net89));
 sky130_fd_sc_hd__buf_2 fanout90 (.A(net91),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net90));
 sky130_fd_sc_hd__clkbuf_2 fanout91 (.A(\data_to_write[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net91));
 sky130_fd_sc_hd__clkbuf_2 fanout92 (.A(net94),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net92));
 sky130_fd_sc_hd__buf_2 fanout93 (.A(net94),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net93));
 sky130_fd_sc_hd__clkbuf_2 fanout94 (.A(net95),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net94));
 sky130_fd_sc_hd__buf_2 fanout95 (.A(\data_to_write[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net95));
 sky130_fd_sc_hd__and2_2 \genblk1[0].lm_gate  (.A(net21),
    .B(\genblk1[0].sel_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[0].wr_en_this_byte ));
 sky130_fd_sc_hd__and2_2 \genblk1[10].lm_gate  (.A(net20),
    .B(\genblk1[10].sel_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[10].wr_en_this_byte ));
 sky130_fd_sc_hd__and2_2 \genblk1[11].lm_gate  (.A(net20),
    .B(\genblk1[11].sel_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[11].wr_en_this_byte ));
 sky130_fd_sc_hd__and2_2 \genblk1[12].lm_gate  (.A(net20),
    .B(\genblk1[12].sel_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[12].wr_en_this_byte ));
 sky130_fd_sc_hd__and2_2 \genblk1[13].lm_gate  (.A(net20),
    .B(\genblk1[13].sel_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[13].wr_en_this_byte ));
 sky130_fd_sc_hd__and2_2 \genblk1[14].lm_gate  (.A(net21),
    .B(\genblk1[14].sel_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[14].wr_en_this_byte ));
 sky130_fd_sc_hd__and2_2 \genblk1[15].lm_gate  (.A(net22),
    .B(\genblk1[15].sel_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[15].wr_en_this_byte ));
 sky130_fd_sc_hd__and2_2 \genblk1[16].lm_gate  (.A(net19),
    .B(\genblk1[16].sel_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[16].wr_en_this_byte ));
 sky130_fd_sc_hd__and2_2 \genblk1[17].lm_gate  (.A(net17),
    .B(\genblk1[17].sel_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[17].wr_en_this_byte ));
 sky130_fd_sc_hd__and2_2 \genblk1[18].lm_gate  (.A(net17),
    .B(\genblk1[18].sel_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[18].wr_en_this_byte ));
 sky130_fd_sc_hd__and2_2 \genblk1[19].lm_gate  (.A(net18),
    .B(\genblk1[19].sel_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[19].wr_en_this_byte ));
 sky130_fd_sc_hd__and2_2 \genblk1[1].lm_gate  (.A(net21),
    .B(\genblk1[1].sel_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[1].wr_en_this_byte ));
 sky130_fd_sc_hd__and2_2 \genblk1[20].lm_gate  (.A(net17),
    .B(\genblk1[20].sel_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[20].wr_en_this_byte ));
 sky130_fd_sc_hd__and2_2 \genblk1[21].lm_gate  (.A(net18),
    .B(\genblk1[21].sel_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[21].wr_en_this_byte ));
 sky130_fd_sc_hd__and2_2 \genblk1[22].lm_gate  (.A(net17),
    .B(\genblk1[22].sel_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[22].wr_en_this_byte ));
 sky130_fd_sc_hd__and2_2 \genblk1[23].lm_gate  (.A(net17),
    .B(\genblk1[23].sel_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[23].wr_en_this_byte ));
 sky130_fd_sc_hd__and2_2 \genblk1[24].lm_gate  (.A(net17),
    .B(\genblk1[24].sel_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[24].wr_en_this_byte ));
 sky130_fd_sc_hd__and2_2 \genblk1[25].lm_gate  (.A(net17),
    .B(\genblk1[25].sel_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[25].wr_en_this_byte ));
 sky130_fd_sc_hd__and2_2 \genblk1[26].lm_gate  (.A(net18),
    .B(\genblk1[26].sel_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[26].wr_en_this_byte ));
 sky130_fd_sc_hd__and2_2 \genblk1[27].lm_gate  (.A(net19),
    .B(\genblk1[27].sel_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[27].wr_en_this_byte ));
 sky130_fd_sc_hd__and2_2 \genblk1[28].lm_gate  (.A(net18),
    .B(\genblk1[28].sel_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[28].wr_en_this_byte ));
 sky130_fd_sc_hd__and2_2 \genblk1[29].lm_gate  (.A(net19),
    .B(\genblk1[29].sel_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[29].wr_en_this_byte ));
 sky130_fd_sc_hd__and2_2 \genblk1[2].lm_gate  (.A(net20),
    .B(\genblk1[2].sel_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[2].wr_en_this_byte ));
 sky130_fd_sc_hd__and2_2 \genblk1[30].lm_gate  (.A(net19),
    .B(\genblk1[30].sel_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[30].wr_en_this_byte ));
 sky130_fd_sc_hd__and2_2 \genblk1[31].lm_gate  (.A(net20),
    .B(\genblk1[31].sel_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[31].wr_en_this_byte ));
 sky130_fd_sc_hd__and2_2 \genblk1[32].lm_gate  (.A(net18),
    .B(\genblk1[32].sel_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[32].wr_en_this_byte ));
 sky130_fd_sc_hd__and2_2 \genblk1[33].lm_gate  (.A(net19),
    .B(\genblk1[33].sel_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[33].wr_en_this_byte ));
 sky130_fd_sc_hd__and2_2 \genblk1[34].lm_gate  (.A(net17),
    .B(\genblk1[34].sel_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[34].wr_en_this_byte ));
 sky130_fd_sc_hd__and2_2 \genblk1[35].lm_gate  (.A(net18),
    .B(\genblk1[35].sel_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[35].wr_en_this_byte ));
 sky130_fd_sc_hd__and2_2 \genblk1[36].lm_gate  (.A(net17),
    .B(\genblk1[36].sel_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[36].wr_en_this_byte ));
 sky130_fd_sc_hd__and2_2 \genblk1[37].lm_gate  (.A(net19),
    .B(\genblk1[37].sel_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[37].wr_en_this_byte ));
 sky130_fd_sc_hd__and2_2 \genblk1[38].lm_gate  (.A(net17),
    .B(\genblk1[38].sel_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[38].wr_en_this_byte ));
 sky130_fd_sc_hd__and2_2 \genblk1[39].lm_gate  (.A(net18),
    .B(\genblk1[39].sel_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[39].wr_en_this_byte ));
 sky130_fd_sc_hd__and2_2 \genblk1[3].lm_gate  (.A(net21),
    .B(\genblk1[3].sel_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[3].wr_en_this_byte ));
 sky130_fd_sc_hd__and2_2 \genblk1[40].lm_gate  (.A(net18),
    .B(\genblk1[40].sel_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[40].wr_en_this_byte ));
 sky130_fd_sc_hd__and2_2 \genblk1[41].lm_gate  (.A(net18),
    .B(\genblk1[41].sel_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[41].wr_en_this_byte ));
 sky130_fd_sc_hd__and2_2 \genblk1[42].lm_gate  (.A(net19),
    .B(\genblk1[42].sel_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[42].wr_en_this_byte ));
 sky130_fd_sc_hd__and2_2 \genblk1[43].lm_gate  (.A(net22),
    .B(\genblk1[43].sel_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[43].wr_en_this_byte ));
 sky130_fd_sc_hd__and2_2 \genblk1[44].lm_gate  (.A(net23),
    .B(\genblk1[44].sel_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[44].wr_en_this_byte ));
 sky130_fd_sc_hd__and2_2 \genblk1[45].lm_gate  (.A(net23),
    .B(\genblk1[45].sel_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[45].wr_en_this_byte ));
 sky130_fd_sc_hd__and2_2 \genblk1[46].lm_gate  (.A(net23),
    .B(\genblk1[46].sel_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[46].wr_en_this_byte ));
 sky130_fd_sc_hd__and2_2 \genblk1[47].lm_gate  (.A(net22),
    .B(\genblk1[47].sel_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[47].wr_en_this_byte ));
 sky130_fd_sc_hd__and2_2 \genblk1[48].lm_gate  (.A(net23),
    .B(\genblk1[48].sel_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[48].wr_en_this_byte ));
 sky130_fd_sc_hd__and2_2 \genblk1[49].lm_gate  (.A(net23),
    .B(\genblk1[49].sel_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[49].wr_en_this_byte ));
 sky130_fd_sc_hd__and2_2 \genblk1[4].lm_gate  (.A(net20),
    .B(\genblk1[4].sel_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[4].wr_en_this_byte ));
 sky130_fd_sc_hd__and2_2 \genblk1[50].lm_gate  (.A(net23),
    .B(\genblk1[50].sel_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[50].wr_en_this_byte ));
 sky130_fd_sc_hd__and2_2 \genblk1[51].lm_gate  (.A(net24),
    .B(\genblk1[51].sel_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[51].wr_en_this_byte ));
 sky130_fd_sc_hd__and2_2 \genblk1[52].lm_gate  (.A(net22),
    .B(\genblk1[52].sel_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[52].wr_en_this_byte ));
 sky130_fd_sc_hd__and2_2 \genblk1[53].lm_gate  (.A(net23),
    .B(\genblk1[53].sel_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[53].wr_en_this_byte ));
 sky130_fd_sc_hd__and2_2 \genblk1[54].lm_gate  (.A(net22),
    .B(\genblk1[54].sel_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[54].wr_en_this_byte ));
 sky130_fd_sc_hd__and2_2 \genblk1[55].lm_gate  (.A(net23),
    .B(\genblk1[55].sel_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[55].wr_en_this_byte ));
 sky130_fd_sc_hd__and2_2 \genblk1[56].lm_gate  (.A(net22),
    .B(\genblk1[56].sel_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[56].wr_en_this_byte ));
 sky130_fd_sc_hd__and2_2 \genblk1[57].lm_gate  (.A(net22),
    .B(\genblk1[57].sel_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[57].wr_en_this_byte ));
 sky130_fd_sc_hd__and2_2 \genblk1[58].lm_gate  (.A(net22),
    .B(\genblk1[58].sel_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[58].wr_en_this_byte ));
 sky130_fd_sc_hd__and2_2 \genblk1[59].lm_gate  (.A(net22),
    .B(\genblk1[59].sel_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[59].wr_en_this_byte ));
 sky130_fd_sc_hd__and2_2 \genblk1[5].lm_gate  (.A(net21),
    .B(\genblk1[5].sel_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[5].wr_en_this_byte ));
 sky130_fd_sc_hd__and2_2 \genblk1[60].lm_gate  (.A(net24),
    .B(\genblk1[60].sel_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[60].wr_en_this_byte ));
 sky130_fd_sc_hd__and2_2 \genblk1[61].lm_gate  (.A(net22),
    .B(\genblk1[61].sel_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[61].wr_en_this_byte ));
 sky130_fd_sc_hd__and2_2 \genblk1[62].lm_gate  (.A(net24),
    .B(\genblk1[62].sel_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[62].wr_en_this_byte ));
 sky130_fd_sc_hd__and2_2 \genblk1[63].lm_gate  (.A(net23),
    .B(\genblk1[63].sel_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[63].wr_en_this_byte ));
 sky130_fd_sc_hd__and2_2 \genblk1[6].lm_gate  (.A(net20),
    .B(\genblk1[6].sel_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[6].wr_en_this_byte ));
 sky130_fd_sc_hd__and2_2 \genblk1[7].lm_gate  (.A(net20),
    .B(\genblk1[7].sel_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[7].wr_en_this_byte ));
 sky130_fd_sc_hd__and2_2 \genblk1[8].lm_gate  (.A(net21),
    .B(\genblk1[8].sel_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[8].wr_en_this_byte ));
 sky130_fd_sc_hd__and2_2 \genblk1[9].lm_gate  (.A(net20),
    .B(\genblk1[9].sel_byte ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[9].wr_en_this_byte ));
 sky130_fd_sc_hd__ebufn_4 \genblk2[0].lm_dt_out_buf[0]  (.A(\genblk2[0].selected_out[0] ),
    .TE_B(\genblk2[0].partition_sel_n ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\combined_out[0] ));
 sky130_fd_sc_hd__ebufn_4 \genblk2[0].lm_dt_out_buf[1]  (.A(\genblk2[0].selected_out[1] ),
    .TE_B(\genblk2[0].partition_sel_n ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\combined_out[1] ));
 sky130_fd_sc_hd__ebufn_4 \genblk2[0].lm_dt_out_buf[2]  (.A(\genblk2[0].selected_out[2] ),
    .TE_B(\genblk2[0].partition_sel_n ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\combined_out[2] ));
 sky130_fd_sc_hd__ebufn_4 \genblk2[0].lm_dt_out_buf[3]  (.A(\genblk2[0].selected_out[3] ),
    .TE_B(\genblk2[0].partition_sel_n ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\combined_out[3] ));
 sky130_fd_sc_hd__ebufn_4 \genblk2[0].lm_dt_out_buf[4]  (.A(\genblk2[0].selected_out[4] ),
    .TE_B(\genblk2[0].partition_sel_n ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\combined_out[4] ));
 sky130_fd_sc_hd__ebufn_4 \genblk2[0].lm_dt_out_buf[5]  (.A(\genblk2[0].selected_out[5] ),
    .TE_B(\genblk2[0].partition_sel_n ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\combined_out[5] ));
 sky130_fd_sc_hd__ebufn_4 \genblk2[0].lm_dt_out_buf[6]  (.A(\genblk2[0].selected_out[6] ),
    .TE_B(\genblk2[0].partition_sel_n ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\combined_out[6] ));
 sky130_fd_sc_hd__ebufn_4 \genblk2[0].lm_dt_out_buf[7]  (.A(\genblk2[0].selected_out[7] ),
    .TE_B(\genblk2[0].partition_sel_n ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\combined_out[7] ));
 sky130_fd_sc_hd__ebufn_4 \genblk2[1].lm_dt_out_buf[0]  (.A(\genblk2[1].selected_out[0] ),
    .TE_B(\genblk2[1].partition_sel_n ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\combined_out[0] ));
 sky130_fd_sc_hd__ebufn_4 \genblk2[1].lm_dt_out_buf[1]  (.A(\genblk2[1].selected_out[1] ),
    .TE_B(\genblk2[1].partition_sel_n ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\combined_out[1] ));
 sky130_fd_sc_hd__ebufn_4 \genblk2[1].lm_dt_out_buf[2]  (.A(\genblk2[1].selected_out[2] ),
    .TE_B(\genblk2[1].partition_sel_n ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\combined_out[2] ));
 sky130_fd_sc_hd__ebufn_4 \genblk2[1].lm_dt_out_buf[3]  (.A(\genblk2[1].selected_out[3] ),
    .TE_B(\genblk2[1].partition_sel_n ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\combined_out[3] ));
 sky130_fd_sc_hd__ebufn_4 \genblk2[1].lm_dt_out_buf[4]  (.A(\genblk2[1].selected_out[4] ),
    .TE_B(\genblk2[1].partition_sel_n ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\combined_out[4] ));
 sky130_fd_sc_hd__ebufn_4 \genblk2[1].lm_dt_out_buf[5]  (.A(\genblk2[1].selected_out[5] ),
    .TE_B(\genblk2[1].partition_sel_n ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\combined_out[5] ));
 sky130_fd_sc_hd__ebufn_4 \genblk2[1].lm_dt_out_buf[6]  (.A(\genblk2[1].selected_out[6] ),
    .TE_B(\genblk2[1].partition_sel_n ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\combined_out[6] ));
 sky130_fd_sc_hd__ebufn_4 \genblk2[1].lm_dt_out_buf[7]  (.A(\genblk2[1].selected_out[7] ),
    .TE_B(\genblk2[1].partition_sel_n ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\combined_out[7] ));
 sky130_fd_sc_hd__ebufn_4 \genblk2[2].lm_dt_out_buf[0]  (.A(\genblk2[2].selected_out[0] ),
    .TE_B(\genblk2[2].partition_sel_n ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\combined_out[0] ));
 sky130_fd_sc_hd__ebufn_4 \genblk2[2].lm_dt_out_buf[1]  (.A(\genblk2[2].selected_out[1] ),
    .TE_B(\genblk2[2].partition_sel_n ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\combined_out[1] ));
 sky130_fd_sc_hd__ebufn_4 \genblk2[2].lm_dt_out_buf[2]  (.A(\genblk2[2].selected_out[2] ),
    .TE_B(\genblk2[2].partition_sel_n ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\combined_out[2] ));
 sky130_fd_sc_hd__ebufn_4 \genblk2[2].lm_dt_out_buf[3]  (.A(\genblk2[2].selected_out[3] ),
    .TE_B(\genblk2[2].partition_sel_n ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\combined_out[3] ));
 sky130_fd_sc_hd__ebufn_4 \genblk2[2].lm_dt_out_buf[4]  (.A(\genblk2[2].selected_out[4] ),
    .TE_B(\genblk2[2].partition_sel_n ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\combined_out[4] ));
 sky130_fd_sc_hd__ebufn_4 \genblk2[2].lm_dt_out_buf[5]  (.A(\genblk2[2].selected_out[5] ),
    .TE_B(\genblk2[2].partition_sel_n ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\combined_out[5] ));
 sky130_fd_sc_hd__ebufn_4 \genblk2[2].lm_dt_out_buf[6]  (.A(\genblk2[2].selected_out[6] ),
    .TE_B(\genblk2[2].partition_sel_n ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\combined_out[6] ));
 sky130_fd_sc_hd__ebufn_4 \genblk2[2].lm_dt_out_buf[7]  (.A(\genblk2[2].selected_out[7] ),
    .TE_B(\genblk2[2].partition_sel_n ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\combined_out[7] ));
 sky130_fd_sc_hd__ebufn_4 \genblk2[3].lm_dt_out_buf[0]  (.A(\genblk2[3].selected_out[0] ),
    .TE_B(\genblk2[3].partition_sel_n ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\combined_out[0] ));
 sky130_fd_sc_hd__ebufn_4 \genblk2[3].lm_dt_out_buf[1]  (.A(\genblk2[3].selected_out[1] ),
    .TE_B(\genblk2[3].partition_sel_n ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\combined_out[1] ));
 sky130_fd_sc_hd__ebufn_4 \genblk2[3].lm_dt_out_buf[2]  (.A(\genblk2[3].selected_out[2] ),
    .TE_B(\genblk2[3].partition_sel_n ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\combined_out[2] ));
 sky130_fd_sc_hd__ebufn_4 \genblk2[3].lm_dt_out_buf[3]  (.A(\genblk2[3].selected_out[3] ),
    .TE_B(\genblk2[3].partition_sel_n ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\combined_out[3] ));
 sky130_fd_sc_hd__ebufn_4 \genblk2[3].lm_dt_out_buf[4]  (.A(\genblk2[3].selected_out[4] ),
    .TE_B(\genblk2[3].partition_sel_n ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\combined_out[4] ));
 sky130_fd_sc_hd__ebufn_4 \genblk2[3].lm_dt_out_buf[5]  (.A(\genblk2[3].selected_out[5] ),
    .TE_B(\genblk2[3].partition_sel_n ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\combined_out[5] ));
 sky130_fd_sc_hd__ebufn_4 \genblk2[3].lm_dt_out_buf[6]  (.A(\genblk2[3].selected_out[6] ),
    .TE_B(\genblk2[3].partition_sel_n ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\combined_out[6] ));
 sky130_fd_sc_hd__ebufn_4 \genblk2[3].lm_dt_out_buf[7]  (.A(\genblk2[3].selected_out[7] ),
    .TE_B(\genblk2[3].partition_sel_n ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Z(\combined_out[7] ));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(wr_en_next),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net113));
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(rst_n),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(uio_in[1]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(uio_in[2]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_1 input12 (.A(uio_in[3]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_1 input13 (.A(uio_in[4]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_1 input14 (.A(uio_in[5]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_1 input15 (.A(uio_in[6]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_1 input16 (.A(uio_in[7]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(ui_in[0]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(ui_in[1]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(ui_in[2]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(ui_in[3]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net5));
 sky130_fd_sc_hd__dlymetal6s2s_1 input6 (.A(ui_in[4]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net6));
 sky130_fd_sc_hd__dlymetal6s2s_1 input7 (.A(ui_in[5]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(ui_in[7]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_1 input9 (.A(uio_in[0]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_4 \lm_dt_final_buf[0]  (.A(\combined_out[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[0]));
 sky130_fd_sc_hd__clkbuf_4 \lm_dt_final_buf[1]  (.A(\combined_out[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[1]));
 sky130_fd_sc_hd__clkbuf_4 \lm_dt_final_buf[2]  (.A(\combined_out[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[2]));
 sky130_fd_sc_hd__clkbuf_4 \lm_dt_final_buf[3]  (.A(\combined_out[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[3]));
 sky130_fd_sc_hd__clkbuf_4 \lm_dt_final_buf[4]  (.A(\combined_out[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[4]));
 sky130_fd_sc_hd__clkbuf_4 \lm_dt_final_buf[5]  (.A(\combined_out[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[5]));
 sky130_fd_sc_hd__clkbuf_4 \lm_dt_final_buf[6]  (.A(\combined_out[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[6]));
 sky130_fd_sc_hd__clkbuf_4 \lm_dt_final_buf[7]  (.A(\combined_out[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[7]));
 sky130_fd_sc_hd__clkbuf_1 max_cap2 (.A(_0264_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net115));
 sky130_fd_sc_hd__clkbuf_2 max_cap25 (.A(net114),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net25));
 sky130_fd_sc_hd__buf_1 max_cap27 (.A(_0268_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net27));
 sky130_fd_sc_hd__conb_1 tt_um_MichaelBell_latch_mem_100 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net100));
 sky130_fd_sc_hd__conb_1 tt_um_MichaelBell_latch_mem_101 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net101));
 sky130_fd_sc_hd__conb_1 tt_um_MichaelBell_latch_mem_102 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net102));
 sky130_fd_sc_hd__conb_1 tt_um_MichaelBell_latch_mem_103 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net103));
 sky130_fd_sc_hd__conb_1 tt_um_MichaelBell_latch_mem_104 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net104));
 sky130_fd_sc_hd__conb_1 tt_um_MichaelBell_latch_mem_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net105));
 sky130_fd_sc_hd__conb_1 tt_um_MichaelBell_latch_mem_106 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net106));
 sky130_fd_sc_hd__conb_1 tt_um_MichaelBell_latch_mem_107 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net107));
 sky130_fd_sc_hd__conb_1 tt_um_MichaelBell_latch_mem_108 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net108));
 sky130_fd_sc_hd__conb_1 tt_um_MichaelBell_latch_mem_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net109));
 sky130_fd_sc_hd__conb_1 tt_um_MichaelBell_latch_mem_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net110));
 sky130_fd_sc_hd__conb_1 tt_um_MichaelBell_latch_mem_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net111));
 sky130_fd_sc_hd__conb_1 tt_um_MichaelBell_latch_mem_96 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net96));
 sky130_fd_sc_hd__conb_1 tt_um_MichaelBell_latch_mem_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net97));
 sky130_fd_sc_hd__conb_1 tt_um_MichaelBell_latch_mem_98 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net98));
 sky130_fd_sc_hd__conb_1 tt_um_MichaelBell_latch_mem_99 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net99));
 sky130_fd_sc_hd__buf_1 wire1 (.A(_0280_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net114));
 sky130_fd_sc_hd__clkbuf_2 wire26 (.A(_0277_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net26));
 sky130_fd_sc_hd__buf_2 wire28 (.A(_0264_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net28));
 assign uio_oe[0] = net96;
 assign uio_oe[1] = net97;
 assign uio_oe[2] = net98;
 assign uio_oe[3] = net99;
 assign uio_oe[4] = net100;
 assign uio_oe[5] = net101;
 assign uio_oe[6] = net102;
 assign uio_oe[7] = net103;
 assign uio_out[0] = net104;
 assign uio_out[1] = net105;
 assign uio_out[2] = net106;
 assign uio_out[3] = net107;
 assign uio_out[4] = net108;
 assign uio_out[5] = net109;
 assign uio_out[6] = net110;
 assign uio_out[7] = net111;
endmodule
