module tt_um_hpretl_tt06_tdc (VGND,
    VPWR,
    clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input VGND;
 input VPWR;
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire clknet_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire net1;
 wire net2;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire \tdc0.o_result[0] ;
 wire \tdc0.o_result[100] ;
 wire \tdc0.o_result[101] ;
 wire \tdc0.o_result[102] ;
 wire \tdc0.o_result[103] ;
 wire \tdc0.o_result[104] ;
 wire \tdc0.o_result[105] ;
 wire \tdc0.o_result[106] ;
 wire \tdc0.o_result[107] ;
 wire \tdc0.o_result[108] ;
 wire \tdc0.o_result[109] ;
 wire \tdc0.o_result[10] ;
 wire \tdc0.o_result[110] ;
 wire \tdc0.o_result[111] ;
 wire \tdc0.o_result[112] ;
 wire \tdc0.o_result[113] ;
 wire \tdc0.o_result[114] ;
 wire \tdc0.o_result[115] ;
 wire \tdc0.o_result[116] ;
 wire \tdc0.o_result[117] ;
 wire \tdc0.o_result[118] ;
 wire \tdc0.o_result[119] ;
 wire \tdc0.o_result[11] ;
 wire \tdc0.o_result[120] ;
 wire \tdc0.o_result[121] ;
 wire \tdc0.o_result[122] ;
 wire \tdc0.o_result[123] ;
 wire \tdc0.o_result[124] ;
 wire \tdc0.o_result[125] ;
 wire \tdc0.o_result[126] ;
 wire \tdc0.o_result[127] ;
 wire \tdc0.o_result[128] ;
 wire \tdc0.o_result[129] ;
 wire \tdc0.o_result[12] ;
 wire \tdc0.o_result[130] ;
 wire \tdc0.o_result[131] ;
 wire \tdc0.o_result[132] ;
 wire \tdc0.o_result[133] ;
 wire \tdc0.o_result[134] ;
 wire \tdc0.o_result[135] ;
 wire \tdc0.o_result[136] ;
 wire \tdc0.o_result[137] ;
 wire \tdc0.o_result[138] ;
 wire \tdc0.o_result[139] ;
 wire \tdc0.o_result[13] ;
 wire \tdc0.o_result[140] ;
 wire \tdc0.o_result[141] ;
 wire \tdc0.o_result[142] ;
 wire \tdc0.o_result[143] ;
 wire \tdc0.o_result[144] ;
 wire \tdc0.o_result[145] ;
 wire \tdc0.o_result[146] ;
 wire \tdc0.o_result[147] ;
 wire \tdc0.o_result[148] ;
 wire \tdc0.o_result[149] ;
 wire \tdc0.o_result[14] ;
 wire \tdc0.o_result[150] ;
 wire \tdc0.o_result[151] ;
 wire \tdc0.o_result[152] ;
 wire \tdc0.o_result[153] ;
 wire \tdc0.o_result[154] ;
 wire \tdc0.o_result[155] ;
 wire \tdc0.o_result[156] ;
 wire \tdc0.o_result[157] ;
 wire \tdc0.o_result[158] ;
 wire \tdc0.o_result[159] ;
 wire \tdc0.o_result[15] ;
 wire \tdc0.o_result[160] ;
 wire \tdc0.o_result[161] ;
 wire \tdc0.o_result[162] ;
 wire \tdc0.o_result[163] ;
 wire \tdc0.o_result[164] ;
 wire \tdc0.o_result[165] ;
 wire \tdc0.o_result[166] ;
 wire \tdc0.o_result[167] ;
 wire \tdc0.o_result[168] ;
 wire \tdc0.o_result[169] ;
 wire \tdc0.o_result[16] ;
 wire \tdc0.o_result[170] ;
 wire \tdc0.o_result[171] ;
 wire \tdc0.o_result[172] ;
 wire \tdc0.o_result[173] ;
 wire \tdc0.o_result[174] ;
 wire \tdc0.o_result[175] ;
 wire \tdc0.o_result[176] ;
 wire \tdc0.o_result[177] ;
 wire \tdc0.o_result[178] ;
 wire \tdc0.o_result[179] ;
 wire \tdc0.o_result[17] ;
 wire \tdc0.o_result[180] ;
 wire \tdc0.o_result[181] ;
 wire \tdc0.o_result[182] ;
 wire \tdc0.o_result[183] ;
 wire \tdc0.o_result[184] ;
 wire \tdc0.o_result[185] ;
 wire \tdc0.o_result[186] ;
 wire \tdc0.o_result[187] ;
 wire \tdc0.o_result[188] ;
 wire \tdc0.o_result[189] ;
 wire \tdc0.o_result[18] ;
 wire \tdc0.o_result[190] ;
 wire \tdc0.o_result[191] ;
 wire \tdc0.o_result[19] ;
 wire \tdc0.o_result[1] ;
 wire \tdc0.o_result[20] ;
 wire \tdc0.o_result[21] ;
 wire \tdc0.o_result[22] ;
 wire \tdc0.o_result[23] ;
 wire \tdc0.o_result[24] ;
 wire \tdc0.o_result[25] ;
 wire \tdc0.o_result[26] ;
 wire \tdc0.o_result[27] ;
 wire \tdc0.o_result[28] ;
 wire \tdc0.o_result[29] ;
 wire \tdc0.o_result[2] ;
 wire \tdc0.o_result[30] ;
 wire \tdc0.o_result[31] ;
 wire \tdc0.o_result[32] ;
 wire \tdc0.o_result[33] ;
 wire \tdc0.o_result[34] ;
 wire \tdc0.o_result[35] ;
 wire \tdc0.o_result[36] ;
 wire \tdc0.o_result[37] ;
 wire \tdc0.o_result[38] ;
 wire \tdc0.o_result[39] ;
 wire \tdc0.o_result[3] ;
 wire \tdc0.o_result[40] ;
 wire \tdc0.o_result[41] ;
 wire \tdc0.o_result[42] ;
 wire \tdc0.o_result[43] ;
 wire \tdc0.o_result[44] ;
 wire \tdc0.o_result[45] ;
 wire \tdc0.o_result[46] ;
 wire \tdc0.o_result[47] ;
 wire \tdc0.o_result[48] ;
 wire \tdc0.o_result[49] ;
 wire \tdc0.o_result[4] ;
 wire \tdc0.o_result[50] ;
 wire \tdc0.o_result[51] ;
 wire \tdc0.o_result[52] ;
 wire \tdc0.o_result[53] ;
 wire \tdc0.o_result[54] ;
 wire \tdc0.o_result[55] ;
 wire \tdc0.o_result[56] ;
 wire \tdc0.o_result[57] ;
 wire \tdc0.o_result[58] ;
 wire \tdc0.o_result[59] ;
 wire \tdc0.o_result[5] ;
 wire \tdc0.o_result[60] ;
 wire \tdc0.o_result[61] ;
 wire \tdc0.o_result[62] ;
 wire \tdc0.o_result[63] ;
 wire \tdc0.o_result[64] ;
 wire \tdc0.o_result[65] ;
 wire \tdc0.o_result[66] ;
 wire \tdc0.o_result[67] ;
 wire \tdc0.o_result[68] ;
 wire \tdc0.o_result[69] ;
 wire \tdc0.o_result[6] ;
 wire \tdc0.o_result[70] ;
 wire \tdc0.o_result[71] ;
 wire \tdc0.o_result[72] ;
 wire \tdc0.o_result[73] ;
 wire \tdc0.o_result[74] ;
 wire \tdc0.o_result[75] ;
 wire \tdc0.o_result[76] ;
 wire \tdc0.o_result[77] ;
 wire \tdc0.o_result[78] ;
 wire \tdc0.o_result[79] ;
 wire \tdc0.o_result[7] ;
 wire \tdc0.o_result[80] ;
 wire \tdc0.o_result[81] ;
 wire \tdc0.o_result[82] ;
 wire \tdc0.o_result[83] ;
 wire \tdc0.o_result[84] ;
 wire \tdc0.o_result[85] ;
 wire \tdc0.o_result[86] ;
 wire \tdc0.o_result[87] ;
 wire \tdc0.o_result[88] ;
 wire \tdc0.o_result[89] ;
 wire \tdc0.o_result[8] ;
 wire \tdc0.o_result[90] ;
 wire \tdc0.o_result[91] ;
 wire \tdc0.o_result[92] ;
 wire \tdc0.o_result[93] ;
 wire \tdc0.o_result[94] ;
 wire \tdc0.o_result[95] ;
 wire \tdc0.o_result[96] ;
 wire \tdc0.o_result[97] ;
 wire \tdc0.o_result[98] ;
 wire \tdc0.o_result[99] ;
 wire \tdc0.o_result[9] ;
 wire \tdc0.w_dly_sig[0] ;
 wire \tdc0.w_dly_sig[100] ;
 wire \tdc0.w_dly_sig[101] ;
 wire \tdc0.w_dly_sig[102] ;
 wire \tdc0.w_dly_sig[103] ;
 wire \tdc0.w_dly_sig[104] ;
 wire \tdc0.w_dly_sig[105] ;
 wire \tdc0.w_dly_sig[106] ;
 wire \tdc0.w_dly_sig[107] ;
 wire \tdc0.w_dly_sig[108] ;
 wire \tdc0.w_dly_sig[109] ;
 wire \tdc0.w_dly_sig[10] ;
 wire \tdc0.w_dly_sig[110] ;
 wire \tdc0.w_dly_sig[111] ;
 wire \tdc0.w_dly_sig[112] ;
 wire \tdc0.w_dly_sig[113] ;
 wire \tdc0.w_dly_sig[114] ;
 wire \tdc0.w_dly_sig[115] ;
 wire \tdc0.w_dly_sig[116] ;
 wire \tdc0.w_dly_sig[117] ;
 wire \tdc0.w_dly_sig[118] ;
 wire \tdc0.w_dly_sig[119] ;
 wire \tdc0.w_dly_sig[11] ;
 wire \tdc0.w_dly_sig[120] ;
 wire \tdc0.w_dly_sig[121] ;
 wire \tdc0.w_dly_sig[122] ;
 wire \tdc0.w_dly_sig[123] ;
 wire \tdc0.w_dly_sig[124] ;
 wire \tdc0.w_dly_sig[125] ;
 wire \tdc0.w_dly_sig[126] ;
 wire \tdc0.w_dly_sig[127] ;
 wire \tdc0.w_dly_sig[128] ;
 wire \tdc0.w_dly_sig[129] ;
 wire \tdc0.w_dly_sig[12] ;
 wire \tdc0.w_dly_sig[130] ;
 wire \tdc0.w_dly_sig[131] ;
 wire \tdc0.w_dly_sig[132] ;
 wire \tdc0.w_dly_sig[133] ;
 wire \tdc0.w_dly_sig[134] ;
 wire \tdc0.w_dly_sig[135] ;
 wire \tdc0.w_dly_sig[136] ;
 wire \tdc0.w_dly_sig[137] ;
 wire \tdc0.w_dly_sig[138] ;
 wire \tdc0.w_dly_sig[139] ;
 wire \tdc0.w_dly_sig[13] ;
 wire \tdc0.w_dly_sig[140] ;
 wire \tdc0.w_dly_sig[141] ;
 wire \tdc0.w_dly_sig[142] ;
 wire \tdc0.w_dly_sig[143] ;
 wire \tdc0.w_dly_sig[144] ;
 wire \tdc0.w_dly_sig[145] ;
 wire \tdc0.w_dly_sig[146] ;
 wire \tdc0.w_dly_sig[147] ;
 wire \tdc0.w_dly_sig[148] ;
 wire \tdc0.w_dly_sig[149] ;
 wire \tdc0.w_dly_sig[14] ;
 wire \tdc0.w_dly_sig[150] ;
 wire \tdc0.w_dly_sig[151] ;
 wire \tdc0.w_dly_sig[152] ;
 wire \tdc0.w_dly_sig[153] ;
 wire \tdc0.w_dly_sig[154] ;
 wire \tdc0.w_dly_sig[155] ;
 wire \tdc0.w_dly_sig[156] ;
 wire \tdc0.w_dly_sig[157] ;
 wire \tdc0.w_dly_sig[158] ;
 wire \tdc0.w_dly_sig[159] ;
 wire \tdc0.w_dly_sig[15] ;
 wire \tdc0.w_dly_sig[160] ;
 wire \tdc0.w_dly_sig[161] ;
 wire \tdc0.w_dly_sig[162] ;
 wire \tdc0.w_dly_sig[163] ;
 wire \tdc0.w_dly_sig[164] ;
 wire \tdc0.w_dly_sig[165] ;
 wire \tdc0.w_dly_sig[166] ;
 wire \tdc0.w_dly_sig[167] ;
 wire \tdc0.w_dly_sig[168] ;
 wire \tdc0.w_dly_sig[169] ;
 wire \tdc0.w_dly_sig[16] ;
 wire \tdc0.w_dly_sig[170] ;
 wire \tdc0.w_dly_sig[171] ;
 wire \tdc0.w_dly_sig[172] ;
 wire \tdc0.w_dly_sig[173] ;
 wire \tdc0.w_dly_sig[174] ;
 wire \tdc0.w_dly_sig[175] ;
 wire \tdc0.w_dly_sig[176] ;
 wire \tdc0.w_dly_sig[177] ;
 wire \tdc0.w_dly_sig[178] ;
 wire \tdc0.w_dly_sig[179] ;
 wire \tdc0.w_dly_sig[17] ;
 wire \tdc0.w_dly_sig[180] ;
 wire \tdc0.w_dly_sig[181] ;
 wire \tdc0.w_dly_sig[182] ;
 wire \tdc0.w_dly_sig[183] ;
 wire \tdc0.w_dly_sig[184] ;
 wire \tdc0.w_dly_sig[185] ;
 wire \tdc0.w_dly_sig[186] ;
 wire \tdc0.w_dly_sig[187] ;
 wire \tdc0.w_dly_sig[188] ;
 wire \tdc0.w_dly_sig[189] ;
 wire \tdc0.w_dly_sig[18] ;
 wire \tdc0.w_dly_sig[190] ;
 wire \tdc0.w_dly_sig[191] ;
 wire \tdc0.w_dly_sig[192] ;
 wire \tdc0.w_dly_sig[193] ;
 wire \tdc0.w_dly_sig[19] ;
 wire \tdc0.w_dly_sig[1] ;
 wire \tdc0.w_dly_sig[20] ;
 wire \tdc0.w_dly_sig[21] ;
 wire \tdc0.w_dly_sig[22] ;
 wire \tdc0.w_dly_sig[23] ;
 wire \tdc0.w_dly_sig[24] ;
 wire \tdc0.w_dly_sig[25] ;
 wire \tdc0.w_dly_sig[26] ;
 wire \tdc0.w_dly_sig[27] ;
 wire \tdc0.w_dly_sig[28] ;
 wire \tdc0.w_dly_sig[29] ;
 wire \tdc0.w_dly_sig[2] ;
 wire \tdc0.w_dly_sig[30] ;
 wire \tdc0.w_dly_sig[31] ;
 wire \tdc0.w_dly_sig[32] ;
 wire \tdc0.w_dly_sig[33] ;
 wire \tdc0.w_dly_sig[34] ;
 wire \tdc0.w_dly_sig[35] ;
 wire \tdc0.w_dly_sig[36] ;
 wire \tdc0.w_dly_sig[37] ;
 wire \tdc0.w_dly_sig[38] ;
 wire \tdc0.w_dly_sig[39] ;
 wire \tdc0.w_dly_sig[3] ;
 wire \tdc0.w_dly_sig[40] ;
 wire \tdc0.w_dly_sig[41] ;
 wire \tdc0.w_dly_sig[42] ;
 wire \tdc0.w_dly_sig[43] ;
 wire \tdc0.w_dly_sig[44] ;
 wire \tdc0.w_dly_sig[45] ;
 wire \tdc0.w_dly_sig[46] ;
 wire \tdc0.w_dly_sig[47] ;
 wire \tdc0.w_dly_sig[48] ;
 wire \tdc0.w_dly_sig[49] ;
 wire \tdc0.w_dly_sig[4] ;
 wire \tdc0.w_dly_sig[50] ;
 wire \tdc0.w_dly_sig[51] ;
 wire \tdc0.w_dly_sig[52] ;
 wire \tdc0.w_dly_sig[53] ;
 wire \tdc0.w_dly_sig[54] ;
 wire \tdc0.w_dly_sig[55] ;
 wire \tdc0.w_dly_sig[56] ;
 wire \tdc0.w_dly_sig[57] ;
 wire \tdc0.w_dly_sig[58] ;
 wire \tdc0.w_dly_sig[59] ;
 wire \tdc0.w_dly_sig[5] ;
 wire \tdc0.w_dly_sig[60] ;
 wire \tdc0.w_dly_sig[61] ;
 wire \tdc0.w_dly_sig[62] ;
 wire \tdc0.w_dly_sig[63] ;
 wire \tdc0.w_dly_sig[64] ;
 wire \tdc0.w_dly_sig[65] ;
 wire \tdc0.w_dly_sig[66] ;
 wire \tdc0.w_dly_sig[67] ;
 wire \tdc0.w_dly_sig[68] ;
 wire \tdc0.w_dly_sig[69] ;
 wire \tdc0.w_dly_sig[6] ;
 wire \tdc0.w_dly_sig[70] ;
 wire \tdc0.w_dly_sig[71] ;
 wire \tdc0.w_dly_sig[72] ;
 wire \tdc0.w_dly_sig[73] ;
 wire \tdc0.w_dly_sig[74] ;
 wire \tdc0.w_dly_sig[75] ;
 wire \tdc0.w_dly_sig[76] ;
 wire \tdc0.w_dly_sig[77] ;
 wire \tdc0.w_dly_sig[78] ;
 wire \tdc0.w_dly_sig[79] ;
 wire \tdc0.w_dly_sig[7] ;
 wire \tdc0.w_dly_sig[80] ;
 wire \tdc0.w_dly_sig[81] ;
 wire \tdc0.w_dly_sig[82] ;
 wire \tdc0.w_dly_sig[83] ;
 wire \tdc0.w_dly_sig[84] ;
 wire \tdc0.w_dly_sig[85] ;
 wire \tdc0.w_dly_sig[86] ;
 wire \tdc0.w_dly_sig[87] ;
 wire \tdc0.w_dly_sig[88] ;
 wire \tdc0.w_dly_sig[89] ;
 wire \tdc0.w_dly_sig[8] ;
 wire \tdc0.w_dly_sig[90] ;
 wire \tdc0.w_dly_sig[91] ;
 wire \tdc0.w_dly_sig[92] ;
 wire \tdc0.w_dly_sig[93] ;
 wire \tdc0.w_dly_sig[94] ;
 wire \tdc0.w_dly_sig[95] ;
 wire \tdc0.w_dly_sig[96] ;
 wire \tdc0.w_dly_sig[97] ;
 wire \tdc0.w_dly_sig[98] ;
 wire \tdc0.w_dly_sig[99] ;
 wire \tdc0.w_dly_sig[9] ;
 wire \tdc0.w_dly_sig_n[0] ;
 wire \tdc0.w_dly_sig_n[100] ;
 wire \tdc0.w_dly_sig_n[101] ;
 wire \tdc0.w_dly_sig_n[102] ;
 wire \tdc0.w_dly_sig_n[103] ;
 wire \tdc0.w_dly_sig_n[104] ;
 wire \tdc0.w_dly_sig_n[105] ;
 wire \tdc0.w_dly_sig_n[106] ;
 wire \tdc0.w_dly_sig_n[107] ;
 wire \tdc0.w_dly_sig_n[108] ;
 wire \tdc0.w_dly_sig_n[109] ;
 wire \tdc0.w_dly_sig_n[10] ;
 wire \tdc0.w_dly_sig_n[110] ;
 wire \tdc0.w_dly_sig_n[111] ;
 wire \tdc0.w_dly_sig_n[112] ;
 wire \tdc0.w_dly_sig_n[113] ;
 wire \tdc0.w_dly_sig_n[114] ;
 wire \tdc0.w_dly_sig_n[115] ;
 wire \tdc0.w_dly_sig_n[116] ;
 wire \tdc0.w_dly_sig_n[117] ;
 wire \tdc0.w_dly_sig_n[118] ;
 wire \tdc0.w_dly_sig_n[119] ;
 wire \tdc0.w_dly_sig_n[11] ;
 wire \tdc0.w_dly_sig_n[120] ;
 wire \tdc0.w_dly_sig_n[121] ;
 wire \tdc0.w_dly_sig_n[122] ;
 wire \tdc0.w_dly_sig_n[123] ;
 wire \tdc0.w_dly_sig_n[124] ;
 wire \tdc0.w_dly_sig_n[125] ;
 wire \tdc0.w_dly_sig_n[126] ;
 wire \tdc0.w_dly_sig_n[127] ;
 wire \tdc0.w_dly_sig_n[128] ;
 wire \tdc0.w_dly_sig_n[129] ;
 wire \tdc0.w_dly_sig_n[12] ;
 wire \tdc0.w_dly_sig_n[130] ;
 wire \tdc0.w_dly_sig_n[131] ;
 wire \tdc0.w_dly_sig_n[132] ;
 wire \tdc0.w_dly_sig_n[133] ;
 wire \tdc0.w_dly_sig_n[134] ;
 wire \tdc0.w_dly_sig_n[135] ;
 wire \tdc0.w_dly_sig_n[136] ;
 wire \tdc0.w_dly_sig_n[137] ;
 wire \tdc0.w_dly_sig_n[138] ;
 wire \tdc0.w_dly_sig_n[139] ;
 wire \tdc0.w_dly_sig_n[13] ;
 wire \tdc0.w_dly_sig_n[140] ;
 wire \tdc0.w_dly_sig_n[141] ;
 wire \tdc0.w_dly_sig_n[142] ;
 wire \tdc0.w_dly_sig_n[143] ;
 wire \tdc0.w_dly_sig_n[144] ;
 wire \tdc0.w_dly_sig_n[145] ;
 wire \tdc0.w_dly_sig_n[146] ;
 wire \tdc0.w_dly_sig_n[147] ;
 wire \tdc0.w_dly_sig_n[148] ;
 wire \tdc0.w_dly_sig_n[149] ;
 wire \tdc0.w_dly_sig_n[14] ;
 wire \tdc0.w_dly_sig_n[150] ;
 wire \tdc0.w_dly_sig_n[151] ;
 wire \tdc0.w_dly_sig_n[152] ;
 wire \tdc0.w_dly_sig_n[153] ;
 wire \tdc0.w_dly_sig_n[154] ;
 wire \tdc0.w_dly_sig_n[155] ;
 wire \tdc0.w_dly_sig_n[156] ;
 wire \tdc0.w_dly_sig_n[157] ;
 wire \tdc0.w_dly_sig_n[158] ;
 wire \tdc0.w_dly_sig_n[159] ;
 wire \tdc0.w_dly_sig_n[15] ;
 wire \tdc0.w_dly_sig_n[160] ;
 wire \tdc0.w_dly_sig_n[161] ;
 wire \tdc0.w_dly_sig_n[162] ;
 wire \tdc0.w_dly_sig_n[163] ;
 wire \tdc0.w_dly_sig_n[164] ;
 wire \tdc0.w_dly_sig_n[165] ;
 wire \tdc0.w_dly_sig_n[166] ;
 wire \tdc0.w_dly_sig_n[167] ;
 wire \tdc0.w_dly_sig_n[168] ;
 wire \tdc0.w_dly_sig_n[169] ;
 wire \tdc0.w_dly_sig_n[16] ;
 wire \tdc0.w_dly_sig_n[170] ;
 wire \tdc0.w_dly_sig_n[171] ;
 wire \tdc0.w_dly_sig_n[172] ;
 wire \tdc0.w_dly_sig_n[173] ;
 wire \tdc0.w_dly_sig_n[174] ;
 wire \tdc0.w_dly_sig_n[175] ;
 wire \tdc0.w_dly_sig_n[176] ;
 wire \tdc0.w_dly_sig_n[177] ;
 wire \tdc0.w_dly_sig_n[178] ;
 wire \tdc0.w_dly_sig_n[179] ;
 wire \tdc0.w_dly_sig_n[17] ;
 wire \tdc0.w_dly_sig_n[180] ;
 wire \tdc0.w_dly_sig_n[181] ;
 wire \tdc0.w_dly_sig_n[182] ;
 wire \tdc0.w_dly_sig_n[183] ;
 wire \tdc0.w_dly_sig_n[184] ;
 wire \tdc0.w_dly_sig_n[185] ;
 wire \tdc0.w_dly_sig_n[186] ;
 wire \tdc0.w_dly_sig_n[187] ;
 wire \tdc0.w_dly_sig_n[188] ;
 wire \tdc0.w_dly_sig_n[189] ;
 wire \tdc0.w_dly_sig_n[18] ;
 wire \tdc0.w_dly_sig_n[190] ;
 wire \tdc0.w_dly_sig_n[191] ;
 wire \tdc0.w_dly_sig_n[192] ;
 wire \tdc0.w_dly_sig_n[19] ;
 wire \tdc0.w_dly_sig_n[1] ;
 wire \tdc0.w_dly_sig_n[20] ;
 wire \tdc0.w_dly_sig_n[21] ;
 wire \tdc0.w_dly_sig_n[22] ;
 wire \tdc0.w_dly_sig_n[23] ;
 wire \tdc0.w_dly_sig_n[24] ;
 wire \tdc0.w_dly_sig_n[25] ;
 wire \tdc0.w_dly_sig_n[26] ;
 wire \tdc0.w_dly_sig_n[27] ;
 wire \tdc0.w_dly_sig_n[28] ;
 wire \tdc0.w_dly_sig_n[29] ;
 wire \tdc0.w_dly_sig_n[2] ;
 wire \tdc0.w_dly_sig_n[30] ;
 wire \tdc0.w_dly_sig_n[31] ;
 wire \tdc0.w_dly_sig_n[32] ;
 wire \tdc0.w_dly_sig_n[33] ;
 wire \tdc0.w_dly_sig_n[34] ;
 wire \tdc0.w_dly_sig_n[35] ;
 wire \tdc0.w_dly_sig_n[36] ;
 wire \tdc0.w_dly_sig_n[37] ;
 wire \tdc0.w_dly_sig_n[38] ;
 wire \tdc0.w_dly_sig_n[39] ;
 wire \tdc0.w_dly_sig_n[3] ;
 wire \tdc0.w_dly_sig_n[40] ;
 wire \tdc0.w_dly_sig_n[41] ;
 wire \tdc0.w_dly_sig_n[42] ;
 wire \tdc0.w_dly_sig_n[43] ;
 wire \tdc0.w_dly_sig_n[44] ;
 wire \tdc0.w_dly_sig_n[45] ;
 wire \tdc0.w_dly_sig_n[46] ;
 wire \tdc0.w_dly_sig_n[47] ;
 wire \tdc0.w_dly_sig_n[48] ;
 wire \tdc0.w_dly_sig_n[49] ;
 wire \tdc0.w_dly_sig_n[4] ;
 wire \tdc0.w_dly_sig_n[50] ;
 wire \tdc0.w_dly_sig_n[51] ;
 wire \tdc0.w_dly_sig_n[52] ;
 wire \tdc0.w_dly_sig_n[53] ;
 wire \tdc0.w_dly_sig_n[54] ;
 wire \tdc0.w_dly_sig_n[55] ;
 wire \tdc0.w_dly_sig_n[56] ;
 wire \tdc0.w_dly_sig_n[57] ;
 wire \tdc0.w_dly_sig_n[58] ;
 wire \tdc0.w_dly_sig_n[59] ;
 wire \tdc0.w_dly_sig_n[5] ;
 wire \tdc0.w_dly_sig_n[60] ;
 wire \tdc0.w_dly_sig_n[61] ;
 wire \tdc0.w_dly_sig_n[62] ;
 wire \tdc0.w_dly_sig_n[63] ;
 wire \tdc0.w_dly_sig_n[64] ;
 wire \tdc0.w_dly_sig_n[65] ;
 wire \tdc0.w_dly_sig_n[66] ;
 wire \tdc0.w_dly_sig_n[67] ;
 wire \tdc0.w_dly_sig_n[68] ;
 wire \tdc0.w_dly_sig_n[69] ;
 wire \tdc0.w_dly_sig_n[6] ;
 wire \tdc0.w_dly_sig_n[70] ;
 wire \tdc0.w_dly_sig_n[71] ;
 wire \tdc0.w_dly_sig_n[72] ;
 wire \tdc0.w_dly_sig_n[73] ;
 wire \tdc0.w_dly_sig_n[74] ;
 wire \tdc0.w_dly_sig_n[75] ;
 wire \tdc0.w_dly_sig_n[76] ;
 wire \tdc0.w_dly_sig_n[77] ;
 wire \tdc0.w_dly_sig_n[78] ;
 wire \tdc0.w_dly_sig_n[79] ;
 wire \tdc0.w_dly_sig_n[7] ;
 wire \tdc0.w_dly_sig_n[80] ;
 wire \tdc0.w_dly_sig_n[81] ;
 wire \tdc0.w_dly_sig_n[82] ;
 wire \tdc0.w_dly_sig_n[83] ;
 wire \tdc0.w_dly_sig_n[84] ;
 wire \tdc0.w_dly_sig_n[85] ;
 wire \tdc0.w_dly_sig_n[86] ;
 wire \tdc0.w_dly_sig_n[87] ;
 wire \tdc0.w_dly_sig_n[88] ;
 wire \tdc0.w_dly_sig_n[89] ;
 wire \tdc0.w_dly_sig_n[8] ;
 wire \tdc0.w_dly_sig_n[90] ;
 wire \tdc0.w_dly_sig_n[91] ;
 wire \tdc0.w_dly_sig_n[92] ;
 wire \tdc0.w_dly_sig_n[93] ;
 wire \tdc0.w_dly_sig_n[94] ;
 wire \tdc0.w_dly_sig_n[95] ;
 wire \tdc0.w_dly_sig_n[96] ;
 wire \tdc0.w_dly_sig_n[97] ;
 wire \tdc0.w_dly_sig_n[98] ;
 wire \tdc0.w_dly_sig_n[99] ;
 wire \tdc0.w_dly_sig_n[9] ;

 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(\tdc0.o_result[101] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_113 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_125 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_141 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_153 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_165 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_169 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_181 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_193 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_197 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_209 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_221 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_225 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_237 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_249 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_253 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_265 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_277 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_281 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_293 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_305 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_309 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_321 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_0_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_41 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_69 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_85 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_97 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_106 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_10_118 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_124 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_10_136 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_10_148 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_10_168 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_10_202 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_10_215 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_10_229 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_10_240 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_10_249 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_259 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_271 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_294 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_306 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_309 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_321 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_53 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_10_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_10_73 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_94 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_11_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_11_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_135 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_11_144 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_155 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_11_186 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_11_199 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_11_239 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_27 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_11_274 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_11_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_289 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_306 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_318 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_11_330 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_39 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_11_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_57 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_101 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_107 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_125 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_12_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_148 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_160 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_172 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_188 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_12_211 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_215 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_12_221 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_229 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_12_240 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_12_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_259 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_12_275 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_283 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_290 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_12_301 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_12_325 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_12_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_50 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_67 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_85 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_12_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_13_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_13_131 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_155 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_13_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_13_191 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_13_199 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_13_213 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_13_221 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_13_241 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_263 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_13_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_13_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_13_332 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_13_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_60 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_13_70 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_13_78 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_13_87 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_13_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_14_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_119 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_14_158 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_172 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_14_193 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_14_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_14_209 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_14_218 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_14_224 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_237 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_14_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_253 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_14_265 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_273 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_285 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_300 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_14_324 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_14_332 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_14_48 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_14_75 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_118 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_15_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_15_155 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_15_163 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_190 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_240 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_266 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_297 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_15_313 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_15_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_15_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_92 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_16_123 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_127 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_16_131 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_16_164 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_170 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_16_174 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_180 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_16_184 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_188 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_16_192 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_16_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_16_22 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_16_222 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_237 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_16_249 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_16_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_16_273 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_16_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_29 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_16_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_16_303 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_16_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_50 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_67 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_16_79 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_16_96 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_17_108 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_17_147 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_163 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_174 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_17_199 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_207 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_17_22 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_17_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_229 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_17_246 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_258 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_17_277 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_295 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_17_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_31 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_17_312 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_17_330 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_17_38 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_46 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_17_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_64 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_76 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_96 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_18_116 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_124 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_18_134 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_18_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_18_160 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_18_171 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_177 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_18_189 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_18_20 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_234 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_246 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_268 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_18_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_306 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_18_315 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_18_38 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_104 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_19_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_143 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_19_155 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_19_165 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_19_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_19_203 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_207 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_19_216 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_19_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_19_239 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_19_247 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_19_258 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_19_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_285 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_19_289 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_19_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_41 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_19_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_19_73 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_19_90 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_19_98 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_1_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_113 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_125 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_137 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_149 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_1_161 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_169 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_181 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_193 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_205 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_1_217 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_225 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_237 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_249 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_261 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_1_273 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_281 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_293 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_305 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_317 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_1_329 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_39 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_81 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_93 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_102 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_114 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_20_121 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_20_130 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_134 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_20_148 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_20_168 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_181 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_20_193 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_20_221 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_233 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_245 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_269 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_281 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_29 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_20_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_321 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_20_59 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_63 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_20_80 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_20_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_91 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_95 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_21_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_116 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_21_140 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_146 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_17 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_21_196 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_21_204 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_21_216 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_21_236 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_21_254 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_272 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_21_278 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_297 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_21_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_318 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_21_34 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_40 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_21_73 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_22_101 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_123 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_22_135 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_22_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_149 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_22_160 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_164 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_22_180 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_202 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_22_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_22_218 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_235 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_22_256 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_22_264 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_22_285 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_22_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_22_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_22_305 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_22_313 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_317 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_22_330 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_22_37 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_22_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_23_107 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_23_121 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_132 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_149 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_23_163 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_23_17 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_23_179 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_185 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_23_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_203 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_215 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_22 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_23_220 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_23_236 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_23_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_261 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_267 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_23_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_285 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_23_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_23_302 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_23_310 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_23_319 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_46 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_23_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_23_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_23_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_23_99 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_24_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_24_119 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_130 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_24_136 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_141 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_24_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_157 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_173 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_24_179 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_187 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_24_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_24_202 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_219 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_228 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_24_241 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_24_247 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_24_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_24_258 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_24_288 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_24_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_38 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_24_42 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_24_63 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_24_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_24_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_25_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_25_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_135 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_25_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_25_164 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_25_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_25_177 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_25_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_209 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_222 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_225 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_25_237 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_25_24 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_25_270 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_278 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_25_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_30 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_25_300 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_308 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_25_34 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_46 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_50 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_25_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_61 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_25_90 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_26_117 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_26_127 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_26_151 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_26_168 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_172 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_26_179 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_187 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_26_203 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_26_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_26_233 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_26_259 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_26_286 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_26_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_26_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_26_45 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_26_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_79 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_92 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_27_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_27_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_117 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_27_143 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_27_158 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_27_165 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_27_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_27_201 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_27_209 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_27_217 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_23 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_27_241 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_27_255 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_263 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_27_297 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_27_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_27_311 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_27_328 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_27_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_27_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_27_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_27_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_27_88 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_27_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_100 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_28_117 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_28_124 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_28_136 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_28_146 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_150 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_28_156 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_164 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_28_176 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_28_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_28_211 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_28_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_28_231 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_240 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_28_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_28_256 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_28_263 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_28_271 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_28_284 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_28_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_28_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_28_302 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_28_315 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_28_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_28_79 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_28_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_29_140 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_29_147 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_155 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_29_165 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_29_202 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_206 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_29_236 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_28 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_287 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_29_299 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_29_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_305 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_29_324 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_29_332 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_29_52 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_29_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_29_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_109 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_121 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_2_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_141 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_153 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_165 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_177 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_2_189 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_197 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_209 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_221 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_233 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_2_245 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_253 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_265 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_277 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_289 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_2_301 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_309 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_321 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_97 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_30_100 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_128 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_30_152 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_30_171 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_179 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_30_189 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_30_213 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_30_22 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_30_274 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_30_282 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_30_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_301 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_32 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_30_331 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_30_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_31_103 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_31_119 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_31_131 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_135 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_151 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_31_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_31_206 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_214 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_222 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_240 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_31_267 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_271 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_299 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_31_46 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_31_57 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_31_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_31_91 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_112 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_32_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_32_193 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_32_213 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_219 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_32_22 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_32_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_32_260 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_32_279 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_32_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_32_291 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_32_299 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_32_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_32_318 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_32_330 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_32_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_32_64 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_32_69 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_32_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_32_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_89 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_33_108 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_33_122 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_33_134 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_33_152 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_158 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_33_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_177 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_33_193 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_33_20 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_33_215 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_33_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_263 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_33_281 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_33_293 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_297 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_33_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_33_314 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_33_32 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_33_332 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_33_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_33_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_61 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_33_90 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_34_102 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_130 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_34_158 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_34_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_207 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_34_242 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_34_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_34_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_258 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_34_271 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_34_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_34_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_298 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_34_315 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_34_63 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_67 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_34_80 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_34_94 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_35_103 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_35_122 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_35_134 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_35_165 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_35_169 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_35_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_35_221 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_233 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_35_25 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_35_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_35_272 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_298 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_35_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_305 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_35_322 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_33 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_37 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_35_50 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_35_57 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_35_80 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_84 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_36_102 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_108 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_36_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_36_200 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_36_231 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_36_249 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_36_263 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_36_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_287 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_36_291 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_36_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_36_306 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_36_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_36_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_36_63 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_71 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_104 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_37_122 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_37_134 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_146 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_37_150 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_37_162 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_37_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_191 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_37_214 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_22 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_241 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_274 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_37_293 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_297 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_313 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_37_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_37_90 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_99 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_10 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_38_102 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_106 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_38_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_38_14 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_38_159 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_18 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_38_185 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_38_200 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_38_207 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_211 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_38_215 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_38_22 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_38_237 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_38_249 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_38_277 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_301 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_38_314 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_38_32 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_38_38 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_42 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_38_46 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_50 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_38_6 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_38_62 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_66 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_38_70 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_74 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_38_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_38_88 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_38_94 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_98 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_113 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_125 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_137 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_149 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_153 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_3_165 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_172 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_176 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_181 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_3_193 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_201 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_208 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_3_220 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_225 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_237 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_249 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_261 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_3_273 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_281 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_293 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_305 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_317 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_3_329 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_93 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_109 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_121 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_4_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_179 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_228 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_240 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_253 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_265 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_277 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_289 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_4_301 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_309 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_321 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_97 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_5_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_130 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_156 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_5_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_177 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_5_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_209 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_5_228 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_237 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_249 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_261 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_5_273 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_281 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_293 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_305 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_317 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_5_329 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_81 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_93 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_107 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_6_112 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_6_131 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_6_157 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_179 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_6_191 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_226 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_6_244 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_253 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_265 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_277 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_289 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_6_301 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_309 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_321 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_65 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_6_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_6_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_94 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_6_99 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_7_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_7_134 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_7_142 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_157 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_172 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_7_189 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_7_209 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_217 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_7_256 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_27 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_7_275 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_281 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_293 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_305 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_317 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_7_329 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_39 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_7_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_57 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_69 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_7_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_87 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_154 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_166 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_197 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_8_209 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_8_231 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_8_240 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_8_249 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_8_271 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_275 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_279 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_291 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_8_303 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_309 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_321 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_41 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_53 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_65 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_90 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_98 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_9_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_118 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_185 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_9_213 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_9_221 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_9_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_9_249 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_9_257 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_263 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_27 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_297 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_309 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_321 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_39 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_9_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_9_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_73 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_86 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_49 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_50 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_52 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_56 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_58 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_40 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_59 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_60 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_61 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_62 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_63 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_64 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_66 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_67 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_68 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_70 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_71 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_72 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_73 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_74 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_75 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_76 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_42 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_43 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_44 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_45 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_46 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_47 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_48 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_78 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_79 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_80 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_81 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_82 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_83 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_84 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_85 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_86 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_87 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_88 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_138 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_139 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_140 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_141 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_142 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_143 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_144 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_145 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_146 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_147 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_148 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_149 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_150 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_151 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_152 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_153 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_154 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_155 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_156 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_157 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_158 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_159 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_160 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_161 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_162 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_163 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_164 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_165 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_166 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_167 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_168 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_169 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_170 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_171 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_172 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_173 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_174 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_175 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_176 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_177 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_178 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_179 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_180 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_181 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_182 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_183 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_184 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_185 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_186 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_187 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_188 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_189 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_190 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_191 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_192 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_89 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_90 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_91 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_92 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_93 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_193 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_194 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_195 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_196 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_197 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_198 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_199 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_200 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_201 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_202 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_203 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_204 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_205 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_206 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_207 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_208 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_209 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_210 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_211 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_212 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_213 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_214 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_215 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_216 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_217 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_218 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_219 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_220 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_221 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_222 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_223 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_224 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_225 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_226 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_227 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_228 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_229 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_230 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_231 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_232 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_233 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_234 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_235 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_236 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_237 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_238 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_239 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_240 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_241 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_242 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_243 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_244 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_245 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_246 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_247 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_94 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_95 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_96 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_97 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_98 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_99 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_248 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_249 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_250 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_251 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_252 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_253 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_254 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_255 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_256 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_257 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_258 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_259 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_260 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_261 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_262 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_263 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_264 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_265 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_266 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_267 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_268 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_269 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_270 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_271 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_272 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_273 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_274 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_275 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_276 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_277 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_278 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_279 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_280 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_281 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_282 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_283 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_284 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_285 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_286 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_287 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_288 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_289 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_290 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_291 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_292 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_293 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_294 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_295 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_296 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_297 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_298 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_299 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_300 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_301 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_302 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_100 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_101 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_102 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_103 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_104 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_105 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_106 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_107 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_108 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_109 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_110 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_111 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_112 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_113 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_114 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_115 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_116 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_117 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_118 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_119 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_120 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_121 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_122 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_123 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_124 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_125 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_126 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_127 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_128 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_129 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_130 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_131 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_132 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_133 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_134 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_135 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_136 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_137 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__nor3_1 _211_ (.A(net3),
    .B(net2),
    .C(net6),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_000_));
 sky130_fd_sc_hd__buf_2 _212_ (.A(_000_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_001_));
 sky130_fd_sc_hd__and2b_1 _213_ (.A_N(net5),
    .B(net4),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_002_));
 sky130_fd_sc_hd__clkbuf_2 _214_ (.A(_002_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_003_));
 sky130_fd_sc_hd__and2_2 _215_ (.A(_001_),
    .B(_003_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_004_));
 sky130_fd_sc_hd__and2b_1 _216_ (.A_N(net2),
    .B(net3),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_005_));
 sky130_fd_sc_hd__nor3b_1 _217_ (.A(net5),
    .B(net4),
    .C_N(net6),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_006_));
 sky130_fd_sc_hd__clkbuf_2 _218_ (.A(_006_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_007_));
 sky130_fd_sc_hd__and2_2 _219_ (.A(_005_),
    .B(_007_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_008_));
 sky130_fd_sc_hd__nor2_1 _220_ (.A(net5),
    .B(net4),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_009_));
 sky130_fd_sc_hd__clkbuf_4 _221_ (.A(_009_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_010_));
 sky130_fd_sc_hd__nor3b_2 _222_ (.A(net3),
    .B(net6),
    .C_N(net2),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_011_));
 sky130_fd_sc_hd__clkbuf_4 _223_ (.A(_011_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_012_));
 sky130_fd_sc_hd__nor3b_1 _224_ (.A(net2),
    .B(net6),
    .C_N(net3),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_013_));
 sky130_fd_sc_hd__and2_2 _225_ (.A(_002_),
    .B(_013_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_014_));
 sky130_fd_sc_hd__a32o_1 _226_ (.A1(\tdc0.o_result[8] ),
    .A2(_010_),
    .A3(_012_),
    .B1(_014_),
    .B2(\tdc0.o_result[48] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_015_));
 sky130_fd_sc_hd__a221o_1 _227_ (.A1(\tdc0.o_result[32] ),
    .A2(_004_),
    .B1(_008_),
    .B2(\tdc0.o_result[144] ),
    .C1(_015_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_016_));
 sky130_fd_sc_hd__and2_2 _228_ (.A(_011_),
    .B(_003_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_017_));
 sky130_fd_sc_hd__and2b_1 _229_ (.A_N(net4),
    .B(net5),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_018_));
 sky130_fd_sc_hd__and3b_1 _230_ (.A_N(net6),
    .B(net2),
    .C(net3),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_019_));
 sky130_fd_sc_hd__and2_1 _231_ (.A(_018_),
    .B(_019_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_020_));
 sky130_fd_sc_hd__and2_1 _232_ (.A(net5),
    .B(net4),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_021_));
 sky130_fd_sc_hd__clkbuf_2 _233_ (.A(_021_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_022_));
 sky130_fd_sc_hd__and2_2 _234_ (.A(_022_),
    .B(_013_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_023_));
 sky130_fd_sc_hd__nor2_1 _235_ (.A(net3),
    .B(net2),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_024_));
 sky130_fd_sc_hd__clkbuf_2 _236_ (.A(_024_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_025_));
 sky130_fd_sc_hd__buf_2 _237_ (.A(_006_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_026_));
 sky130_fd_sc_hd__and2_1 _238_ (.A(_025_),
    .B(_026_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_027_));
 sky130_fd_sc_hd__a22o_1 _239_ (.A1(\tdc0.o_result[112] ),
    .A2(_023_),
    .B1(_027_),
    .B2(\tdc0.o_result[128] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_028_));
 sky130_fd_sc_hd__a221o_1 _240_ (.A1(\tdc0.o_result[40] ),
    .A2(_017_),
    .B1(_020_),
    .B2(\tdc0.o_result[88] ),
    .C1(_028_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_029_));
 sky130_fd_sc_hd__buf_2 _241_ (.A(_009_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_030_));
 sky130_fd_sc_hd__and2_2 _242_ (.A(_030_),
    .B(_019_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_031_));
 sky130_fd_sc_hd__and3_1 _243_ (.A(\tdc0.o_result[120] ),
    .B(_022_),
    .C(_019_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_032_));
 sky130_fd_sc_hd__a22o_2 _244_ (.A1(net5),
    .A2(net6),
    .B1(_000_),
    .B2(_030_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_033_));
 sky130_fd_sc_hd__clkbuf_2 _245_ (.A(_018_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_034_));
 sky130_fd_sc_hd__buf_2 _246_ (.A(_013_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_035_));
 sky130_fd_sc_hd__and3_1 _247_ (.A(\tdc0.o_result[80] ),
    .B(_034_),
    .C(_035_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_036_));
 sky130_fd_sc_hd__a2111o_1 _248_ (.A1(\tdc0.o_result[24] ),
    .A2(_031_),
    .B1(_032_),
    .C1(_033_),
    .D1(_036_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_037_));
 sky130_fd_sc_hd__and2b_2 _249_ (.A_N(net3),
    .B(net2),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_038_));
 sky130_fd_sc_hd__and2_2 _250_ (.A(_038_),
    .B(_007_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_039_));
 sky130_fd_sc_hd__and2_1 _251_ (.A(net3),
    .B(net2),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_040_));
 sky130_fd_sc_hd__and3_1 _252_ (.A(\tdc0.o_result[152] ),
    .B(_007_),
    .C(_040_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_041_));
 sky130_fd_sc_hd__and3b_1 _253_ (.A_N(net5),
    .B(net4),
    .C(net6),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_042_));
 sky130_fd_sc_hd__buf_2 _254_ (.A(_042_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_043_));
 sky130_fd_sc_hd__and3_1 _255_ (.A(\tdc0.o_result[160] ),
    .B(_025_),
    .C(_043_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_044_));
 sky130_fd_sc_hd__and3_1 _256_ (.A(\tdc0.o_result[16] ),
    .B(_010_),
    .C(_035_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_045_));
 sky130_fd_sc_hd__a2111o_1 _257_ (.A1(\tdc0.o_result[136] ),
    .A2(_039_),
    .B1(_041_),
    .C1(_044_),
    .D1(_045_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_046_));
 sky130_fd_sc_hd__and2_2 _258_ (.A(_022_),
    .B(_011_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_047_));
 sky130_fd_sc_hd__and3_1 _259_ (.A(\tdc0.o_result[96] ),
    .B(_001_),
    .C(_022_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_048_));
 sky130_fd_sc_hd__and3_1 _260_ (.A(\tdc0.o_result[64] ),
    .B(_001_),
    .C(_034_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_049_));
 sky130_fd_sc_hd__buf_2 _261_ (.A(_042_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_050_));
 sky130_fd_sc_hd__buf_2 _262_ (.A(_040_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_051_));
 sky130_fd_sc_hd__and3_1 _263_ (.A(\tdc0.o_result[184] ),
    .B(_050_),
    .C(_051_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_052_));
 sky130_fd_sc_hd__a2111o_1 _264_ (.A1(\tdc0.o_result[104] ),
    .A2(_047_),
    .B1(_048_),
    .C1(_049_),
    .D1(_052_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_053_));
 sky130_fd_sc_hd__buf_2 _265_ (.A(_019_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_054_));
 sky130_fd_sc_hd__and2_2 _266_ (.A(_003_),
    .B(_054_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_055_));
 sky130_fd_sc_hd__clkbuf_2 _267_ (.A(_042_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_056_));
 sky130_fd_sc_hd__and3_1 _268_ (.A(\tdc0.o_result[168] ),
    .B(_038_),
    .C(_056_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_057_));
 sky130_fd_sc_hd__clkbuf_2 _269_ (.A(_018_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_058_));
 sky130_fd_sc_hd__and3_1 _270_ (.A(\tdc0.o_result[72] ),
    .B(_012_),
    .C(_058_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_059_));
 sky130_fd_sc_hd__buf_2 _271_ (.A(_005_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_060_));
 sky130_fd_sc_hd__and3_1 _272_ (.A(\tdc0.o_result[176] ),
    .B(_060_),
    .C(_050_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_061_));
 sky130_fd_sc_hd__a2111o_1 _273_ (.A1(\tdc0.o_result[56] ),
    .A2(_055_),
    .B1(_057_),
    .C1(_059_),
    .D1(_061_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_062_));
 sky130_fd_sc_hd__or4_1 _274_ (.A(_037_),
    .B(_046_),
    .C(_053_),
    .D(_062_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_063_));
 sky130_fd_sc_hd__a22oi_4 _275_ (.A1(net5),
    .A2(net6),
    .B1(_001_),
    .B2(_010_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_064_));
 sky130_fd_sc_hd__o32a_4 _276_ (.A1(_016_),
    .A2(_029_),
    .A3(_063_),
    .B1(_064_),
    .B2(\tdc0.o_result[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[0]));
 sky130_fd_sc_hd__and2_2 _277_ (.A(_021_),
    .B(_019_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_065_));
 sky130_fd_sc_hd__a22o_1 _278_ (.A1(\tdc0.o_result[57] ),
    .A2(_055_),
    .B1(_065_),
    .B2(\tdc0.o_result[121] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_066_));
 sky130_fd_sc_hd__a221o_1 _279_ (.A1(\tdc0.o_result[41] ),
    .A2(_017_),
    .B1(_014_),
    .B2(\tdc0.o_result[49] ),
    .C1(_066_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_067_));
 sky130_fd_sc_hd__and2_1 _280_ (.A(_001_),
    .B(_058_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_068_));
 sky130_fd_sc_hd__and2_1 _281_ (.A(_043_),
    .B(_040_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_069_));
 sky130_fd_sc_hd__a32o_1 _282_ (.A1(\tdc0.o_result[9] ),
    .A2(_010_),
    .A3(_012_),
    .B1(_039_),
    .B2(\tdc0.o_result[137] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_070_));
 sky130_fd_sc_hd__a221o_1 _283_ (.A1(\tdc0.o_result[65] ),
    .A2(_068_),
    .B1(_069_),
    .B2(\tdc0.o_result[185] ),
    .C1(_070_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_071_));
 sky130_fd_sc_hd__and2_2 _284_ (.A(_001_),
    .B(_022_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_072_));
 sky130_fd_sc_hd__and3_1 _285_ (.A(\tdc0.o_result[169] ),
    .B(_038_),
    .C(_043_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_073_));
 sky130_fd_sc_hd__and3_1 _286_ (.A(\tdc0.o_result[89] ),
    .B(_034_),
    .C(_054_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_074_));
 sky130_fd_sc_hd__a2111o_1 _287_ (.A1(\tdc0.o_result[97] ),
    .A2(_072_),
    .B1(_073_),
    .C1(_074_),
    .D1(_033_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_075_));
 sky130_fd_sc_hd__buf_2 _288_ (.A(_013_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_076_));
 sky130_fd_sc_hd__and3_1 _289_ (.A(\tdc0.o_result[113] ),
    .B(_022_),
    .C(_076_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_077_));
 sky130_fd_sc_hd__and3_1 _290_ (.A(\tdc0.o_result[17] ),
    .B(_010_),
    .C(_076_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_078_));
 sky130_fd_sc_hd__and3_1 _291_ (.A(\tdc0.o_result[161] ),
    .B(_025_),
    .C(_056_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_079_));
 sky130_fd_sc_hd__a2111o_1 _292_ (.A1(\tdc0.o_result[25] ),
    .A2(_031_),
    .B1(_077_),
    .C1(_078_),
    .D1(_079_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_080_));
 sky130_fd_sc_hd__and3_1 _293_ (.A(\tdc0.o_result[105] ),
    .B(_022_),
    .C(_011_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_081_));
 sky130_fd_sc_hd__and3_1 _294_ (.A(\tdc0.o_result[177] ),
    .B(_060_),
    .C(_056_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_082_));
 sky130_fd_sc_hd__and3_1 _295_ (.A(\tdc0.o_result[145] ),
    .B(_060_),
    .C(_026_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_083_));
 sky130_fd_sc_hd__a2111o_1 _296_ (.A1(\tdc0.o_result[33] ),
    .A2(_004_),
    .B1(_081_),
    .C1(_082_),
    .D1(_083_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_084_));
 sky130_fd_sc_hd__and2_2 _297_ (.A(_012_),
    .B(_034_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_085_));
 sky130_fd_sc_hd__and3_1 _298_ (.A(\tdc0.o_result[81] ),
    .B(_034_),
    .C(_076_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_086_));
 sky130_fd_sc_hd__and3_1 _299_ (.A(\tdc0.o_result[129] ),
    .B(_025_),
    .C(_026_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_087_));
 sky130_fd_sc_hd__and3_1 _300_ (.A(\tdc0.o_result[153] ),
    .B(_026_),
    .C(_051_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_088_));
 sky130_fd_sc_hd__a2111o_1 _301_ (.A1(\tdc0.o_result[73] ),
    .A2(_085_),
    .B1(_086_),
    .C1(_087_),
    .D1(_088_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_089_));
 sky130_fd_sc_hd__or4_1 _302_ (.A(_075_),
    .B(_080_),
    .C(_084_),
    .D(_089_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_090_));
 sky130_fd_sc_hd__o32a_4 _303_ (.A1(_067_),
    .A2(_071_),
    .A3(_090_),
    .B1(_064_),
    .B2(\tdc0.o_result[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[1]));
 sky130_fd_sc_hd__a32o_1 _304_ (.A1(\tdc0.o_result[82] ),
    .A2(_058_),
    .A3(_035_),
    .B1(_004_),
    .B2(\tdc0.o_result[34] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_091_));
 sky130_fd_sc_hd__a221o_1 _305_ (.A1(\tdc0.o_result[98] ),
    .A2(_072_),
    .B1(_023_),
    .B2(\tdc0.o_result[114] ),
    .C1(_091_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_092_));
 sky130_fd_sc_hd__a22o_1 _306_ (.A1(\tdc0.o_result[106] ),
    .A2(_047_),
    .B1(_085_),
    .B2(\tdc0.o_result[74] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_093_));
 sky130_fd_sc_hd__a221o_1 _307_ (.A1(\tdc0.o_result[42] ),
    .A2(_017_),
    .B1(_008_),
    .B2(\tdc0.o_result[146] ),
    .C1(_093_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_094_));
 sky130_fd_sc_hd__and3_1 _308_ (.A(\tdc0.o_result[58] ),
    .B(_002_),
    .C(_019_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_095_));
 sky130_fd_sc_hd__and3_1 _309_ (.A(\tdc0.o_result[18] ),
    .B(_030_),
    .C(_076_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_096_));
 sky130_fd_sc_hd__a2111o_1 _310_ (.A1(\tdc0.o_result[122] ),
    .A2(_065_),
    .B1(_095_),
    .C1(_096_),
    .D1(_033_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_097_));
 sky130_fd_sc_hd__and3_1 _311_ (.A(\tdc0.o_result[162] ),
    .B(_024_),
    .C(_043_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_098_));
 sky130_fd_sc_hd__and3_1 _312_ (.A(\tdc0.o_result[130] ),
    .B(_025_),
    .C(_007_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_099_));
 sky130_fd_sc_hd__and3_1 _313_ (.A(\tdc0.o_result[90] ),
    .B(_058_),
    .C(_054_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_100_));
 sky130_fd_sc_hd__a2111o_1 _314_ (.A1(\tdc0.o_result[50] ),
    .A2(_014_),
    .B1(_098_),
    .C1(_099_),
    .D1(_100_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_101_));
 sky130_fd_sc_hd__and3_1 _315_ (.A(\tdc0.o_result[154] ),
    .B(_007_),
    .C(_040_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_102_));
 sky130_fd_sc_hd__and3_1 _316_ (.A(\tdc0.o_result[178] ),
    .B(_060_),
    .C(_056_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_103_));
 sky130_fd_sc_hd__and3_1 _317_ (.A(\tdc0.o_result[170] ),
    .B(_038_),
    .C(_050_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_104_));
 sky130_fd_sc_hd__a2111o_1 _318_ (.A1(\tdc0.o_result[138] ),
    .A2(_039_),
    .B1(_102_),
    .C1(_103_),
    .D1(_104_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_105_));
 sky130_fd_sc_hd__and3_1 _319_ (.A(\tdc0.o_result[10] ),
    .B(_010_),
    .C(_012_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_106_));
 sky130_fd_sc_hd__and3_1 _320_ (.A(\tdc0.o_result[66] ),
    .B(_001_),
    .C(_058_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_107_));
 sky130_fd_sc_hd__and3_1 _321_ (.A(\tdc0.o_result[186] ),
    .B(_050_),
    .C(_051_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_108_));
 sky130_fd_sc_hd__a2111o_1 _322_ (.A1(\tdc0.o_result[26] ),
    .A2(_031_),
    .B1(_106_),
    .C1(_107_),
    .D1(_108_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_109_));
 sky130_fd_sc_hd__or4_1 _323_ (.A(_097_),
    .B(_101_),
    .C(_105_),
    .D(_109_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_110_));
 sky130_fd_sc_hd__o32a_4 _324_ (.A1(_092_),
    .A2(_094_),
    .A3(_110_),
    .B1(_064_),
    .B2(\tdc0.o_result[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[2]));
 sky130_fd_sc_hd__a32o_1 _325_ (.A1(\tdc0.o_result[11] ),
    .A2(_010_),
    .A3(_012_),
    .B1(_047_),
    .B2(\tdc0.o_result[107] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_111_));
 sky130_fd_sc_hd__a221o_1 _326_ (.A1(\tdc0.o_result[99] ),
    .A2(_072_),
    .B1(_055_),
    .B2(\tdc0.o_result[59] ),
    .C1(_111_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_112_));
 sky130_fd_sc_hd__a32o_1 _327_ (.A1(\tdc0.o_result[155] ),
    .A2(_026_),
    .A3(_051_),
    .B1(_068_),
    .B2(\tdc0.o_result[67] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_113_));
 sky130_fd_sc_hd__a221o_1 _328_ (.A1(\tdc0.o_result[75] ),
    .A2(_085_),
    .B1(_031_),
    .B2(\tdc0.o_result[27] ),
    .C1(_113_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_114_));
 sky130_fd_sc_hd__and3_1 _329_ (.A(\tdc0.o_result[19] ),
    .B(_030_),
    .C(_076_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_115_));
 sky130_fd_sc_hd__and3_1 _330_ (.A(\tdc0.o_result[163] ),
    .B(_025_),
    .C(_043_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_116_));
 sky130_fd_sc_hd__a2111o_1 _331_ (.A1(\tdc0.o_result[91] ),
    .A2(_020_),
    .B1(_115_),
    .C1(_116_),
    .D1(_033_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_117_));
 sky130_fd_sc_hd__and3_1 _332_ (.A(\tdc0.o_result[43] ),
    .B(_011_),
    .C(_003_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_118_));
 sky130_fd_sc_hd__and3_1 _333_ (.A(\tdc0.o_result[123] ),
    .B(_022_),
    .C(_054_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_119_));
 sky130_fd_sc_hd__and3_1 _334_ (.A(\tdc0.o_result[83] ),
    .B(_058_),
    .C(_035_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_120_));
 sky130_fd_sc_hd__a2111o_1 _335_ (.A1(\tdc0.o_result[139] ),
    .A2(_039_),
    .B1(_118_),
    .C1(_119_),
    .D1(_120_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_121_));
 sky130_fd_sc_hd__and3_1 _336_ (.A(\tdc0.o_result[147] ),
    .B(_060_),
    .C(_007_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_122_));
 sky130_fd_sc_hd__and3_1 _337_ (.A(\tdc0.o_result[171] ),
    .B(_038_),
    .C(_056_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_123_));
 sky130_fd_sc_hd__and3_1 _338_ (.A(\tdc0.o_result[131] ),
    .B(_025_),
    .C(_026_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_124_));
 sky130_fd_sc_hd__a2111o_1 _339_ (.A1(\tdc0.o_result[115] ),
    .A2(_023_),
    .B1(_122_),
    .C1(_123_),
    .D1(_124_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_125_));
 sky130_fd_sc_hd__and3_1 _340_ (.A(\tdc0.o_result[187] ),
    .B(_056_),
    .C(_051_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_126_));
 sky130_fd_sc_hd__and3_1 _341_ (.A(\tdc0.o_result[51] ),
    .B(_003_),
    .C(_035_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_127_));
 sky130_fd_sc_hd__and3_1 _342_ (.A(\tdc0.o_result[179] ),
    .B(_060_),
    .C(_050_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_128_));
 sky130_fd_sc_hd__a2111o_1 _343_ (.A1(\tdc0.o_result[35] ),
    .A2(_004_),
    .B1(_126_),
    .C1(_127_),
    .D1(_128_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_129_));
 sky130_fd_sc_hd__or4_1 _344_ (.A(_117_),
    .B(_121_),
    .C(_125_),
    .D(_129_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_130_));
 sky130_fd_sc_hd__o32a_4 _345_ (.A1(_112_),
    .A2(_114_),
    .A3(_130_),
    .B1(_064_),
    .B2(\tdc0.o_result[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[3]));
 sky130_fd_sc_hd__a22o_1 _346_ (.A1(\tdc0.o_result[108] ),
    .A2(_047_),
    .B1(_027_),
    .B2(\tdc0.o_result[132] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_131_));
 sky130_fd_sc_hd__a221o_1 _347_ (.A1(\tdc0.o_result[100] ),
    .A2(_072_),
    .B1(_023_),
    .B2(\tdc0.o_result[116] ),
    .C1(_131_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_132_));
 sky130_fd_sc_hd__a32o_1 _348_ (.A1(\tdc0.o_result[180] ),
    .A2(_060_),
    .A3(_050_),
    .B1(_031_),
    .B2(\tdc0.o_result[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_133_));
 sky130_fd_sc_hd__a221o_1 _349_ (.A1(\tdc0.o_result[76] ),
    .A2(_085_),
    .B1(_020_),
    .B2(\tdc0.o_result[92] ),
    .C1(_133_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_134_));
 sky130_fd_sc_hd__and3_1 _350_ (.A(\tdc0.o_result[164] ),
    .B(_024_),
    .C(_043_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_135_));
 sky130_fd_sc_hd__and3_1 _351_ (.A(\tdc0.o_result[20] ),
    .B(_030_),
    .C(_076_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_136_));
 sky130_fd_sc_hd__a2111o_1 _352_ (.A1(\tdc0.o_result[188] ),
    .A2(_069_),
    .B1(_135_),
    .C1(_136_),
    .D1(_033_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_137_));
 sky130_fd_sc_hd__and3_1 _353_ (.A(\tdc0.o_result[84] ),
    .B(_034_),
    .C(_076_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_138_));
 sky130_fd_sc_hd__and3_1 _354_ (.A(\tdc0.o_result[124] ),
    .B(_022_),
    .C(_054_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_139_));
 sky130_fd_sc_hd__and3_1 _355_ (.A(\tdc0.o_result[60] ),
    .B(_003_),
    .C(_054_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_140_));
 sky130_fd_sc_hd__a2111o_1 _356_ (.A1(\tdc0.o_result[140] ),
    .A2(_039_),
    .B1(_138_),
    .C1(_139_),
    .D1(_140_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_141_));
 sky130_fd_sc_hd__and3_1 _357_ (.A(\tdc0.o_result[12] ),
    .B(_030_),
    .C(_011_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_142_));
 sky130_fd_sc_hd__and3_1 _358_ (.A(\tdc0.o_result[156] ),
    .B(_026_),
    .C(_051_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_143_));
 sky130_fd_sc_hd__and3_1 _359_ (.A(\tdc0.o_result[172] ),
    .B(_038_),
    .C(_050_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_144_));
 sky130_fd_sc_hd__a2111o_1 _360_ (.A1(\tdc0.o_result[148] ),
    .A2(_008_),
    .B1(_142_),
    .C1(_143_),
    .D1(_144_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_145_));
 sky130_fd_sc_hd__and3_1 _361_ (.A(\tdc0.o_result[44] ),
    .B(_012_),
    .C(_003_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_146_));
 sky130_fd_sc_hd__and3_1 _362_ (.A(\tdc0.o_result[52] ),
    .B(_003_),
    .C(_035_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_147_));
 sky130_fd_sc_hd__and3_1 _363_ (.A(\tdc0.o_result[68] ),
    .B(_001_),
    .C(_058_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_148_));
 sky130_fd_sc_hd__a2111o_1 _364_ (.A1(\tdc0.o_result[36] ),
    .A2(_004_),
    .B1(_146_),
    .C1(_147_),
    .D1(_148_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_149_));
 sky130_fd_sc_hd__or4_1 _365_ (.A(_137_),
    .B(_141_),
    .C(_145_),
    .D(_149_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_150_));
 sky130_fd_sc_hd__o32a_4 _366_ (.A1(_132_),
    .A2(_134_),
    .A3(_150_),
    .B1(_064_),
    .B2(\tdc0.o_result[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[4]));
 sky130_fd_sc_hd__a22o_1 _367_ (.A1(\tdc0.o_result[69] ),
    .A2(_068_),
    .B1(_065_),
    .B2(\tdc0.o_result[125] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_151_));
 sky130_fd_sc_hd__a221o_1 _368_ (.A1(\tdc0.o_result[45] ),
    .A2(_017_),
    .B1(_014_),
    .B2(\tdc0.o_result[53] ),
    .C1(_151_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_152_));
 sky130_fd_sc_hd__a32o_1 _369_ (.A1(\tdc0.o_result[165] ),
    .A2(_025_),
    .A3(_050_),
    .B1(_039_),
    .B2(\tdc0.o_result[141] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_153_));
 sky130_fd_sc_hd__a221o_1 _370_ (.A1(\tdc0.o_result[61] ),
    .A2(_055_),
    .B1(_004_),
    .B2(\tdc0.o_result[37] ),
    .C1(_153_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_154_));
 sky130_fd_sc_hd__and3_1 _371_ (.A(\tdc0.o_result[133] ),
    .B(_024_),
    .C(_007_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_155_));
 sky130_fd_sc_hd__and3_1 _372_ (.A(\tdc0.o_result[85] ),
    .B(_034_),
    .C(_076_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_156_));
 sky130_fd_sc_hd__a2111o_1 _373_ (.A1(\tdc0.o_result[117] ),
    .A2(_023_),
    .B1(_155_),
    .C1(_156_),
    .D1(_033_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_157_));
 sky130_fd_sc_hd__and3_1 _374_ (.A(\tdc0.o_result[13] ),
    .B(_030_),
    .C(_011_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_158_));
 sky130_fd_sc_hd__and3_1 _375_ (.A(\tdc0.o_result[29] ),
    .B(_030_),
    .C(_054_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_159_));
 sky130_fd_sc_hd__and3_1 _376_ (.A(\tdc0.o_result[21] ),
    .B(_010_),
    .C(_035_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_160_));
 sky130_fd_sc_hd__a2111o_1 _377_ (.A1(\tdc0.o_result[101] ),
    .A2(_072_),
    .B1(_158_),
    .C1(_159_),
    .D1(_160_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_161_));
 sky130_fd_sc_hd__and3_1 _378_ (.A(\tdc0.o_result[181] ),
    .B(_005_),
    .C(_043_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_162_));
 sky130_fd_sc_hd__and3_1 _379_ (.A(\tdc0.o_result[189] ),
    .B(_056_),
    .C(_051_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_163_));
 sky130_fd_sc_hd__and3_1 _380_ (.A(\tdc0.o_result[149] ),
    .B(_060_),
    .C(_026_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_164_));
 sky130_fd_sc_hd__a2111o_1 _381_ (.A1(\tdc0.o_result[109] ),
    .A2(_047_),
    .B1(_162_),
    .C1(_163_),
    .D1(_164_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_165_));
 sky130_fd_sc_hd__and3_1 _382_ (.A(\tdc0.o_result[93] ),
    .B(_034_),
    .C(_054_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_166_));
 sky130_fd_sc_hd__and3_1 _383_ (.A(\tdc0.o_result[157] ),
    .B(_026_),
    .C(_051_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_167_));
 sky130_fd_sc_hd__and3_1 _384_ (.A(\tdc0.o_result[173] ),
    .B(_038_),
    .C(_050_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_168_));
 sky130_fd_sc_hd__a2111o_1 _385_ (.A1(\tdc0.o_result[77] ),
    .A2(_085_),
    .B1(_166_),
    .C1(_167_),
    .D1(_168_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_169_));
 sky130_fd_sc_hd__or4_1 _386_ (.A(_157_),
    .B(_161_),
    .C(_165_),
    .D(_169_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_170_));
 sky130_fd_sc_hd__o32a_4 _387_ (.A1(_152_),
    .A2(_154_),
    .A3(_170_),
    .B1(_064_),
    .B2(\tdc0.o_result[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[5]));
 sky130_fd_sc_hd__a22o_1 _388_ (.A1(\tdc0.o_result[110] ),
    .A2(_047_),
    .B1(_008_),
    .B2(\tdc0.o_result[150] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_171_));
 sky130_fd_sc_hd__a221o_1 _389_ (.A1(\tdc0.o_result[102] ),
    .A2(_072_),
    .B1(_023_),
    .B2(\tdc0.o_result[118] ),
    .C1(_171_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_172_));
 sky130_fd_sc_hd__a32o_1 _390_ (.A1(\tdc0.o_result[86] ),
    .A2(_058_),
    .A3(_035_),
    .B1(_020_),
    .B2(\tdc0.o_result[94] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_173_));
 sky130_fd_sc_hd__a221o_1 _391_ (.A1(\tdc0.o_result[142] ),
    .A2(_039_),
    .B1(_004_),
    .B2(\tdc0.o_result[38] ),
    .C1(_173_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_174_));
 sky130_fd_sc_hd__and3_1 _392_ (.A(\tdc0.o_result[70] ),
    .B(_001_),
    .C(_018_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_175_));
 sky130_fd_sc_hd__and3_1 _393_ (.A(\tdc0.o_result[190] ),
    .B(_043_),
    .C(_051_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_176_));
 sky130_fd_sc_hd__a2111o_1 _394_ (.A1(\tdc0.o_result[54] ),
    .A2(_014_),
    .B1(_175_),
    .C1(_176_),
    .D1(_033_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_177_));
 sky130_fd_sc_hd__and3_1 _395_ (.A(\tdc0.o_result[134] ),
    .B(_024_),
    .C(_007_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_178_));
 sky130_fd_sc_hd__and3_1 _396_ (.A(\tdc0.o_result[166] ),
    .B(_025_),
    .C(_043_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_179_));
 sky130_fd_sc_hd__and3_1 _397_ (.A(\tdc0.o_result[78] ),
    .B(_012_),
    .C(_058_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_180_));
 sky130_fd_sc_hd__a2111o_1 _398_ (.A1(\tdc0.o_result[126] ),
    .A2(_065_),
    .B1(_178_),
    .C1(_179_),
    .D1(_180_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_181_));
 sky130_fd_sc_hd__and3_1 _399_ (.A(\tdc0.o_result[158] ),
    .B(_007_),
    .C(_040_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_182_));
 sky130_fd_sc_hd__and3_1 _400_ (.A(\tdc0.o_result[182] ),
    .B(_060_),
    .C(_056_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_183_));
 sky130_fd_sc_hd__and3_1 _401_ (.A(\tdc0.o_result[174] ),
    .B(_038_),
    .C(_056_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_184_));
 sky130_fd_sc_hd__a2111o_1 _402_ (.A1(\tdc0.o_result[46] ),
    .A2(_017_),
    .B1(_182_),
    .C1(_183_),
    .D1(_184_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_185_));
 sky130_fd_sc_hd__and3_1 _403_ (.A(\tdc0.o_result[14] ),
    .B(_010_),
    .C(_012_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_186_));
 sky130_fd_sc_hd__and3_1 _404_ (.A(\tdc0.o_result[62] ),
    .B(_003_),
    .C(_054_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_187_));
 sky130_fd_sc_hd__and3_1 _405_ (.A(\tdc0.o_result[22] ),
    .B(_010_),
    .C(_035_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_188_));
 sky130_fd_sc_hd__a2111o_1 _406_ (.A1(\tdc0.o_result[30] ),
    .A2(_031_),
    .B1(_186_),
    .C1(_187_),
    .D1(_188_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_189_));
 sky130_fd_sc_hd__or4_1 _407_ (.A(_177_),
    .B(_181_),
    .C(_185_),
    .D(_189_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_190_));
 sky130_fd_sc_hd__o32a_4 _408_ (.A1(_172_),
    .A2(_174_),
    .A3(_190_),
    .B1(_064_),
    .B2(\tdc0.o_result[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[6]));
 sky130_fd_sc_hd__a22o_1 _409_ (.A1(\tdc0.o_result[79] ),
    .A2(_085_),
    .B1(_027_),
    .B2(\tdc0.o_result[135] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_191_));
 sky130_fd_sc_hd__a221o_1 _410_ (.A1(\tdc0.o_result[103] ),
    .A2(_072_),
    .B1(_023_),
    .B2(\tdc0.o_result[119] ),
    .C1(_191_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_192_));
 sky130_fd_sc_hd__a32o_1 _411_ (.A1(\tdc0.o_result[183] ),
    .A2(_060_),
    .A3(_050_),
    .B1(_031_),
    .B2(\tdc0.o_result[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_193_));
 sky130_fd_sc_hd__a221o_1 _412_ (.A1(\tdc0.o_result[47] ),
    .A2(_017_),
    .B1(_055_),
    .B2(\tdc0.o_result[63] ),
    .C1(_193_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_194_));
 sky130_fd_sc_hd__and3_1 _413_ (.A(\tdc0.o_result[143] ),
    .B(_038_),
    .C(_007_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_195_));
 sky130_fd_sc_hd__and3_1 _414_ (.A(\tdc0.o_result[23] ),
    .B(_030_),
    .C(_076_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_196_));
 sky130_fd_sc_hd__a2111o_1 _415_ (.A1(\tdc0.o_result[191] ),
    .A2(_069_),
    .B1(_195_),
    .C1(_196_),
    .D1(_033_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_197_));
 sky130_fd_sc_hd__and3_1 _416_ (.A(\tdc0.o_result[87] ),
    .B(_034_),
    .C(_076_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_198_));
 sky130_fd_sc_hd__and3_1 _417_ (.A(\tdc0.o_result[167] ),
    .B(_025_),
    .C(_043_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_199_));
 sky130_fd_sc_hd__and3_1 _418_ (.A(\tdc0.o_result[71] ),
    .B(_001_),
    .C(_034_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_200_));
 sky130_fd_sc_hd__a2111o_1 _419_ (.A1(\tdc0.o_result[127] ),
    .A2(_065_),
    .B1(_198_),
    .C1(_199_),
    .D1(_200_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_201_));
 sky130_fd_sc_hd__and3_1 _420_ (.A(\tdc0.o_result[15] ),
    .B(_030_),
    .C(_011_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_202_));
 sky130_fd_sc_hd__and3_1 _421_ (.A(\tdc0.o_result[159] ),
    .B(_026_),
    .C(_051_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_203_));
 sky130_fd_sc_hd__and3_1 _422_ (.A(\tdc0.o_result[175] ),
    .B(_038_),
    .C(_056_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_204_));
 sky130_fd_sc_hd__a2111o_1 _423_ (.A1(\tdc0.o_result[151] ),
    .A2(_008_),
    .B1(_202_),
    .C1(_203_),
    .D1(_204_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_205_));
 sky130_fd_sc_hd__and3_1 _424_ (.A(\tdc0.o_result[111] ),
    .B(_022_),
    .C(_012_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_206_));
 sky130_fd_sc_hd__and3_1 _425_ (.A(\tdc0.o_result[55] ),
    .B(_003_),
    .C(_035_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_207_));
 sky130_fd_sc_hd__and3_1 _426_ (.A(\tdc0.o_result[95] ),
    .B(_058_),
    .C(_054_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_208_));
 sky130_fd_sc_hd__a2111o_1 _427_ (.A1(\tdc0.o_result[39] ),
    .A2(_004_),
    .B1(_206_),
    .C1(_207_),
    .D1(_208_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_209_));
 sky130_fd_sc_hd__or4_1 _428_ (.A(_197_),
    .B(_201_),
    .C(_205_),
    .D(_209_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_210_));
 sky130_fd_sc_hd__o32a_4 _429_ (.A1(_192_),
    .A2(_194_),
    .A3(_210_),
    .B1(_064_),
    .B2(\tdc0.o_result[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[7]));
 sky130_fd_sc_hd__dfxtp_1 _430_ (.CLK(clknet_4_15_0_clk),
    .D(\tdc0.w_dly_sig[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[0] ));
 sky130_fd_sc_hd__dfxtp_1 _431_ (.CLK(clknet_4_15_0_clk),
    .D(\tdc0.w_dly_sig[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[1] ));
 sky130_fd_sc_hd__dfxtp_1 _432_ (.CLK(clknet_4_15_0_clk),
    .D(\tdc0.w_dly_sig[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[2] ));
 sky130_fd_sc_hd__dfxtp_1 _433_ (.CLK(clknet_4_15_0_clk),
    .D(\tdc0.w_dly_sig[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[3] ));
 sky130_fd_sc_hd__dfxtp_1 _434_ (.CLK(clknet_4_7_0_clk),
    .D(net23),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[4] ));
 sky130_fd_sc_hd__dfxtp_1 _435_ (.CLK(clknet_4_15_0_clk),
    .D(\tdc0.w_dly_sig[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[5] ));
 sky130_fd_sc_hd__dfxtp_1 _436_ (.CLK(clknet_4_15_0_clk),
    .D(\tdc0.w_dly_sig[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[6] ));
 sky130_fd_sc_hd__dfxtp_1 _437_ (.CLK(clknet_4_15_0_clk),
    .D(\tdc0.w_dly_sig[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[7] ));
 sky130_fd_sc_hd__dfxtp_1 _438_ (.CLK(clknet_4_15_0_clk),
    .D(\tdc0.w_dly_sig[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[8] ));
 sky130_fd_sc_hd__dfxtp_1 _439_ (.CLK(clknet_4_15_0_clk),
    .D(\tdc0.w_dly_sig[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[9] ));
 sky130_fd_sc_hd__dfxtp_1 _440_ (.CLK(clknet_4_15_0_clk),
    .D(\tdc0.w_dly_sig[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[10] ));
 sky130_fd_sc_hd__dfxtp_1 _441_ (.CLK(clknet_4_15_0_clk),
    .D(\tdc0.w_dly_sig[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[11] ));
 sky130_fd_sc_hd__dfxtp_1 _442_ (.CLK(clknet_4_14_0_clk),
    .D(\tdc0.w_dly_sig[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[12] ));
 sky130_fd_sc_hd__dfxtp_1 _443_ (.CLK(clknet_4_14_0_clk),
    .D(\tdc0.w_dly_sig[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[13] ));
 sky130_fd_sc_hd__dfxtp_1 _444_ (.CLK(clknet_4_14_0_clk),
    .D(\tdc0.w_dly_sig[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[14] ));
 sky130_fd_sc_hd__dfxtp_1 _445_ (.CLK(clknet_4_14_0_clk),
    .D(\tdc0.w_dly_sig[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[15] ));
 sky130_fd_sc_hd__dfxtp_1 _446_ (.CLK(clknet_4_14_0_clk),
    .D(net26),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[16] ));
 sky130_fd_sc_hd__dfxtp_1 _447_ (.CLK(clknet_4_11_0_clk),
    .D(net25),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[17] ));
 sky130_fd_sc_hd__dfxtp_1 _448_ (.CLK(clknet_4_14_0_clk),
    .D(\tdc0.w_dly_sig[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[18] ));
 sky130_fd_sc_hd__dfxtp_1 _449_ (.CLK(clknet_4_14_0_clk),
    .D(net27),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[19] ));
 sky130_fd_sc_hd__dfxtp_1 _450_ (.CLK(clknet_4_11_0_clk),
    .D(\tdc0.w_dly_sig[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[20] ));
 sky130_fd_sc_hd__dfxtp_1 _451_ (.CLK(clknet_4_14_0_clk),
    .D(net24),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[21] ));
 sky130_fd_sc_hd__dfxtp_1 _452_ (.CLK(clknet_4_14_0_clk),
    .D(\tdc0.w_dly_sig[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[22] ));
 sky130_fd_sc_hd__dfxtp_1 _453_ (.CLK(clknet_4_11_0_clk),
    .D(\tdc0.w_dly_sig[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[23] ));
 sky130_fd_sc_hd__dfxtp_1 _454_ (.CLK(clknet_4_11_0_clk),
    .D(\tdc0.w_dly_sig[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[24] ));
 sky130_fd_sc_hd__dfxtp_1 _455_ (.CLK(clknet_4_11_0_clk),
    .D(\tdc0.w_dly_sig[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[25] ));
 sky130_fd_sc_hd__dfxtp_1 _456_ (.CLK(clknet_4_11_0_clk),
    .D(\tdc0.w_dly_sig[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[26] ));
 sky130_fd_sc_hd__dfxtp_1 _457_ (.CLK(clknet_4_10_0_clk),
    .D(\tdc0.w_dly_sig[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[27] ));
 sky130_fd_sc_hd__dfxtp_1 _458_ (.CLK(clknet_4_10_0_clk),
    .D(\tdc0.w_dly_sig[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[28] ));
 sky130_fd_sc_hd__dfxtp_1 _459_ (.CLK(clknet_4_11_0_clk),
    .D(\tdc0.w_dly_sig[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[29] ));
 sky130_fd_sc_hd__dfxtp_1 _460_ (.CLK(clknet_4_11_0_clk),
    .D(\tdc0.w_dly_sig[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[30] ));
 sky130_fd_sc_hd__dfxtp_1 _461_ (.CLK(clknet_4_10_0_clk),
    .D(\tdc0.w_dly_sig[32] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[31] ));
 sky130_fd_sc_hd__dfxtp_1 _462_ (.CLK(clknet_4_12_0_clk),
    .D(\tdc0.w_dly_sig[33] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[32] ));
 sky130_fd_sc_hd__dfxtp_1 _463_ (.CLK(clknet_4_14_0_clk),
    .D(\tdc0.w_dly_sig[34] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[33] ));
 sky130_fd_sc_hd__dfxtp_1 _464_ (.CLK(clknet_4_12_0_clk),
    .D(\tdc0.w_dly_sig[35] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[34] ));
 sky130_fd_sc_hd__dfxtp_1 _465_ (.CLK(clknet_4_14_0_clk),
    .D(\tdc0.w_dly_sig[36] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[35] ));
 sky130_fd_sc_hd__dfxtp_1 _466_ (.CLK(clknet_4_12_0_clk),
    .D(\tdc0.w_dly_sig[37] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[36] ));
 sky130_fd_sc_hd__dfxtp_1 _467_ (.CLK(clknet_4_12_0_clk),
    .D(\tdc0.w_dly_sig[38] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[37] ));
 sky130_fd_sc_hd__dfxtp_1 _468_ (.CLK(clknet_4_13_0_clk),
    .D(\tdc0.w_dly_sig[39] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[38] ));
 sky130_fd_sc_hd__dfxtp_1 _469_ (.CLK(clknet_4_7_0_clk),
    .D(\tdc0.w_dly_sig[40] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[39] ));
 sky130_fd_sc_hd__dfxtp_1 _470_ (.CLK(clknet_4_13_0_clk),
    .D(\tdc0.w_dly_sig[41] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[40] ));
 sky130_fd_sc_hd__dfxtp_1 _471_ (.CLK(clknet_4_12_0_clk),
    .D(\tdc0.w_dly_sig[42] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[41] ));
 sky130_fd_sc_hd__dfxtp_1 _472_ (.CLK(clknet_4_13_0_clk),
    .D(\tdc0.w_dly_sig[43] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[42] ));
 sky130_fd_sc_hd__dfxtp_1 _473_ (.CLK(clknet_4_13_0_clk),
    .D(\tdc0.w_dly_sig[44] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[43] ));
 sky130_fd_sc_hd__dfxtp_1 _474_ (.CLK(clknet_4_12_0_clk),
    .D(\tdc0.w_dly_sig[45] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[44] ));
 sky130_fd_sc_hd__dfxtp_1 _475_ (.CLK(clknet_4_12_0_clk),
    .D(\tdc0.w_dly_sig[46] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[45] ));
 sky130_fd_sc_hd__dfxtp_1 _476_ (.CLK(clknet_4_15_0_clk),
    .D(\tdc0.w_dly_sig[47] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[46] ));
 sky130_fd_sc_hd__dfxtp_1 _477_ (.CLK(clknet_4_15_0_clk),
    .D(\tdc0.w_dly_sig[48] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[47] ));
 sky130_fd_sc_hd__dfxtp_1 _478_ (.CLK(clknet_4_15_0_clk),
    .D(\tdc0.w_dly_sig[49] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[48] ));
 sky130_fd_sc_hd__dfxtp_1 _479_ (.CLK(clknet_4_15_0_clk),
    .D(\tdc0.w_dly_sig[50] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[49] ));
 sky130_fd_sc_hd__dfxtp_1 _480_ (.CLK(clknet_4_13_0_clk),
    .D(\tdc0.w_dly_sig[51] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[50] ));
 sky130_fd_sc_hd__dfxtp_1 _481_ (.CLK(clknet_4_15_0_clk),
    .D(\tdc0.w_dly_sig[52] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[51] ));
 sky130_fd_sc_hd__dfxtp_1 _482_ (.CLK(clknet_4_12_0_clk),
    .D(\tdc0.w_dly_sig[53] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[52] ));
 sky130_fd_sc_hd__dfxtp_1 _483_ (.CLK(clknet_4_13_0_clk),
    .D(\tdc0.w_dly_sig[54] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[53] ));
 sky130_fd_sc_hd__dfxtp_1 _484_ (.CLK(clknet_4_13_0_clk),
    .D(\tdc0.w_dly_sig[55] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[54] ));
 sky130_fd_sc_hd__dfxtp_1 _485_ (.CLK(clknet_4_7_0_clk),
    .D(\tdc0.w_dly_sig[56] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[55] ));
 sky130_fd_sc_hd__dfxtp_1 _486_ (.CLK(clknet_4_7_0_clk),
    .D(\tdc0.w_dly_sig[57] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[56] ));
 sky130_fd_sc_hd__dfxtp_1 _487_ (.CLK(clknet_4_13_0_clk),
    .D(\tdc0.w_dly_sig[58] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[57] ));
 sky130_fd_sc_hd__dfxtp_1 _488_ (.CLK(clknet_4_13_0_clk),
    .D(\tdc0.w_dly_sig[59] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[58] ));
 sky130_fd_sc_hd__dfxtp_1 _489_ (.CLK(clknet_4_7_0_clk),
    .D(\tdc0.w_dly_sig[60] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[59] ));
 sky130_fd_sc_hd__dfxtp_1 _490_ (.CLK(clknet_4_7_0_clk),
    .D(\tdc0.w_dly_sig[61] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[60] ));
 sky130_fd_sc_hd__dfxtp_1 _491_ (.CLK(clknet_4_7_0_clk),
    .D(\tdc0.w_dly_sig[62] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[61] ));
 sky130_fd_sc_hd__dfxtp_1 _492_ (.CLK(clknet_4_12_0_clk),
    .D(\tdc0.w_dly_sig[63] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[62] ));
 sky130_fd_sc_hd__dfxtp_1 _493_ (.CLK(clknet_4_13_0_clk),
    .D(\tdc0.w_dly_sig[64] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[63] ));
 sky130_fd_sc_hd__dfxtp_1 _494_ (.CLK(clknet_4_6_0_clk),
    .D(\tdc0.w_dly_sig[65] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[64] ));
 sky130_fd_sc_hd__dfxtp_1 _495_ (.CLK(clknet_4_9_0_clk),
    .D(\tdc0.w_dly_sig[66] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[65] ));
 sky130_fd_sc_hd__dfxtp_1 _496_ (.CLK(clknet_4_6_0_clk),
    .D(\tdc0.w_dly_sig[67] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[66] ));
 sky130_fd_sc_hd__dfxtp_1 _497_ (.CLK(clknet_4_3_0_clk),
    .D(\tdc0.w_dly_sig[68] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[67] ));
 sky130_fd_sc_hd__dfxtp_1 _498_ (.CLK(clknet_4_6_0_clk),
    .D(\tdc0.w_dly_sig[69] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[68] ));
 sky130_fd_sc_hd__dfxtp_1 _499_ (.CLK(clknet_4_3_0_clk),
    .D(\tdc0.w_dly_sig[70] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[69] ));
 sky130_fd_sc_hd__dfxtp_1 _500_ (.CLK(clknet_4_3_0_clk),
    .D(\tdc0.w_dly_sig[71] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[70] ));
 sky130_fd_sc_hd__dfxtp_1 _501_ (.CLK(clknet_4_3_0_clk),
    .D(\tdc0.w_dly_sig[72] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[71] ));
 sky130_fd_sc_hd__dfxtp_1 _502_ (.CLK(clknet_4_1_0_clk),
    .D(\tdc0.w_dly_sig[73] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[72] ));
 sky130_fd_sc_hd__dfxtp_1 _503_ (.CLK(clknet_4_1_0_clk),
    .D(\tdc0.w_dly_sig[74] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[73] ));
 sky130_fd_sc_hd__dfxtp_1 _504_ (.CLK(clknet_4_4_0_clk),
    .D(\tdc0.w_dly_sig[75] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[74] ));
 sky130_fd_sc_hd__dfxtp_1 _505_ (.CLK(clknet_4_1_0_clk),
    .D(\tdc0.w_dly_sig[76] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[75] ));
 sky130_fd_sc_hd__dfxtp_1 _506_ (.CLK(clknet_4_1_0_clk),
    .D(\tdc0.w_dly_sig[77] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[76] ));
 sky130_fd_sc_hd__dfxtp_1 _507_ (.CLK(clknet_4_1_0_clk),
    .D(\tdc0.w_dly_sig[78] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[77] ));
 sky130_fd_sc_hd__dfxtp_1 _508_ (.CLK(clknet_4_1_0_clk),
    .D(\tdc0.w_dly_sig[79] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[78] ));
 sky130_fd_sc_hd__dfxtp_1 _509_ (.CLK(clknet_4_1_0_clk),
    .D(\tdc0.w_dly_sig[80] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[79] ));
 sky130_fd_sc_hd__dfxtp_1 _510_ (.CLK(clknet_4_1_0_clk),
    .D(\tdc0.w_dly_sig[81] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[80] ));
 sky130_fd_sc_hd__dfxtp_1 _511_ (.CLK(clknet_4_1_0_clk),
    .D(\tdc0.w_dly_sig[82] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[81] ));
 sky130_fd_sc_hd__dfxtp_1 _512_ (.CLK(clknet_4_4_0_clk),
    .D(\tdc0.w_dly_sig[83] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[82] ));
 sky130_fd_sc_hd__dfxtp_1 _513_ (.CLK(clknet_4_4_0_clk),
    .D(\tdc0.w_dly_sig[84] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[83] ));
 sky130_fd_sc_hd__dfxtp_1 _514_ (.CLK(clknet_4_4_0_clk),
    .D(\tdc0.w_dly_sig[85] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[84] ));
 sky130_fd_sc_hd__dfxtp_1 _515_ (.CLK(clknet_4_4_0_clk),
    .D(\tdc0.w_dly_sig[86] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[85] ));
 sky130_fd_sc_hd__dfxtp_1 _516_ (.CLK(clknet_4_4_0_clk),
    .D(\tdc0.w_dly_sig[87] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[86] ));
 sky130_fd_sc_hd__dfxtp_1 _517_ (.CLK(clknet_4_4_0_clk),
    .D(\tdc0.w_dly_sig[88] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[87] ));
 sky130_fd_sc_hd__dfxtp_1 _518_ (.CLK(clknet_4_5_0_clk),
    .D(\tdc0.w_dly_sig[89] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[88] ));
 sky130_fd_sc_hd__dfxtp_1 _519_ (.CLK(clknet_4_4_0_clk),
    .D(\tdc0.w_dly_sig[90] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[89] ));
 sky130_fd_sc_hd__dfxtp_1 _520_ (.CLK(clknet_4_4_0_clk),
    .D(\tdc0.w_dly_sig[91] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[90] ));
 sky130_fd_sc_hd__dfxtp_1 _521_ (.CLK(clknet_4_4_0_clk),
    .D(\tdc0.w_dly_sig[92] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[91] ));
 sky130_fd_sc_hd__dfxtp_1 _522_ (.CLK(clknet_4_6_0_clk),
    .D(\tdc0.w_dly_sig[93] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[92] ));
 sky130_fd_sc_hd__dfxtp_1 _523_ (.CLK(clknet_4_6_0_clk),
    .D(\tdc0.w_dly_sig[94] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[93] ));
 sky130_fd_sc_hd__dfxtp_1 _524_ (.CLK(clknet_4_6_0_clk),
    .D(\tdc0.w_dly_sig[95] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[94] ));
 sky130_fd_sc_hd__dfxtp_1 _525_ (.CLK(clknet_4_6_0_clk),
    .D(\tdc0.w_dly_sig[96] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[95] ));
 sky130_fd_sc_hd__dfxtp_1 _526_ (.CLK(clknet_4_6_0_clk),
    .D(\tdc0.w_dly_sig[97] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[96] ));
 sky130_fd_sc_hd__dfxtp_1 _527_ (.CLK(clknet_4_7_0_clk),
    .D(\tdc0.w_dly_sig[98] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[97] ));
 sky130_fd_sc_hd__dfxtp_1 _528_ (.CLK(clknet_4_7_0_clk),
    .D(\tdc0.w_dly_sig[99] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[98] ));
 sky130_fd_sc_hd__dfxtp_1 _529_ (.CLK(clknet_4_7_0_clk),
    .D(\tdc0.w_dly_sig[100] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[99] ));
 sky130_fd_sc_hd__dfxtp_1 _530_ (.CLK(clknet_4_5_0_clk),
    .D(\tdc0.w_dly_sig[101] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[100] ));
 sky130_fd_sc_hd__dfxtp_1 _531_ (.CLK(clknet_4_7_0_clk),
    .D(\tdc0.w_dly_sig[102] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[101] ));
 sky130_fd_sc_hd__dfxtp_1 _532_ (.CLK(clknet_4_5_0_clk),
    .D(\tdc0.w_dly_sig[103] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[102] ));
 sky130_fd_sc_hd__dfxtp_1 _533_ (.CLK(clknet_4_5_0_clk),
    .D(\tdc0.w_dly_sig[104] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[103] ));
 sky130_fd_sc_hd__dfxtp_1 _534_ (.CLK(clknet_4_7_0_clk),
    .D(\tdc0.w_dly_sig[105] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[104] ));
 sky130_fd_sc_hd__dfxtp_1 _535_ (.CLK(clknet_4_5_0_clk),
    .D(\tdc0.w_dly_sig[106] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[105] ));
 sky130_fd_sc_hd__dfxtp_1 _536_ (.CLK(clknet_4_5_0_clk),
    .D(\tdc0.w_dly_sig[107] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[106] ));
 sky130_fd_sc_hd__dfxtp_1 _537_ (.CLK(clknet_4_6_0_clk),
    .D(\tdc0.w_dly_sig[108] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[107] ));
 sky130_fd_sc_hd__dfxtp_1 _538_ (.CLK(clknet_4_5_0_clk),
    .D(\tdc0.w_dly_sig[109] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[108] ));
 sky130_fd_sc_hd__dfxtp_1 _539_ (.CLK(clknet_4_5_0_clk),
    .D(\tdc0.w_dly_sig[110] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[109] ));
 sky130_fd_sc_hd__dfxtp_1 _540_ (.CLK(clknet_4_5_0_clk),
    .D(\tdc0.w_dly_sig[111] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[110] ));
 sky130_fd_sc_hd__dfxtp_1 _541_ (.CLK(clknet_4_5_0_clk),
    .D(\tdc0.w_dly_sig[112] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[111] ));
 sky130_fd_sc_hd__dfxtp_1 _542_ (.CLK(clknet_4_5_0_clk),
    .D(\tdc0.w_dly_sig[113] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[112] ));
 sky130_fd_sc_hd__dfxtp_1 _543_ (.CLK(clknet_4_5_0_clk),
    .D(\tdc0.w_dly_sig[114] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[113] ));
 sky130_fd_sc_hd__dfxtp_1 _544_ (.CLK(clknet_4_5_0_clk),
    .D(\tdc0.w_dly_sig[115] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[114] ));
 sky130_fd_sc_hd__dfxtp_1 _545_ (.CLK(clknet_4_5_0_clk),
    .D(\tdc0.w_dly_sig[116] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[115] ));
 sky130_fd_sc_hd__dfxtp_1 _546_ (.CLK(clknet_4_5_0_clk),
    .D(\tdc0.w_dly_sig[117] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[116] ));
 sky130_fd_sc_hd__dfxtp_1 _547_ (.CLK(clknet_4_5_0_clk),
    .D(\tdc0.w_dly_sig[118] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[117] ));
 sky130_fd_sc_hd__dfxtp_1 _548_ (.CLK(clknet_4_5_0_clk),
    .D(\tdc0.w_dly_sig[119] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[118] ));
 sky130_fd_sc_hd__dfxtp_1 _549_ (.CLK(clknet_4_5_0_clk),
    .D(\tdc0.w_dly_sig[120] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[119] ));
 sky130_fd_sc_hd__dfxtp_1 _550_ (.CLK(clknet_4_5_0_clk),
    .D(\tdc0.w_dly_sig[121] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[120] ));
 sky130_fd_sc_hd__dfxtp_1 _551_ (.CLK(clknet_4_5_0_clk),
    .D(\tdc0.w_dly_sig[122] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[121] ));
 sky130_fd_sc_hd__dfxtp_1 _552_ (.CLK(clknet_4_4_0_clk),
    .D(\tdc0.w_dly_sig[123] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[122] ));
 sky130_fd_sc_hd__dfxtp_1 _553_ (.CLK(clknet_4_4_0_clk),
    .D(\tdc0.w_dly_sig[124] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[123] ));
 sky130_fd_sc_hd__dfxtp_1 _554_ (.CLK(clknet_4_4_0_clk),
    .D(\tdc0.w_dly_sig[125] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[124] ));
 sky130_fd_sc_hd__dfxtp_1 _555_ (.CLK(clknet_4_1_0_clk),
    .D(\tdc0.w_dly_sig[126] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[125] ));
 sky130_fd_sc_hd__dfxtp_1 _556_ (.CLK(clknet_4_1_0_clk),
    .D(\tdc0.w_dly_sig[127] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[126] ));
 sky130_fd_sc_hd__dfxtp_1 _557_ (.CLK(clknet_4_1_0_clk),
    .D(\tdc0.w_dly_sig[128] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[127] ));
 sky130_fd_sc_hd__dfxtp_1 _558_ (.CLK(clknet_4_4_0_clk),
    .D(\tdc0.w_dly_sig[129] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[128] ));
 sky130_fd_sc_hd__dfxtp_1 _559_ (.CLK(clknet_4_1_0_clk),
    .D(\tdc0.w_dly_sig[130] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[129] ));
 sky130_fd_sc_hd__dfxtp_1 _560_ (.CLK(clknet_4_0_0_clk),
    .D(\tdc0.w_dly_sig[131] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[130] ));
 sky130_fd_sc_hd__dfxtp_1 _561_ (.CLK(clknet_4_1_0_clk),
    .D(\tdc0.w_dly_sig[132] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[131] ));
 sky130_fd_sc_hd__dfxtp_1 _562_ (.CLK(clknet_4_0_0_clk),
    .D(\tdc0.w_dly_sig[133] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[132] ));
 sky130_fd_sc_hd__dfxtp_1 _563_ (.CLK(clknet_4_0_0_clk),
    .D(\tdc0.w_dly_sig[134] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[133] ));
 sky130_fd_sc_hd__dfxtp_1 _564_ (.CLK(clknet_4_0_0_clk),
    .D(\tdc0.w_dly_sig[135] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[134] ));
 sky130_fd_sc_hd__dfxtp_1 _565_ (.CLK(clknet_4_0_0_clk),
    .D(\tdc0.w_dly_sig[136] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[135] ));
 sky130_fd_sc_hd__dfxtp_1 _566_ (.CLK(clknet_4_2_0_clk),
    .D(\tdc0.w_dly_sig[137] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[136] ));
 sky130_fd_sc_hd__dfxtp_1 _567_ (.CLK(clknet_4_9_0_clk),
    .D(\tdc0.w_dly_sig[138] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[137] ));
 sky130_fd_sc_hd__dfxtp_1 _568_ (.CLK(clknet_4_2_0_clk),
    .D(\tdc0.w_dly_sig[139] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[138] ));
 sky130_fd_sc_hd__dfxtp_1 _569_ (.CLK(clknet_4_3_0_clk),
    .D(\tdc0.w_dly_sig[140] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[139] ));
 sky130_fd_sc_hd__dfxtp_1 _570_ (.CLK(clknet_4_3_0_clk),
    .D(\tdc0.w_dly_sig[141] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[140] ));
 sky130_fd_sc_hd__dfxtp_1 _571_ (.CLK(clknet_4_3_0_clk),
    .D(\tdc0.w_dly_sig[142] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[141] ));
 sky130_fd_sc_hd__dfxtp_1 _572_ (.CLK(clknet_4_9_0_clk),
    .D(\tdc0.w_dly_sig[143] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[142] ));
 sky130_fd_sc_hd__dfxtp_1 _573_ (.CLK(clknet_4_9_0_clk),
    .D(\tdc0.w_dly_sig[144] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[143] ));
 sky130_fd_sc_hd__dfxtp_1 _574_ (.CLK(clknet_4_9_0_clk),
    .D(\tdc0.w_dly_sig[145] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[144] ));
 sky130_fd_sc_hd__dfxtp_1 _575_ (.CLK(clknet_4_9_0_clk),
    .D(\tdc0.w_dly_sig[146] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[145] ));
 sky130_fd_sc_hd__dfxtp_1 _576_ (.CLK(clknet_4_9_0_clk),
    .D(\tdc0.w_dly_sig[147] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[146] ));
 sky130_fd_sc_hd__dfxtp_1 _577_ (.CLK(clknet_4_3_0_clk),
    .D(\tdc0.w_dly_sig[148] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[147] ));
 sky130_fd_sc_hd__dfxtp_1 _578_ (.CLK(clknet_4_9_0_clk),
    .D(\tdc0.w_dly_sig[149] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[148] ));
 sky130_fd_sc_hd__dfxtp_1 _579_ (.CLK(clknet_4_8_0_clk),
    .D(\tdc0.w_dly_sig[150] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[149] ));
 sky130_fd_sc_hd__dfxtp_1 _580_ (.CLK(clknet_4_0_0_clk),
    .D(\tdc0.w_dly_sig[151] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[150] ));
 sky130_fd_sc_hd__dfxtp_1 _581_ (.CLK(clknet_4_2_0_clk),
    .D(\tdc0.w_dly_sig[152] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[151] ));
 sky130_fd_sc_hd__dfxtp_1 _582_ (.CLK(clknet_4_2_0_clk),
    .D(\tdc0.w_dly_sig[153] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[152] ));
 sky130_fd_sc_hd__dfxtp_1 _583_ (.CLK(clknet_4_0_0_clk),
    .D(\tdc0.w_dly_sig[154] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[153] ));
 sky130_fd_sc_hd__dfxtp_1 _584_ (.CLK(clknet_4_0_0_clk),
    .D(\tdc0.w_dly_sig[155] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[154] ));
 sky130_fd_sc_hd__dfxtp_1 _585_ (.CLK(clknet_4_0_0_clk),
    .D(\tdc0.w_dly_sig[156] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[155] ));
 sky130_fd_sc_hd__dfxtp_1 _586_ (.CLK(clknet_4_2_0_clk),
    .D(\tdc0.w_dly_sig[157] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[156] ));
 sky130_fd_sc_hd__dfxtp_1 _587_ (.CLK(clknet_4_0_0_clk),
    .D(\tdc0.w_dly_sig[158] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[157] ));
 sky130_fd_sc_hd__dfxtp_1 _588_ (.CLK(clknet_4_9_0_clk),
    .D(\tdc0.w_dly_sig[159] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[158] ));
 sky130_fd_sc_hd__dfxtp_1 _589_ (.CLK(clknet_4_2_0_clk),
    .D(\tdc0.w_dly_sig[160] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[159] ));
 sky130_fd_sc_hd__dfxtp_1 _590_ (.CLK(clknet_4_2_0_clk),
    .D(\tdc0.w_dly_sig[161] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[160] ));
 sky130_fd_sc_hd__dfxtp_1 _591_ (.CLK(clknet_4_8_0_clk),
    .D(\tdc0.w_dly_sig[162] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[161] ));
 sky130_fd_sc_hd__dfxtp_1 _592_ (.CLK(clknet_4_2_0_clk),
    .D(\tdc0.w_dly_sig[163] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[162] ));
 sky130_fd_sc_hd__dfxtp_1 _593_ (.CLK(clknet_4_2_0_clk),
    .D(\tdc0.w_dly_sig[164] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[163] ));
 sky130_fd_sc_hd__dfxtp_1 _594_ (.CLK(clknet_4_8_0_clk),
    .D(\tdc0.w_dly_sig[165] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[164] ));
 sky130_fd_sc_hd__dfxtp_1 _595_ (.CLK(clknet_4_8_0_clk),
    .D(\tdc0.w_dly_sig[166] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[165] ));
 sky130_fd_sc_hd__dfxtp_1 _596_ (.CLK(clknet_4_2_0_clk),
    .D(\tdc0.w_dly_sig[167] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[166] ));
 sky130_fd_sc_hd__dfxtp_1 _597_ (.CLK(clknet_4_2_0_clk),
    .D(\tdc0.w_dly_sig[168] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[167] ));
 sky130_fd_sc_hd__dfxtp_1 _598_ (.CLK(clknet_4_2_0_clk),
    .D(\tdc0.w_dly_sig[169] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[168] ));
 sky130_fd_sc_hd__dfxtp_1 _599_ (.CLK(clknet_4_2_0_clk),
    .D(\tdc0.w_dly_sig[170] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[169] ));
 sky130_fd_sc_hd__dfxtp_1 _600_ (.CLK(clknet_4_8_0_clk),
    .D(\tdc0.w_dly_sig[171] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[170] ));
 sky130_fd_sc_hd__dfxtp_1 _601_ (.CLK(clknet_4_8_0_clk),
    .D(\tdc0.w_dly_sig[172] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[171] ));
 sky130_fd_sc_hd__dfxtp_1 _602_ (.CLK(clknet_4_8_0_clk),
    .D(\tdc0.w_dly_sig[173] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[172] ));
 sky130_fd_sc_hd__dfxtp_1 _603_ (.CLK(clknet_4_8_0_clk),
    .D(\tdc0.w_dly_sig[174] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[173] ));
 sky130_fd_sc_hd__dfxtp_1 _604_ (.CLK(clknet_4_8_0_clk),
    .D(\tdc0.w_dly_sig[175] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[174] ));
 sky130_fd_sc_hd__dfxtp_1 _605_ (.CLK(clknet_4_8_0_clk),
    .D(\tdc0.w_dly_sig[176] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[175] ));
 sky130_fd_sc_hd__dfxtp_1 _606_ (.CLK(clknet_4_8_0_clk),
    .D(\tdc0.w_dly_sig[177] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[176] ));
 sky130_fd_sc_hd__dfxtp_1 _607_ (.CLK(clknet_4_8_0_clk),
    .D(\tdc0.w_dly_sig[178] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[177] ));
 sky130_fd_sc_hd__dfxtp_1 _608_ (.CLK(clknet_4_8_0_clk),
    .D(\tdc0.w_dly_sig[179] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[178] ));
 sky130_fd_sc_hd__dfxtp_1 _609_ (.CLK(clknet_4_10_0_clk),
    .D(\tdc0.w_dly_sig[180] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[179] ));
 sky130_fd_sc_hd__dfxtp_1 _610_ (.CLK(clknet_4_10_0_clk),
    .D(\tdc0.w_dly_sig[181] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[180] ));
 sky130_fd_sc_hd__dfxtp_1 _611_ (.CLK(clknet_4_10_0_clk),
    .D(\tdc0.w_dly_sig[182] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[181] ));
 sky130_fd_sc_hd__dfxtp_1 _612_ (.CLK(clknet_4_10_0_clk),
    .D(\tdc0.w_dly_sig[183] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[182] ));
 sky130_fd_sc_hd__dfxtp_1 _613_ (.CLK(clknet_4_10_0_clk),
    .D(\tdc0.w_dly_sig[184] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[183] ));
 sky130_fd_sc_hd__dfxtp_1 _614_ (.CLK(clknet_4_10_0_clk),
    .D(\tdc0.w_dly_sig[185] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[184] ));
 sky130_fd_sc_hd__dfxtp_1 _615_ (.CLK(clknet_4_11_0_clk),
    .D(\tdc0.w_dly_sig[186] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[185] ));
 sky130_fd_sc_hd__dfxtp_1 _616_ (.CLK(clknet_4_10_0_clk),
    .D(\tdc0.w_dly_sig[187] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[186] ));
 sky130_fd_sc_hd__dfxtp_1 _617_ (.CLK(clknet_4_10_0_clk),
    .D(\tdc0.w_dly_sig[188] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[187] ));
 sky130_fd_sc_hd__dfxtp_1 _618_ (.CLK(clknet_4_11_0_clk),
    .D(\tdc0.w_dly_sig[189] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[188] ));
 sky130_fd_sc_hd__dfxtp_1 _619_ (.CLK(clknet_4_10_0_clk),
    .D(\tdc0.w_dly_sig[190] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[189] ));
 sky130_fd_sc_hd__dfxtp_1 _620_ (.CLK(clknet_4_10_0_clk),
    .D(\tdc0.w_dly_sig[191] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[190] ));
 sky130_fd_sc_hd__dfxtp_1 _621_ (.CLK(clknet_4_11_0_clk),
    .D(\tdc0.w_dly_sig[192] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tdc0.o_result[191] ));
 sky130_fd_sc_hd__buf_2 _638_ (.A(net1),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tdc0.w_dly_sig[0] ));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_4_0_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_4_10_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_4_11_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_4_12_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_4_13_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_4_14_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_4_15_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_4_1_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_4_2_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_4_3_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_4_4_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_4_5_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_4_6_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_4_7_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_4_8_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_4_9_0_clk));
 sky130_fd_sc_hd__buf_8 input1 (.A(ui_in[0]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net1));
 sky130_fd_sc_hd__buf_2 input2 (.A(ui_in[3]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net2));
 sky130_fd_sc_hd__buf_2 input3 (.A(ui_in[4]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_2 input4 (.A(ui_in[5]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net4));
 sky130_fd_sc_hd__buf_2 input5 (.A(ui_in[6]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_4 input6 (.A(ui_in[7]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net6));
 sky130_fd_sc_hd__buf_1 rebuffer1 (.A(\tdc0.w_dly_sig[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_1 rebuffer2 (.A(\tdc0.w_dly_sig[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_1 rebuffer3 (.A(\tdc0.w_dly_sig[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_1 rebuffer4 (.A(\tdc0.w_dly_sig[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_1 rebuffer5 (.A(\tdc0.w_dly_sig[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net27));
 sky130_fd_sc_hd__inv_4 \tdc0.g_dly_chain_even[0].dly_stg1  (.A(net1),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[0] ));
 sky130_fd_sc_hd__inv_4 \tdc0.g_dly_chain_even[0].dly_stg2  (.A(\tdc0.w_dly_sig_n[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[1] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[100].dly_stg1  (.A(\tdc0.w_dly_sig[100] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[100] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[100].dly_stg2  (.A(\tdc0.w_dly_sig_n[100] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[101] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[101].dly_stg1  (.A(\tdc0.w_dly_sig[101] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[101] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[101].dly_stg2  (.A(\tdc0.w_dly_sig_n[101] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[102] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[102].dly_stg1  (.A(\tdc0.w_dly_sig[102] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[102] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[102].dly_stg2  (.A(\tdc0.w_dly_sig_n[102] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[103] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[103].dly_stg1  (.A(\tdc0.w_dly_sig[103] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[103] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[103].dly_stg2  (.A(\tdc0.w_dly_sig_n[103] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[104] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[104].dly_stg1  (.A(\tdc0.w_dly_sig[104] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[104] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[104].dly_stg2  (.A(\tdc0.w_dly_sig_n[104] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[105] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[105].dly_stg1  (.A(\tdc0.w_dly_sig[105] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[105] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[105].dly_stg2  (.A(\tdc0.w_dly_sig_n[105] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[106] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[106].dly_stg1  (.A(\tdc0.w_dly_sig[106] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[106] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[106].dly_stg2  (.A(\tdc0.w_dly_sig_n[106] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[107] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[107].dly_stg1  (.A(\tdc0.w_dly_sig[107] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[107] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[107].dly_stg2  (.A(\tdc0.w_dly_sig_n[107] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[108] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[108].dly_stg1  (.A(\tdc0.w_dly_sig[108] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[108] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[108].dly_stg2  (.A(\tdc0.w_dly_sig_n[108] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[109] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[109].dly_stg1  (.A(\tdc0.w_dly_sig[109] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[109] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[109].dly_stg2  (.A(\tdc0.w_dly_sig_n[109] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[110] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[10].dly_stg1  (.A(\tdc0.w_dly_sig[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[10] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[10].dly_stg2  (.A(\tdc0.w_dly_sig_n[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[11] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[110].dly_stg1  (.A(\tdc0.w_dly_sig[110] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[110] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[110].dly_stg2  (.A(\tdc0.w_dly_sig_n[110] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[111] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[111].dly_stg1  (.A(\tdc0.w_dly_sig[111] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[111] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[111].dly_stg2  (.A(\tdc0.w_dly_sig_n[111] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[112] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[112].dly_stg1  (.A(\tdc0.w_dly_sig[112] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[112] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[112].dly_stg2  (.A(\tdc0.w_dly_sig_n[112] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[113] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[113].dly_stg1  (.A(\tdc0.w_dly_sig[113] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[113] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[113].dly_stg2  (.A(\tdc0.w_dly_sig_n[113] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[114] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[114].dly_stg1  (.A(\tdc0.w_dly_sig[114] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[114] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[114].dly_stg2  (.A(\tdc0.w_dly_sig_n[114] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[115] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[115].dly_stg1  (.A(\tdc0.w_dly_sig[115] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[115] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[115].dly_stg2  (.A(\tdc0.w_dly_sig_n[115] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[116] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[116].dly_stg1  (.A(\tdc0.w_dly_sig[116] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[116] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[116].dly_stg2  (.A(\tdc0.w_dly_sig_n[116] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[117] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[117].dly_stg1  (.A(\tdc0.w_dly_sig[117] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[117] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[117].dly_stg2  (.A(\tdc0.w_dly_sig_n[117] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[118] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[118].dly_stg1  (.A(\tdc0.w_dly_sig[118] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[118] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[118].dly_stg2  (.A(\tdc0.w_dly_sig_n[118] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[119] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[119].dly_stg1  (.A(\tdc0.w_dly_sig[119] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[119] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[119].dly_stg2  (.A(\tdc0.w_dly_sig_n[119] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[120] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[11].dly_stg1  (.A(\tdc0.w_dly_sig[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[11] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[11].dly_stg2  (.A(\tdc0.w_dly_sig_n[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[12] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[120].dly_stg1  (.A(\tdc0.w_dly_sig[120] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[120] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[120].dly_stg2  (.A(\tdc0.w_dly_sig_n[120] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[121] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[121].dly_stg1  (.A(\tdc0.w_dly_sig[121] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[121] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[121].dly_stg2  (.A(\tdc0.w_dly_sig_n[121] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[122] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[122].dly_stg1  (.A(\tdc0.w_dly_sig[122] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[122] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[122].dly_stg2  (.A(\tdc0.w_dly_sig_n[122] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[123] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[123].dly_stg1  (.A(\tdc0.w_dly_sig[123] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[123] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[123].dly_stg2  (.A(\tdc0.w_dly_sig_n[123] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[124] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[124].dly_stg1  (.A(\tdc0.w_dly_sig[124] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[124] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[124].dly_stg2  (.A(\tdc0.w_dly_sig_n[124] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[125] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[125].dly_stg1  (.A(\tdc0.w_dly_sig[125] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[125] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[125].dly_stg2  (.A(\tdc0.w_dly_sig_n[125] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[126] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[126].dly_stg1  (.A(\tdc0.w_dly_sig[126] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[126] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[126].dly_stg2  (.A(\tdc0.w_dly_sig_n[126] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[127] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[127].dly_stg1  (.A(\tdc0.w_dly_sig[127] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[127] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[127].dly_stg2  (.A(\tdc0.w_dly_sig_n[127] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[128] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[128].dly_stg1  (.A(\tdc0.w_dly_sig[128] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[128] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[128].dly_stg2  (.A(\tdc0.w_dly_sig_n[128] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[129] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[129].dly_stg1  (.A(\tdc0.w_dly_sig[129] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[129] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[129].dly_stg2  (.A(\tdc0.w_dly_sig_n[129] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[130] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[12].dly_stg1  (.A(\tdc0.w_dly_sig[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[12] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[12].dly_stg2  (.A(\tdc0.w_dly_sig_n[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[13] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[130].dly_stg1  (.A(\tdc0.w_dly_sig[130] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[130] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[130].dly_stg2  (.A(\tdc0.w_dly_sig_n[130] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[131] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[131].dly_stg1  (.A(\tdc0.w_dly_sig[131] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[131] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[131].dly_stg2  (.A(\tdc0.w_dly_sig_n[131] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[132] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[132].dly_stg1  (.A(\tdc0.w_dly_sig[132] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[132] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[132].dly_stg2  (.A(\tdc0.w_dly_sig_n[132] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[133] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[133].dly_stg1  (.A(\tdc0.w_dly_sig[133] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[133] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[133].dly_stg2  (.A(\tdc0.w_dly_sig_n[133] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[134] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[134].dly_stg1  (.A(\tdc0.w_dly_sig[134] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[134] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[134].dly_stg2  (.A(\tdc0.w_dly_sig_n[134] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[135] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[135].dly_stg1  (.A(\tdc0.w_dly_sig[135] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[135] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[135].dly_stg2  (.A(\tdc0.w_dly_sig_n[135] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[136] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[136].dly_stg1  (.A(\tdc0.w_dly_sig[136] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[136] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[136].dly_stg2  (.A(\tdc0.w_dly_sig_n[136] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[137] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[137].dly_stg1  (.A(\tdc0.w_dly_sig[137] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[137] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[137].dly_stg2  (.A(\tdc0.w_dly_sig_n[137] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[138] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[138].dly_stg1  (.A(\tdc0.w_dly_sig[138] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[138] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[138].dly_stg2  (.A(\tdc0.w_dly_sig_n[138] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[139] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[139].dly_stg1  (.A(\tdc0.w_dly_sig[139] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[139] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[139].dly_stg2  (.A(\tdc0.w_dly_sig_n[139] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[140] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[13].dly_stg1  (.A(\tdc0.w_dly_sig[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[13] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[13].dly_stg2  (.A(\tdc0.w_dly_sig_n[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[14] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[140].dly_stg1  (.A(\tdc0.w_dly_sig[140] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[140] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[140].dly_stg2  (.A(\tdc0.w_dly_sig_n[140] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[141] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[141].dly_stg1  (.A(\tdc0.w_dly_sig[141] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[141] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[141].dly_stg2  (.A(\tdc0.w_dly_sig_n[141] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[142] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[142].dly_stg1  (.A(\tdc0.w_dly_sig[142] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[142] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[142].dly_stg2  (.A(\tdc0.w_dly_sig_n[142] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[143] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[143].dly_stg1  (.A(\tdc0.w_dly_sig[143] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[143] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[143].dly_stg2  (.A(\tdc0.w_dly_sig_n[143] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[144] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[144].dly_stg1  (.A(\tdc0.w_dly_sig[144] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[144] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[144].dly_stg2  (.A(\tdc0.w_dly_sig_n[144] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[145] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[145].dly_stg1  (.A(\tdc0.w_dly_sig[145] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[145] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[145].dly_stg2  (.A(\tdc0.w_dly_sig_n[145] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[146] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[146].dly_stg1  (.A(\tdc0.w_dly_sig[146] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[146] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[146].dly_stg2  (.A(\tdc0.w_dly_sig_n[146] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[147] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[147].dly_stg1  (.A(\tdc0.w_dly_sig[147] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[147] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[147].dly_stg2  (.A(\tdc0.w_dly_sig_n[147] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[148] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[148].dly_stg1  (.A(\tdc0.w_dly_sig[148] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[148] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[148].dly_stg2  (.A(\tdc0.w_dly_sig_n[148] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[149] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[149].dly_stg1  (.A(\tdc0.w_dly_sig[149] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[149] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[149].dly_stg2  (.A(\tdc0.w_dly_sig_n[149] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[150] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[14].dly_stg1  (.A(\tdc0.w_dly_sig[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[14] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[14].dly_stg2  (.A(\tdc0.w_dly_sig_n[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[15] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[150].dly_stg1  (.A(\tdc0.w_dly_sig[150] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[150] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[150].dly_stg2  (.A(\tdc0.w_dly_sig_n[150] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[151] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[151].dly_stg1  (.A(\tdc0.w_dly_sig[151] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[151] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[151].dly_stg2  (.A(\tdc0.w_dly_sig_n[151] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[152] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[152].dly_stg1  (.A(\tdc0.w_dly_sig[152] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[152] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[152].dly_stg2  (.A(\tdc0.w_dly_sig_n[152] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[153] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[153].dly_stg1  (.A(\tdc0.w_dly_sig[153] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[153] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[153].dly_stg2  (.A(\tdc0.w_dly_sig_n[153] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[154] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[154].dly_stg1  (.A(\tdc0.w_dly_sig[154] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[154] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[154].dly_stg2  (.A(\tdc0.w_dly_sig_n[154] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[155] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[155].dly_stg1  (.A(\tdc0.w_dly_sig[155] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[155] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[155].dly_stg2  (.A(\tdc0.w_dly_sig_n[155] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[156] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[156].dly_stg1  (.A(\tdc0.w_dly_sig[156] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[156] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[156].dly_stg2  (.A(\tdc0.w_dly_sig_n[156] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[157] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[157].dly_stg1  (.A(\tdc0.w_dly_sig[157] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[157] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[157].dly_stg2  (.A(\tdc0.w_dly_sig_n[157] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[158] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[158].dly_stg1  (.A(\tdc0.w_dly_sig[158] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[158] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[158].dly_stg2  (.A(\tdc0.w_dly_sig_n[158] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[159] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[159].dly_stg1  (.A(\tdc0.w_dly_sig[159] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[159] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[159].dly_stg2  (.A(\tdc0.w_dly_sig_n[159] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[160] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[15].dly_stg1  (.A(\tdc0.w_dly_sig[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[15] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[15].dly_stg2  (.A(\tdc0.w_dly_sig_n[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[16] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[160].dly_stg1  (.A(\tdc0.w_dly_sig[160] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[160] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[160].dly_stg2  (.A(\tdc0.w_dly_sig_n[160] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[161] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[161].dly_stg1  (.A(\tdc0.w_dly_sig[161] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[161] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[161].dly_stg2  (.A(\tdc0.w_dly_sig_n[161] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[162] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[162].dly_stg1  (.A(\tdc0.w_dly_sig[162] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[162] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[162].dly_stg2  (.A(\tdc0.w_dly_sig_n[162] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[163] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[163].dly_stg1  (.A(\tdc0.w_dly_sig[163] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[163] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[163].dly_stg2  (.A(\tdc0.w_dly_sig_n[163] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[164] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[164].dly_stg1  (.A(\tdc0.w_dly_sig[164] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[164] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[164].dly_stg2  (.A(\tdc0.w_dly_sig_n[164] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[165] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[165].dly_stg1  (.A(\tdc0.w_dly_sig[165] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[165] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[165].dly_stg2  (.A(\tdc0.w_dly_sig_n[165] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[166] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[166].dly_stg1  (.A(\tdc0.w_dly_sig[166] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[166] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[166].dly_stg2  (.A(\tdc0.w_dly_sig_n[166] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[167] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[167].dly_stg1  (.A(\tdc0.w_dly_sig[167] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[167] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[167].dly_stg2  (.A(\tdc0.w_dly_sig_n[167] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[168] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[168].dly_stg1  (.A(\tdc0.w_dly_sig[168] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[168] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[168].dly_stg2  (.A(\tdc0.w_dly_sig_n[168] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[169] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[169].dly_stg1  (.A(\tdc0.w_dly_sig[169] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[169] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[169].dly_stg2  (.A(\tdc0.w_dly_sig_n[169] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[170] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[16].dly_stg1  (.A(\tdc0.w_dly_sig[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[16] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[16].dly_stg2  (.A(\tdc0.w_dly_sig_n[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[17] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[170].dly_stg1  (.A(\tdc0.w_dly_sig[170] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[170] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[170].dly_stg2  (.A(\tdc0.w_dly_sig_n[170] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[171] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[171].dly_stg1  (.A(\tdc0.w_dly_sig[171] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[171] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[171].dly_stg2  (.A(\tdc0.w_dly_sig_n[171] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[172] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[172].dly_stg1  (.A(\tdc0.w_dly_sig[172] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[172] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[172].dly_stg2  (.A(\tdc0.w_dly_sig_n[172] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[173] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[173].dly_stg1  (.A(\tdc0.w_dly_sig[173] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[173] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[173].dly_stg2  (.A(\tdc0.w_dly_sig_n[173] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[174] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[174].dly_stg1  (.A(\tdc0.w_dly_sig[174] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[174] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[174].dly_stg2  (.A(\tdc0.w_dly_sig_n[174] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[175] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[175].dly_stg1  (.A(\tdc0.w_dly_sig[175] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[175] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[175].dly_stg2  (.A(\tdc0.w_dly_sig_n[175] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[176] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[176].dly_stg1  (.A(\tdc0.w_dly_sig[176] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[176] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[176].dly_stg2  (.A(\tdc0.w_dly_sig_n[176] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[177] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[177].dly_stg1  (.A(\tdc0.w_dly_sig[177] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[177] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[177].dly_stg2  (.A(\tdc0.w_dly_sig_n[177] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[178] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[178].dly_stg1  (.A(\tdc0.w_dly_sig[178] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[178] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[178].dly_stg2  (.A(\tdc0.w_dly_sig_n[178] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[179] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[179].dly_stg1  (.A(\tdc0.w_dly_sig[179] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[179] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[179].dly_stg2  (.A(\tdc0.w_dly_sig_n[179] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[180] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[17].dly_stg1  (.A(\tdc0.w_dly_sig[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[17] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[17].dly_stg2  (.A(\tdc0.w_dly_sig_n[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[18] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[180].dly_stg1  (.A(\tdc0.w_dly_sig[180] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[180] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[180].dly_stg2  (.A(\tdc0.w_dly_sig_n[180] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[181] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[181].dly_stg1  (.A(\tdc0.w_dly_sig[181] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[181] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[181].dly_stg2  (.A(\tdc0.w_dly_sig_n[181] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[182] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[182].dly_stg1  (.A(\tdc0.w_dly_sig[182] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[182] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[182].dly_stg2  (.A(\tdc0.w_dly_sig_n[182] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[183] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[183].dly_stg1  (.A(\tdc0.w_dly_sig[183] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[183] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[183].dly_stg2  (.A(\tdc0.w_dly_sig_n[183] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[184] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[184].dly_stg1  (.A(\tdc0.w_dly_sig[184] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[184] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[184].dly_stg2  (.A(\tdc0.w_dly_sig_n[184] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[185] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[185].dly_stg1  (.A(\tdc0.w_dly_sig[185] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[185] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[185].dly_stg2  (.A(\tdc0.w_dly_sig_n[185] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[186] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[186].dly_stg1  (.A(\tdc0.w_dly_sig[186] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[186] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[186].dly_stg2  (.A(\tdc0.w_dly_sig_n[186] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[187] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[187].dly_stg1  (.A(\tdc0.w_dly_sig[187] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[187] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[187].dly_stg2  (.A(\tdc0.w_dly_sig_n[187] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[188] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[188].dly_stg1  (.A(\tdc0.w_dly_sig[188] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[188] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[188].dly_stg2  (.A(\tdc0.w_dly_sig_n[188] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[189] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[189].dly_stg1  (.A(\tdc0.w_dly_sig[189] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[189] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[189].dly_stg2  (.A(\tdc0.w_dly_sig_n[189] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[190] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[18].dly_stg1  (.A(\tdc0.w_dly_sig[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[18] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[18].dly_stg2  (.A(\tdc0.w_dly_sig_n[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[19] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[190].dly_stg1  (.A(\tdc0.w_dly_sig[190] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[190] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[190].dly_stg2  (.A(\tdc0.w_dly_sig_n[190] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[191] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[191].dly_stg1  (.A(\tdc0.w_dly_sig[191] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[191] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[191].dly_stg2  (.A(\tdc0.w_dly_sig_n[191] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[192] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[192].dly_stg1  (.A(\tdc0.w_dly_sig[192] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[192] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[192].dly_stg2  (.A(\tdc0.w_dly_sig_n[192] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[193] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[19].dly_stg1  (.A(\tdc0.w_dly_sig[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[19] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[19].dly_stg2  (.A(\tdc0.w_dly_sig_n[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[20] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[1].dly_stg1  (.A(\tdc0.w_dly_sig[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[1] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[1].dly_stg2  (.A(\tdc0.w_dly_sig_n[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[2] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[20].dly_stg1  (.A(\tdc0.w_dly_sig[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[20] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[20].dly_stg2  (.A(\tdc0.w_dly_sig_n[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[21] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[21].dly_stg1  (.A(\tdc0.w_dly_sig[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[21] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[21].dly_stg2  (.A(\tdc0.w_dly_sig_n[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[22] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[22].dly_stg1  (.A(\tdc0.w_dly_sig[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[22] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[22].dly_stg2  (.A(\tdc0.w_dly_sig_n[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[23] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[23].dly_stg1  (.A(\tdc0.w_dly_sig[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[23] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[23].dly_stg2  (.A(\tdc0.w_dly_sig_n[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[24] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[24].dly_stg1  (.A(\tdc0.w_dly_sig[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[24] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[24].dly_stg2  (.A(\tdc0.w_dly_sig_n[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[25] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[25].dly_stg1  (.A(\tdc0.w_dly_sig[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[25] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[25].dly_stg2  (.A(\tdc0.w_dly_sig_n[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[26] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[26].dly_stg1  (.A(\tdc0.w_dly_sig[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[26] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[26].dly_stg2  (.A(\tdc0.w_dly_sig_n[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[27] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[27].dly_stg1  (.A(\tdc0.w_dly_sig[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[27] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[27].dly_stg2  (.A(\tdc0.w_dly_sig_n[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[28] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[28].dly_stg1  (.A(\tdc0.w_dly_sig[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[28] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[28].dly_stg2  (.A(\tdc0.w_dly_sig_n[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[29] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[29].dly_stg1  (.A(\tdc0.w_dly_sig[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[29] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[29].dly_stg2  (.A(\tdc0.w_dly_sig_n[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[30] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[2].dly_stg1  (.A(\tdc0.w_dly_sig[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[2] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[2].dly_stg2  (.A(\tdc0.w_dly_sig_n[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[3] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[30].dly_stg1  (.A(\tdc0.w_dly_sig[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[30] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[30].dly_stg2  (.A(\tdc0.w_dly_sig_n[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[31] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[31].dly_stg1  (.A(\tdc0.w_dly_sig[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[31] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[31].dly_stg2  (.A(\tdc0.w_dly_sig_n[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[32] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[32].dly_stg1  (.A(\tdc0.w_dly_sig[32] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[32] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[32].dly_stg2  (.A(\tdc0.w_dly_sig_n[32] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[33] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[33].dly_stg1  (.A(\tdc0.w_dly_sig[33] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[33] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[33].dly_stg2  (.A(\tdc0.w_dly_sig_n[33] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[34] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[34].dly_stg1  (.A(\tdc0.w_dly_sig[34] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[34] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[34].dly_stg2  (.A(\tdc0.w_dly_sig_n[34] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[35] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[35].dly_stg1  (.A(\tdc0.w_dly_sig[35] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[35] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[35].dly_stg2  (.A(\tdc0.w_dly_sig_n[35] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[36] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[36].dly_stg1  (.A(\tdc0.w_dly_sig[36] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[36] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[36].dly_stg2  (.A(\tdc0.w_dly_sig_n[36] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[37] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[37].dly_stg1  (.A(\tdc0.w_dly_sig[37] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[37] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[37].dly_stg2  (.A(\tdc0.w_dly_sig_n[37] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[38] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[38].dly_stg1  (.A(\tdc0.w_dly_sig[38] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[38] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[38].dly_stg2  (.A(\tdc0.w_dly_sig_n[38] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[39] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[39].dly_stg1  (.A(\tdc0.w_dly_sig[39] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[39] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[39].dly_stg2  (.A(\tdc0.w_dly_sig_n[39] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[40] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[3].dly_stg1  (.A(\tdc0.w_dly_sig[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[3] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[3].dly_stg2  (.A(\tdc0.w_dly_sig_n[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[4] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[40].dly_stg1  (.A(\tdc0.w_dly_sig[40] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[40] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[40].dly_stg2  (.A(\tdc0.w_dly_sig_n[40] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[41] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[41].dly_stg1  (.A(\tdc0.w_dly_sig[41] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[41] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[41].dly_stg2  (.A(\tdc0.w_dly_sig_n[41] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[42] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[42].dly_stg1  (.A(\tdc0.w_dly_sig[42] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[42] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[42].dly_stg2  (.A(\tdc0.w_dly_sig_n[42] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[43] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[43].dly_stg1  (.A(\tdc0.w_dly_sig[43] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[43] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[43].dly_stg2  (.A(\tdc0.w_dly_sig_n[43] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[44] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[44].dly_stg1  (.A(\tdc0.w_dly_sig[44] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[44] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[44].dly_stg2  (.A(\tdc0.w_dly_sig_n[44] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[45] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[45].dly_stg1  (.A(\tdc0.w_dly_sig[45] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[45] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[45].dly_stg2  (.A(\tdc0.w_dly_sig_n[45] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[46] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[46].dly_stg1  (.A(\tdc0.w_dly_sig[46] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[46] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[46].dly_stg2  (.A(\tdc0.w_dly_sig_n[46] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[47] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[47].dly_stg1  (.A(\tdc0.w_dly_sig[47] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[47] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[47].dly_stg2  (.A(\tdc0.w_dly_sig_n[47] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[48] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[48].dly_stg1  (.A(\tdc0.w_dly_sig[48] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[48] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[48].dly_stg2  (.A(\tdc0.w_dly_sig_n[48] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[49] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[49].dly_stg1  (.A(\tdc0.w_dly_sig[49] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[49] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[49].dly_stg2  (.A(\tdc0.w_dly_sig_n[49] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[50] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[4].dly_stg1  (.A(\tdc0.w_dly_sig[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[4] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[4].dly_stg2  (.A(\tdc0.w_dly_sig_n[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[5] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[50].dly_stg1  (.A(\tdc0.w_dly_sig[50] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[50] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[50].dly_stg2  (.A(\tdc0.w_dly_sig_n[50] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[51] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[51].dly_stg1  (.A(\tdc0.w_dly_sig[51] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[51] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[51].dly_stg2  (.A(\tdc0.w_dly_sig_n[51] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[52] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[52].dly_stg1  (.A(\tdc0.w_dly_sig[52] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[52] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[52].dly_stg2  (.A(\tdc0.w_dly_sig_n[52] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[53] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[53].dly_stg1  (.A(\tdc0.w_dly_sig[53] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[53] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[53].dly_stg2  (.A(\tdc0.w_dly_sig_n[53] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[54] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[54].dly_stg1  (.A(\tdc0.w_dly_sig[54] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[54] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[54].dly_stg2  (.A(\tdc0.w_dly_sig_n[54] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[55] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[55].dly_stg1  (.A(\tdc0.w_dly_sig[55] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[55] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[55].dly_stg2  (.A(\tdc0.w_dly_sig_n[55] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[56] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[56].dly_stg1  (.A(\tdc0.w_dly_sig[56] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[56] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[56].dly_stg2  (.A(\tdc0.w_dly_sig_n[56] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[57] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[57].dly_stg1  (.A(\tdc0.w_dly_sig[57] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[57] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[57].dly_stg2  (.A(\tdc0.w_dly_sig_n[57] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[58] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[58].dly_stg1  (.A(\tdc0.w_dly_sig[58] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[58] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[58].dly_stg2  (.A(\tdc0.w_dly_sig_n[58] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[59] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[59].dly_stg1  (.A(\tdc0.w_dly_sig[59] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[59] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[59].dly_stg2  (.A(\tdc0.w_dly_sig_n[59] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[60] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[5].dly_stg1  (.A(\tdc0.w_dly_sig[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[5] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[5].dly_stg2  (.A(\tdc0.w_dly_sig_n[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[6] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[60].dly_stg1  (.A(\tdc0.w_dly_sig[60] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[60] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[60].dly_stg2  (.A(\tdc0.w_dly_sig_n[60] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[61] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[61].dly_stg1  (.A(\tdc0.w_dly_sig[61] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[61] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[61].dly_stg2  (.A(\tdc0.w_dly_sig_n[61] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[62] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[62].dly_stg1  (.A(\tdc0.w_dly_sig[62] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[62] ));
 sky130_fd_sc_hd__inv_4 \tdc0.g_dly_chain_even[62].dly_stg2  (.A(\tdc0.w_dly_sig_n[62] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[63] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[63].dly_stg1  (.A(\tdc0.w_dly_sig[63] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[63] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[63].dly_stg2  (.A(\tdc0.w_dly_sig_n[63] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[64] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[64].dly_stg1  (.A(\tdc0.w_dly_sig[64] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[64] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[64].dly_stg2  (.A(\tdc0.w_dly_sig_n[64] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[65] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[65].dly_stg1  (.A(\tdc0.w_dly_sig[65] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[65] ));
 sky130_fd_sc_hd__inv_4 \tdc0.g_dly_chain_even[65].dly_stg2  (.A(\tdc0.w_dly_sig_n[65] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[66] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[66].dly_stg1  (.A(\tdc0.w_dly_sig[66] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[66] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[66].dly_stg2  (.A(\tdc0.w_dly_sig_n[66] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[67] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[67].dly_stg1  (.A(\tdc0.w_dly_sig[67] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[67] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[67].dly_stg2  (.A(\tdc0.w_dly_sig_n[67] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[68] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[68].dly_stg1  (.A(\tdc0.w_dly_sig[68] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[68] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[68].dly_stg2  (.A(\tdc0.w_dly_sig_n[68] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[69] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[69].dly_stg1  (.A(\tdc0.w_dly_sig[69] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[69] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[69].dly_stg2  (.A(\tdc0.w_dly_sig_n[69] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[70] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[6].dly_stg1  (.A(\tdc0.w_dly_sig[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[6] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[6].dly_stg2  (.A(\tdc0.w_dly_sig_n[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[7] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[70].dly_stg1  (.A(\tdc0.w_dly_sig[70] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[70] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[70].dly_stg2  (.A(\tdc0.w_dly_sig_n[70] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[71] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[71].dly_stg1  (.A(\tdc0.w_dly_sig[71] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[71] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[71].dly_stg2  (.A(\tdc0.w_dly_sig_n[71] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[72] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[72].dly_stg1  (.A(\tdc0.w_dly_sig[72] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[72] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[72].dly_stg2  (.A(\tdc0.w_dly_sig_n[72] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[73] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[73].dly_stg1  (.A(\tdc0.w_dly_sig[73] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[73] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[73].dly_stg2  (.A(\tdc0.w_dly_sig_n[73] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[74] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[74].dly_stg1  (.A(\tdc0.w_dly_sig[74] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[74] ));
 sky130_fd_sc_hd__inv_4 \tdc0.g_dly_chain_even[74].dly_stg2  (.A(\tdc0.w_dly_sig_n[74] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[75] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[75].dly_stg1  (.A(\tdc0.w_dly_sig[75] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[75] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[75].dly_stg2  (.A(\tdc0.w_dly_sig_n[75] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[76] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[76].dly_stg1  (.A(\tdc0.w_dly_sig[76] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[76] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[76].dly_stg2  (.A(\tdc0.w_dly_sig_n[76] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[77] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[77].dly_stg1  (.A(\tdc0.w_dly_sig[77] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[77] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[77].dly_stg2  (.A(\tdc0.w_dly_sig_n[77] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[78] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[78].dly_stg1  (.A(\tdc0.w_dly_sig[78] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[78] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[78].dly_stg2  (.A(\tdc0.w_dly_sig_n[78] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[79] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[79].dly_stg1  (.A(\tdc0.w_dly_sig[79] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[79] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[79].dly_stg2  (.A(\tdc0.w_dly_sig_n[79] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[80] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[7].dly_stg1  (.A(\tdc0.w_dly_sig[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[7] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[7].dly_stg2  (.A(\tdc0.w_dly_sig_n[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[8] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[80].dly_stg1  (.A(\tdc0.w_dly_sig[80] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[80] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[80].dly_stg2  (.A(\tdc0.w_dly_sig_n[80] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[81] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[81].dly_stg1  (.A(\tdc0.w_dly_sig[81] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[81] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[81].dly_stg2  (.A(\tdc0.w_dly_sig_n[81] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[82] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[82].dly_stg1  (.A(\tdc0.w_dly_sig[82] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[82] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[82].dly_stg2  (.A(\tdc0.w_dly_sig_n[82] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[83] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[83].dly_stg1  (.A(\tdc0.w_dly_sig[83] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[83] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[83].dly_stg2  (.A(\tdc0.w_dly_sig_n[83] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[84] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[84].dly_stg1  (.A(\tdc0.w_dly_sig[84] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[84] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[84].dly_stg2  (.A(\tdc0.w_dly_sig_n[84] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[85] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[85].dly_stg1  (.A(\tdc0.w_dly_sig[85] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[85] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[85].dly_stg2  (.A(\tdc0.w_dly_sig_n[85] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[86] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[86].dly_stg1  (.A(\tdc0.w_dly_sig[86] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[86] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[86].dly_stg2  (.A(\tdc0.w_dly_sig_n[86] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[87] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[87].dly_stg1  (.A(\tdc0.w_dly_sig[87] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[87] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[87].dly_stg2  (.A(\tdc0.w_dly_sig_n[87] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[88] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[88].dly_stg1  (.A(\tdc0.w_dly_sig[88] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[88] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[88].dly_stg2  (.A(\tdc0.w_dly_sig_n[88] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[89] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[89].dly_stg1  (.A(\tdc0.w_dly_sig[89] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[89] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[89].dly_stg2  (.A(\tdc0.w_dly_sig_n[89] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[90] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[8].dly_stg1  (.A(\tdc0.w_dly_sig[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[8] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[8].dly_stg2  (.A(\tdc0.w_dly_sig_n[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[9] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[90].dly_stg1  (.A(\tdc0.w_dly_sig[90] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[90] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[90].dly_stg2  (.A(\tdc0.w_dly_sig_n[90] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[91] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[91].dly_stg1  (.A(\tdc0.w_dly_sig[91] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[91] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[91].dly_stg2  (.A(\tdc0.w_dly_sig_n[91] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[92] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[92].dly_stg1  (.A(\tdc0.w_dly_sig[92] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[92] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[92].dly_stg2  (.A(\tdc0.w_dly_sig_n[92] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[93] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[93].dly_stg1  (.A(\tdc0.w_dly_sig[93] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[93] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[93].dly_stg2  (.A(\tdc0.w_dly_sig_n[93] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[94] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[94].dly_stg1  (.A(\tdc0.w_dly_sig[94] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[94] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[94].dly_stg2  (.A(\tdc0.w_dly_sig_n[94] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[95] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[95].dly_stg1  (.A(\tdc0.w_dly_sig[95] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[95] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[95].dly_stg2  (.A(\tdc0.w_dly_sig_n[95] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[96] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[96].dly_stg1  (.A(\tdc0.w_dly_sig[96] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[96] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[96].dly_stg2  (.A(\tdc0.w_dly_sig_n[96] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[97] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[97].dly_stg1  (.A(\tdc0.w_dly_sig[97] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[97] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[97].dly_stg2  (.A(\tdc0.w_dly_sig_n[97] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[98] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[98].dly_stg1  (.A(\tdc0.w_dly_sig[98] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[98] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[98].dly_stg2  (.A(\tdc0.w_dly_sig_n[98] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[99] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[99].dly_stg1  (.A(\tdc0.w_dly_sig[99] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[99] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[99].dly_stg2  (.A(\tdc0.w_dly_sig_n[99] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[100] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[9].dly_stg1  (.A(\tdc0.w_dly_sig[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[9] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_even[9].dly_stg2  (.A(\tdc0.w_dly_sig_n[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[10] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[0].dly_stg1  (.A(net1),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[1] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[0].dly_stg2  (.A(\tdc0.w_dly_sig_n[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[2] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[100].dly_stg1  (.A(\tdc0.w_dly_sig[100] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[101] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[100].dly_stg2  (.A(\tdc0.w_dly_sig_n[100] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[102] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[101].dly_stg1  (.A(\tdc0.w_dly_sig[101] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[102] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[101].dly_stg2  (.A(\tdc0.w_dly_sig_n[101] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[103] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[102].dly_stg1  (.A(\tdc0.w_dly_sig[102] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[103] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[102].dly_stg2  (.A(\tdc0.w_dly_sig_n[102] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[104] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[103].dly_stg1  (.A(\tdc0.w_dly_sig[103] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[104] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[103].dly_stg2  (.A(\tdc0.w_dly_sig_n[103] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[105] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[104].dly_stg1  (.A(\tdc0.w_dly_sig[104] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[105] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[104].dly_stg2  (.A(\tdc0.w_dly_sig_n[104] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[106] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[105].dly_stg1  (.A(\tdc0.w_dly_sig[105] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[106] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[105].dly_stg2  (.A(\tdc0.w_dly_sig_n[105] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[107] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[106].dly_stg1  (.A(\tdc0.w_dly_sig[106] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[107] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[106].dly_stg2  (.A(\tdc0.w_dly_sig_n[106] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[108] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[107].dly_stg1  (.A(\tdc0.w_dly_sig[107] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[108] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[107].dly_stg2  (.A(\tdc0.w_dly_sig_n[107] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[109] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[108].dly_stg1  (.A(\tdc0.w_dly_sig[108] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[109] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[108].dly_stg2  (.A(\tdc0.w_dly_sig_n[108] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[110] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[109].dly_stg1  (.A(\tdc0.w_dly_sig[109] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[110] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[109].dly_stg2  (.A(\tdc0.w_dly_sig_n[109] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[111] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[10].dly_stg1  (.A(\tdc0.w_dly_sig[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[11] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[10].dly_stg2  (.A(\tdc0.w_dly_sig_n[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[12] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[110].dly_stg1  (.A(\tdc0.w_dly_sig[110] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[111] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[110].dly_stg2  (.A(\tdc0.w_dly_sig_n[110] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[112] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[111].dly_stg1  (.A(\tdc0.w_dly_sig[111] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[112] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[111].dly_stg2  (.A(\tdc0.w_dly_sig_n[111] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[113] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[112].dly_stg1  (.A(\tdc0.w_dly_sig[112] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[113] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[112].dly_stg2  (.A(\tdc0.w_dly_sig_n[112] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[114] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[113].dly_stg1  (.A(\tdc0.w_dly_sig[113] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[114] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[113].dly_stg2  (.A(\tdc0.w_dly_sig_n[113] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[115] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[114].dly_stg1  (.A(\tdc0.w_dly_sig[114] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[115] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[114].dly_stg2  (.A(\tdc0.w_dly_sig_n[114] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[116] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[115].dly_stg1  (.A(\tdc0.w_dly_sig[115] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[116] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[115].dly_stg2  (.A(\tdc0.w_dly_sig_n[115] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[117] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[116].dly_stg1  (.A(\tdc0.w_dly_sig[116] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[117] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[116].dly_stg2  (.A(\tdc0.w_dly_sig_n[116] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[118] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[117].dly_stg1  (.A(\tdc0.w_dly_sig[117] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[118] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[117].dly_stg2  (.A(\tdc0.w_dly_sig_n[117] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[119] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[118].dly_stg1  (.A(\tdc0.w_dly_sig[118] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[119] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[118].dly_stg2  (.A(\tdc0.w_dly_sig_n[118] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[120] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[119].dly_stg1  (.A(\tdc0.w_dly_sig[119] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[120] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[119].dly_stg2  (.A(\tdc0.w_dly_sig_n[119] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[121] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[11].dly_stg1  (.A(\tdc0.w_dly_sig[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[12] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[11].dly_stg2  (.A(\tdc0.w_dly_sig_n[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[13] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[120].dly_stg1  (.A(\tdc0.w_dly_sig[120] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[121] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[120].dly_stg2  (.A(\tdc0.w_dly_sig_n[120] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[122] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[121].dly_stg1  (.A(\tdc0.w_dly_sig[121] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[122] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[121].dly_stg2  (.A(\tdc0.w_dly_sig_n[121] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[123] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[122].dly_stg1  (.A(\tdc0.w_dly_sig[122] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[123] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[122].dly_stg2  (.A(\tdc0.w_dly_sig_n[122] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[124] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[123].dly_stg1  (.A(\tdc0.w_dly_sig[123] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[124] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[123].dly_stg2  (.A(\tdc0.w_dly_sig_n[123] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[125] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[124].dly_stg1  (.A(\tdc0.w_dly_sig[124] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[125] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[124].dly_stg2  (.A(\tdc0.w_dly_sig_n[124] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[126] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[125].dly_stg1  (.A(\tdc0.w_dly_sig[125] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[126] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[125].dly_stg2  (.A(\tdc0.w_dly_sig_n[125] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[127] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[126].dly_stg1  (.A(\tdc0.w_dly_sig[126] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[127] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[126].dly_stg2  (.A(\tdc0.w_dly_sig_n[126] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[128] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[127].dly_stg1  (.A(\tdc0.w_dly_sig[127] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[128] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[127].dly_stg2  (.A(\tdc0.w_dly_sig_n[127] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[129] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[128].dly_stg1  (.A(\tdc0.w_dly_sig[128] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[129] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[128].dly_stg2  (.A(\tdc0.w_dly_sig_n[128] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[130] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[129].dly_stg1  (.A(\tdc0.w_dly_sig[129] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[130] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[129].dly_stg2  (.A(\tdc0.w_dly_sig_n[129] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[131] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[12].dly_stg1  (.A(\tdc0.w_dly_sig[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[13] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[12].dly_stg2  (.A(\tdc0.w_dly_sig_n[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[14] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[130].dly_stg1  (.A(\tdc0.w_dly_sig[130] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[131] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[130].dly_stg2  (.A(\tdc0.w_dly_sig_n[130] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[132] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[131].dly_stg1  (.A(\tdc0.w_dly_sig[131] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[132] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[131].dly_stg2  (.A(\tdc0.w_dly_sig_n[131] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[133] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[132].dly_stg1  (.A(\tdc0.w_dly_sig[132] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[133] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[132].dly_stg2  (.A(\tdc0.w_dly_sig_n[132] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[134] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[133].dly_stg1  (.A(\tdc0.w_dly_sig[133] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[134] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[133].dly_stg2  (.A(\tdc0.w_dly_sig_n[133] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[135] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[134].dly_stg1  (.A(\tdc0.w_dly_sig[134] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[135] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[134].dly_stg2  (.A(\tdc0.w_dly_sig_n[134] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[136] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[135].dly_stg1  (.A(\tdc0.w_dly_sig[135] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[136] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[135].dly_stg2  (.A(\tdc0.w_dly_sig_n[135] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[137] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[136].dly_stg1  (.A(\tdc0.w_dly_sig[136] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[137] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[136].dly_stg2  (.A(\tdc0.w_dly_sig_n[136] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[138] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[137].dly_stg1  (.A(\tdc0.w_dly_sig[137] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[138] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[137].dly_stg2  (.A(\tdc0.w_dly_sig_n[137] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[139] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[138].dly_stg1  (.A(\tdc0.w_dly_sig[138] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[139] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[138].dly_stg2  (.A(\tdc0.w_dly_sig_n[138] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[140] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[139].dly_stg1  (.A(\tdc0.w_dly_sig[139] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[140] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[139].dly_stg2  (.A(\tdc0.w_dly_sig_n[139] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[141] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[13].dly_stg1  (.A(\tdc0.w_dly_sig[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[14] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[13].dly_stg2  (.A(\tdc0.w_dly_sig_n[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[15] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[140].dly_stg1  (.A(\tdc0.w_dly_sig[140] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[141] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[140].dly_stg2  (.A(\tdc0.w_dly_sig_n[140] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[142] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[141].dly_stg1  (.A(\tdc0.w_dly_sig[141] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[142] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[141].dly_stg2  (.A(\tdc0.w_dly_sig_n[141] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[143] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[142].dly_stg1  (.A(\tdc0.w_dly_sig[142] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[143] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[142].dly_stg2  (.A(\tdc0.w_dly_sig_n[142] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[144] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[143].dly_stg1  (.A(\tdc0.w_dly_sig[143] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[144] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[143].dly_stg2  (.A(\tdc0.w_dly_sig_n[143] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[145] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[144].dly_stg1  (.A(\tdc0.w_dly_sig[144] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[145] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[144].dly_stg2  (.A(\tdc0.w_dly_sig_n[144] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[146] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[145].dly_stg1  (.A(\tdc0.w_dly_sig[145] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[146] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[145].dly_stg2  (.A(\tdc0.w_dly_sig_n[145] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[147] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[146].dly_stg1  (.A(\tdc0.w_dly_sig[146] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[147] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[146].dly_stg2  (.A(\tdc0.w_dly_sig_n[146] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[148] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[147].dly_stg1  (.A(\tdc0.w_dly_sig[147] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[148] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[147].dly_stg2  (.A(\tdc0.w_dly_sig_n[147] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[149] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[148].dly_stg1  (.A(\tdc0.w_dly_sig[148] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[149] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[148].dly_stg2  (.A(\tdc0.w_dly_sig_n[148] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[150] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[149].dly_stg1  (.A(\tdc0.w_dly_sig[149] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[150] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[149].dly_stg2  (.A(\tdc0.w_dly_sig_n[149] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[151] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[14].dly_stg1  (.A(\tdc0.w_dly_sig[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[15] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[14].dly_stg2  (.A(\tdc0.w_dly_sig_n[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[16] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[150].dly_stg1  (.A(\tdc0.w_dly_sig[150] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[151] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[150].dly_stg2  (.A(\tdc0.w_dly_sig_n[150] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[152] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[151].dly_stg1  (.A(\tdc0.w_dly_sig[151] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[152] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[151].dly_stg2  (.A(\tdc0.w_dly_sig_n[151] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[153] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[152].dly_stg1  (.A(\tdc0.w_dly_sig[152] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[153] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[152].dly_stg2  (.A(\tdc0.w_dly_sig_n[152] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[154] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[153].dly_stg1  (.A(\tdc0.w_dly_sig[153] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[154] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[153].dly_stg2  (.A(\tdc0.w_dly_sig_n[153] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[155] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[154].dly_stg1  (.A(\tdc0.w_dly_sig[154] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[155] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[154].dly_stg2  (.A(\tdc0.w_dly_sig_n[154] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[156] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[155].dly_stg1  (.A(\tdc0.w_dly_sig[155] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[156] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[155].dly_stg2  (.A(\tdc0.w_dly_sig_n[155] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[157] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[156].dly_stg1  (.A(\tdc0.w_dly_sig[156] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[157] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[156].dly_stg2  (.A(\tdc0.w_dly_sig_n[156] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[158] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[157].dly_stg1  (.A(\tdc0.w_dly_sig[157] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[158] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[157].dly_stg2  (.A(\tdc0.w_dly_sig_n[157] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[159] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[158].dly_stg1  (.A(\tdc0.w_dly_sig[158] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[159] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[158].dly_stg2  (.A(\tdc0.w_dly_sig_n[158] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[160] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[159].dly_stg1  (.A(\tdc0.w_dly_sig[159] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[160] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[159].dly_stg2  (.A(\tdc0.w_dly_sig_n[159] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[161] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[15].dly_stg1  (.A(\tdc0.w_dly_sig[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[16] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[15].dly_stg2  (.A(\tdc0.w_dly_sig_n[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[17] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[160].dly_stg1  (.A(\tdc0.w_dly_sig[160] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[161] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[160].dly_stg2  (.A(\tdc0.w_dly_sig_n[160] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[162] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[161].dly_stg1  (.A(\tdc0.w_dly_sig[161] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[162] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[161].dly_stg2  (.A(\tdc0.w_dly_sig_n[161] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[163] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[162].dly_stg1  (.A(\tdc0.w_dly_sig[162] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[163] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[162].dly_stg2  (.A(\tdc0.w_dly_sig_n[162] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[164] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[163].dly_stg1  (.A(\tdc0.w_dly_sig[163] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[164] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[163].dly_stg2  (.A(\tdc0.w_dly_sig_n[163] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[165] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[164].dly_stg1  (.A(\tdc0.w_dly_sig[164] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[165] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[164].dly_stg2  (.A(\tdc0.w_dly_sig_n[164] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[166] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[165].dly_stg1  (.A(\tdc0.w_dly_sig[165] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[166] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[165].dly_stg2  (.A(\tdc0.w_dly_sig_n[165] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[167] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[166].dly_stg1  (.A(\tdc0.w_dly_sig[166] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[167] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[166].dly_stg2  (.A(\tdc0.w_dly_sig_n[166] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[168] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[167].dly_stg1  (.A(\tdc0.w_dly_sig[167] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[168] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[167].dly_stg2  (.A(\tdc0.w_dly_sig_n[167] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[169] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[168].dly_stg1  (.A(\tdc0.w_dly_sig[168] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[169] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[168].dly_stg2  (.A(\tdc0.w_dly_sig_n[168] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[170] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[169].dly_stg1  (.A(\tdc0.w_dly_sig[169] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[170] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[169].dly_stg2  (.A(\tdc0.w_dly_sig_n[169] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[171] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[16].dly_stg1  (.A(\tdc0.w_dly_sig[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[17] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[16].dly_stg2  (.A(\tdc0.w_dly_sig_n[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[18] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[170].dly_stg1  (.A(\tdc0.w_dly_sig[170] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[171] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[170].dly_stg2  (.A(\tdc0.w_dly_sig_n[170] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[172] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[171].dly_stg1  (.A(\tdc0.w_dly_sig[171] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[172] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[171].dly_stg2  (.A(\tdc0.w_dly_sig_n[171] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[173] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[172].dly_stg1  (.A(\tdc0.w_dly_sig[172] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[173] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[172].dly_stg2  (.A(\tdc0.w_dly_sig_n[172] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[174] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[173].dly_stg1  (.A(\tdc0.w_dly_sig[173] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[174] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[173].dly_stg2  (.A(\tdc0.w_dly_sig_n[173] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[175] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[174].dly_stg1  (.A(\tdc0.w_dly_sig[174] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[175] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[174].dly_stg2  (.A(\tdc0.w_dly_sig_n[174] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[176] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[175].dly_stg1  (.A(\tdc0.w_dly_sig[175] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[176] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[175].dly_stg2  (.A(\tdc0.w_dly_sig_n[175] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[177] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[176].dly_stg1  (.A(\tdc0.w_dly_sig[176] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[177] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[176].dly_stg2  (.A(\tdc0.w_dly_sig_n[176] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[178] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[177].dly_stg1  (.A(\tdc0.w_dly_sig[177] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[178] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[177].dly_stg2  (.A(\tdc0.w_dly_sig_n[177] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[179] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[178].dly_stg1  (.A(\tdc0.w_dly_sig[178] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[179] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[178].dly_stg2  (.A(\tdc0.w_dly_sig_n[178] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[180] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[179].dly_stg1  (.A(\tdc0.w_dly_sig[179] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[180] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[179].dly_stg2  (.A(\tdc0.w_dly_sig_n[179] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[181] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[17].dly_stg1  (.A(\tdc0.w_dly_sig[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[18] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[17].dly_stg2  (.A(\tdc0.w_dly_sig_n[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[19] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[180].dly_stg1  (.A(\tdc0.w_dly_sig[180] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[181] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[180].dly_stg2  (.A(\tdc0.w_dly_sig_n[180] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[182] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[181].dly_stg1  (.A(\tdc0.w_dly_sig[181] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[182] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[181].dly_stg2  (.A(\tdc0.w_dly_sig_n[181] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[183] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[182].dly_stg1  (.A(\tdc0.w_dly_sig[182] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[183] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[182].dly_stg2  (.A(\tdc0.w_dly_sig_n[182] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[184] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[183].dly_stg1  (.A(\tdc0.w_dly_sig[183] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[184] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[183].dly_stg2  (.A(\tdc0.w_dly_sig_n[183] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[185] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[184].dly_stg1  (.A(\tdc0.w_dly_sig[184] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[185] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[184].dly_stg2  (.A(\tdc0.w_dly_sig_n[184] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[186] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[185].dly_stg1  (.A(\tdc0.w_dly_sig[185] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[186] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[185].dly_stg2  (.A(\tdc0.w_dly_sig_n[185] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[187] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[186].dly_stg1  (.A(\tdc0.w_dly_sig[186] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[187] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[186].dly_stg2  (.A(\tdc0.w_dly_sig_n[186] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[188] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[187].dly_stg1  (.A(\tdc0.w_dly_sig[187] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[188] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[187].dly_stg2  (.A(\tdc0.w_dly_sig_n[187] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[189] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[188].dly_stg1  (.A(\tdc0.w_dly_sig[188] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[189] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[188].dly_stg2  (.A(\tdc0.w_dly_sig_n[188] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[190] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[189].dly_stg1  (.A(\tdc0.w_dly_sig[189] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[190] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[189].dly_stg2  (.A(\tdc0.w_dly_sig_n[189] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[191] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[18].dly_stg1  (.A(\tdc0.w_dly_sig[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[19] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[18].dly_stg2  (.A(\tdc0.w_dly_sig_n[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[20] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[190].dly_stg1  (.A(\tdc0.w_dly_sig[190] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[191] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[190].dly_stg2  (.A(\tdc0.w_dly_sig_n[190] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[192] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[191].dly_stg1  (.A(\tdc0.w_dly_sig[191] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[192] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[191].dly_stg2  (.A(\tdc0.w_dly_sig_n[191] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[193] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[19].dly_stg1  (.A(\tdc0.w_dly_sig[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[20] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[19].dly_stg2  (.A(\tdc0.w_dly_sig_n[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[21] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[1].dly_stg1  (.A(\tdc0.w_dly_sig[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[2] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[1].dly_stg2  (.A(\tdc0.w_dly_sig_n[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[3] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[20].dly_stg1  (.A(\tdc0.w_dly_sig[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[21] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[20].dly_stg2  (.A(\tdc0.w_dly_sig_n[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[22] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[21].dly_stg1  (.A(\tdc0.w_dly_sig[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[22] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[21].dly_stg2  (.A(\tdc0.w_dly_sig_n[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[23] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[22].dly_stg1  (.A(\tdc0.w_dly_sig[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[23] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[22].dly_stg2  (.A(\tdc0.w_dly_sig_n[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[24] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[23].dly_stg1  (.A(\tdc0.w_dly_sig[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[24] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[23].dly_stg2  (.A(\tdc0.w_dly_sig_n[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[25] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[24].dly_stg1  (.A(\tdc0.w_dly_sig[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[25] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[24].dly_stg2  (.A(\tdc0.w_dly_sig_n[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[26] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[25].dly_stg1  (.A(\tdc0.w_dly_sig[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[26] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[25].dly_stg2  (.A(\tdc0.w_dly_sig_n[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[27] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[26].dly_stg1  (.A(\tdc0.w_dly_sig[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[27] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[26].dly_stg2  (.A(\tdc0.w_dly_sig_n[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[28] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[27].dly_stg1  (.A(\tdc0.w_dly_sig[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[28] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[27].dly_stg2  (.A(\tdc0.w_dly_sig_n[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[29] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[28].dly_stg1  (.A(\tdc0.w_dly_sig[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[29] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[28].dly_stg2  (.A(\tdc0.w_dly_sig_n[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[30] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[29].dly_stg1  (.A(\tdc0.w_dly_sig[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[30] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[29].dly_stg2  (.A(\tdc0.w_dly_sig_n[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[31] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[2].dly_stg1  (.A(\tdc0.w_dly_sig[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[3] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[2].dly_stg2  (.A(\tdc0.w_dly_sig_n[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[4] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[30].dly_stg1  (.A(\tdc0.w_dly_sig[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[31] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[30].dly_stg2  (.A(\tdc0.w_dly_sig_n[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[32] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[31].dly_stg1  (.A(\tdc0.w_dly_sig[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[32] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[31].dly_stg2  (.A(\tdc0.w_dly_sig_n[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[33] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[32].dly_stg1  (.A(\tdc0.w_dly_sig[32] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[33] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[32].dly_stg2  (.A(\tdc0.w_dly_sig_n[32] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[34] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[33].dly_stg1  (.A(\tdc0.w_dly_sig[33] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[34] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[33].dly_stg2  (.A(\tdc0.w_dly_sig_n[33] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[35] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[34].dly_stg1  (.A(\tdc0.w_dly_sig[34] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[35] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[34].dly_stg2  (.A(\tdc0.w_dly_sig_n[34] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[36] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[35].dly_stg1  (.A(\tdc0.w_dly_sig[35] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[36] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[35].dly_stg2  (.A(\tdc0.w_dly_sig_n[35] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[37] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[36].dly_stg1  (.A(\tdc0.w_dly_sig[36] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[37] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[36].dly_stg2  (.A(\tdc0.w_dly_sig_n[36] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[38] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[37].dly_stg1  (.A(\tdc0.w_dly_sig[37] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[38] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[37].dly_stg2  (.A(\tdc0.w_dly_sig_n[37] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[39] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[38].dly_stg1  (.A(\tdc0.w_dly_sig[38] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[39] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[38].dly_stg2  (.A(\tdc0.w_dly_sig_n[38] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[40] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[39].dly_stg1  (.A(\tdc0.w_dly_sig[39] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[40] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[39].dly_stg2  (.A(\tdc0.w_dly_sig_n[39] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[41] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[3].dly_stg1  (.A(\tdc0.w_dly_sig[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[4] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[3].dly_stg2  (.A(\tdc0.w_dly_sig_n[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[5] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[40].dly_stg1  (.A(\tdc0.w_dly_sig[40] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[41] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[40].dly_stg2  (.A(\tdc0.w_dly_sig_n[40] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[42] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[41].dly_stg1  (.A(\tdc0.w_dly_sig[41] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[42] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[41].dly_stg2  (.A(\tdc0.w_dly_sig_n[41] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[43] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[42].dly_stg1  (.A(\tdc0.w_dly_sig[42] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[43] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[42].dly_stg2  (.A(\tdc0.w_dly_sig_n[42] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[44] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[43].dly_stg1  (.A(\tdc0.w_dly_sig[43] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[44] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[43].dly_stg2  (.A(\tdc0.w_dly_sig_n[43] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[45] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[44].dly_stg1  (.A(\tdc0.w_dly_sig[44] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[45] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[44].dly_stg2  (.A(\tdc0.w_dly_sig_n[44] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[46] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[45].dly_stg1  (.A(\tdc0.w_dly_sig[45] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[46] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[45].dly_stg2  (.A(\tdc0.w_dly_sig_n[45] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[47] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[46].dly_stg1  (.A(\tdc0.w_dly_sig[46] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[47] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[46].dly_stg2  (.A(\tdc0.w_dly_sig_n[46] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[48] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[47].dly_stg1  (.A(\tdc0.w_dly_sig[47] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[48] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[47].dly_stg2  (.A(\tdc0.w_dly_sig_n[47] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[49] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[48].dly_stg1  (.A(\tdc0.w_dly_sig[48] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[49] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[48].dly_stg2  (.A(\tdc0.w_dly_sig_n[48] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[50] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[49].dly_stg1  (.A(\tdc0.w_dly_sig[49] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[50] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[49].dly_stg2  (.A(\tdc0.w_dly_sig_n[49] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[51] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[4].dly_stg1  (.A(\tdc0.w_dly_sig[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[5] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[4].dly_stg2  (.A(\tdc0.w_dly_sig_n[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[6] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[50].dly_stg1  (.A(\tdc0.w_dly_sig[50] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[51] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[50].dly_stg2  (.A(\tdc0.w_dly_sig_n[50] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[52] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[51].dly_stg1  (.A(\tdc0.w_dly_sig[51] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[52] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[51].dly_stg2  (.A(\tdc0.w_dly_sig_n[51] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[53] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[52].dly_stg1  (.A(\tdc0.w_dly_sig[52] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[53] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[52].dly_stg2  (.A(\tdc0.w_dly_sig_n[52] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[54] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[53].dly_stg1  (.A(\tdc0.w_dly_sig[53] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[54] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[53].dly_stg2  (.A(\tdc0.w_dly_sig_n[53] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[55] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[54].dly_stg1  (.A(\tdc0.w_dly_sig[54] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[55] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[54].dly_stg2  (.A(\tdc0.w_dly_sig_n[54] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[56] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[55].dly_stg1  (.A(\tdc0.w_dly_sig[55] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[56] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[55].dly_stg2  (.A(\tdc0.w_dly_sig_n[55] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[57] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[56].dly_stg1  (.A(\tdc0.w_dly_sig[56] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[57] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[56].dly_stg2  (.A(\tdc0.w_dly_sig_n[56] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[58] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[57].dly_stg1  (.A(\tdc0.w_dly_sig[57] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[58] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[57].dly_stg2  (.A(\tdc0.w_dly_sig_n[57] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[59] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[58].dly_stg1  (.A(\tdc0.w_dly_sig[58] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[59] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[58].dly_stg2  (.A(\tdc0.w_dly_sig_n[58] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[60] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[59].dly_stg1  (.A(\tdc0.w_dly_sig[59] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[60] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[59].dly_stg2  (.A(\tdc0.w_dly_sig_n[59] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[61] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[5].dly_stg1  (.A(\tdc0.w_dly_sig[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[6] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[5].dly_stg2  (.A(\tdc0.w_dly_sig_n[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[7] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[60].dly_stg1  (.A(\tdc0.w_dly_sig[60] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[61] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[60].dly_stg2  (.A(\tdc0.w_dly_sig_n[60] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[62] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[61].dly_stg1  (.A(\tdc0.w_dly_sig[61] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[62] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[61].dly_stg2  (.A(\tdc0.w_dly_sig_n[61] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[63] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[62].dly_stg1  (.A(\tdc0.w_dly_sig[62] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[63] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[62].dly_stg2  (.A(\tdc0.w_dly_sig_n[62] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[64] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[63].dly_stg1  (.A(\tdc0.w_dly_sig[63] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[64] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[63].dly_stg2  (.A(\tdc0.w_dly_sig_n[63] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[65] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[64].dly_stg1  (.A(\tdc0.w_dly_sig[64] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[65] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[64].dly_stg2  (.A(\tdc0.w_dly_sig_n[64] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[66] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[65].dly_stg1  (.A(\tdc0.w_dly_sig[65] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[66] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[65].dly_stg2  (.A(\tdc0.w_dly_sig_n[65] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[67] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[66].dly_stg1  (.A(\tdc0.w_dly_sig[66] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[67] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[66].dly_stg2  (.A(\tdc0.w_dly_sig_n[66] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[68] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[67].dly_stg1  (.A(\tdc0.w_dly_sig[67] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[68] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[67].dly_stg2  (.A(\tdc0.w_dly_sig_n[67] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[69] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[68].dly_stg1  (.A(\tdc0.w_dly_sig[68] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[69] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[68].dly_stg2  (.A(\tdc0.w_dly_sig_n[68] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[70] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[69].dly_stg1  (.A(\tdc0.w_dly_sig[69] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[70] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[69].dly_stg2  (.A(\tdc0.w_dly_sig_n[69] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[71] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[6].dly_stg1  (.A(\tdc0.w_dly_sig[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[7] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[6].dly_stg2  (.A(\tdc0.w_dly_sig_n[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[8] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[70].dly_stg1  (.A(\tdc0.w_dly_sig[70] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[71] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[70].dly_stg2  (.A(\tdc0.w_dly_sig_n[70] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[72] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[71].dly_stg1  (.A(\tdc0.w_dly_sig[71] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[72] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[71].dly_stg2  (.A(\tdc0.w_dly_sig_n[71] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[73] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[72].dly_stg1  (.A(\tdc0.w_dly_sig[72] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[73] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[72].dly_stg2  (.A(\tdc0.w_dly_sig_n[72] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[74] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[73].dly_stg1  (.A(\tdc0.w_dly_sig[73] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[74] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[73].dly_stg2  (.A(\tdc0.w_dly_sig_n[73] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[75] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[74].dly_stg1  (.A(\tdc0.w_dly_sig[74] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[75] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[74].dly_stg2  (.A(\tdc0.w_dly_sig_n[74] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[76] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[75].dly_stg1  (.A(\tdc0.w_dly_sig[75] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[76] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[75].dly_stg2  (.A(\tdc0.w_dly_sig_n[75] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[77] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[76].dly_stg1  (.A(\tdc0.w_dly_sig[76] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[77] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[76].dly_stg2  (.A(\tdc0.w_dly_sig_n[76] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[78] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[77].dly_stg1  (.A(\tdc0.w_dly_sig[77] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[78] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[77].dly_stg2  (.A(\tdc0.w_dly_sig_n[77] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[79] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[78].dly_stg1  (.A(\tdc0.w_dly_sig[78] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[79] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[78].dly_stg2  (.A(\tdc0.w_dly_sig_n[78] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[80] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[79].dly_stg1  (.A(\tdc0.w_dly_sig[79] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[80] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[79].dly_stg2  (.A(\tdc0.w_dly_sig_n[79] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[81] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[7].dly_stg1  (.A(\tdc0.w_dly_sig[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[8] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[7].dly_stg2  (.A(\tdc0.w_dly_sig_n[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[9] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[80].dly_stg1  (.A(\tdc0.w_dly_sig[80] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[81] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[80].dly_stg2  (.A(\tdc0.w_dly_sig_n[80] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[82] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[81].dly_stg1  (.A(\tdc0.w_dly_sig[81] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[82] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[81].dly_stg2  (.A(\tdc0.w_dly_sig_n[81] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[83] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[82].dly_stg1  (.A(\tdc0.w_dly_sig[82] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[83] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[82].dly_stg2  (.A(\tdc0.w_dly_sig_n[82] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[84] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[83].dly_stg1  (.A(\tdc0.w_dly_sig[83] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[84] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[83].dly_stg2  (.A(\tdc0.w_dly_sig_n[83] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[85] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[84].dly_stg1  (.A(\tdc0.w_dly_sig[84] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[85] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[84].dly_stg2  (.A(\tdc0.w_dly_sig_n[84] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[86] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[85].dly_stg1  (.A(\tdc0.w_dly_sig[85] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[86] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[85].dly_stg2  (.A(\tdc0.w_dly_sig_n[85] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[87] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[86].dly_stg1  (.A(\tdc0.w_dly_sig[86] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[87] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[86].dly_stg2  (.A(\tdc0.w_dly_sig_n[86] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[88] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[87].dly_stg1  (.A(\tdc0.w_dly_sig[87] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[88] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[87].dly_stg2  (.A(\tdc0.w_dly_sig_n[87] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[89] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[88].dly_stg1  (.A(\tdc0.w_dly_sig[88] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[89] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[88].dly_stg2  (.A(\tdc0.w_dly_sig_n[88] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[90] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[89].dly_stg1  (.A(\tdc0.w_dly_sig[89] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[90] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[89].dly_stg2  (.A(\tdc0.w_dly_sig_n[89] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[91] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[8].dly_stg1  (.A(\tdc0.w_dly_sig[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[9] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[8].dly_stg2  (.A(\tdc0.w_dly_sig_n[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[10] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[90].dly_stg1  (.A(\tdc0.w_dly_sig[90] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[91] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[90].dly_stg2  (.A(\tdc0.w_dly_sig_n[90] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[92] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[91].dly_stg1  (.A(\tdc0.w_dly_sig[91] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[92] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[91].dly_stg2  (.A(\tdc0.w_dly_sig_n[91] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[93] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[92].dly_stg1  (.A(\tdc0.w_dly_sig[92] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[93] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[92].dly_stg2  (.A(\tdc0.w_dly_sig_n[92] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[94] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[93].dly_stg1  (.A(\tdc0.w_dly_sig[93] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[94] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[93].dly_stg2  (.A(\tdc0.w_dly_sig_n[93] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[95] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[94].dly_stg1  (.A(\tdc0.w_dly_sig[94] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[95] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[94].dly_stg2  (.A(\tdc0.w_dly_sig_n[94] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[96] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[95].dly_stg1  (.A(\tdc0.w_dly_sig[95] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[96] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[95].dly_stg2  (.A(\tdc0.w_dly_sig_n[95] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[97] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[96].dly_stg1  (.A(\tdc0.w_dly_sig[96] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[97] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[96].dly_stg2  (.A(\tdc0.w_dly_sig_n[96] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[98] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[97].dly_stg1  (.A(\tdc0.w_dly_sig[97] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[98] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[97].dly_stg2  (.A(\tdc0.w_dly_sig_n[97] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[99] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[98].dly_stg1  (.A(\tdc0.w_dly_sig[98] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[99] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[98].dly_stg2  (.A(\tdc0.w_dly_sig_n[98] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[100] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[99].dly_stg1  (.A(\tdc0.w_dly_sig[99] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[100] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[99].dly_stg2  (.A(\tdc0.w_dly_sig_n[99] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[101] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[9].dly_stg1  (.A(\tdc0.w_dly_sig[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig_n[10] ));
 sky130_fd_sc_hd__inv_2 \tdc0.g_dly_chain_interleave[9].dly_stg2  (.A(\tdc0.w_dly_sig_n[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\tdc0.w_dly_sig[11] ));
 sky130_fd_sc_hd__conb_1 tt_um_hpretl_tt06_tdc_10 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net10));
 sky130_fd_sc_hd__conb_1 tt_um_hpretl_tt06_tdc_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net11));
 sky130_fd_sc_hd__conb_1 tt_um_hpretl_tt06_tdc_12 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net12));
 sky130_fd_sc_hd__conb_1 tt_um_hpretl_tt06_tdc_13 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net13));
 sky130_fd_sc_hd__conb_1 tt_um_hpretl_tt06_tdc_14 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net14));
 sky130_fd_sc_hd__conb_1 tt_um_hpretl_tt06_tdc_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net15));
 sky130_fd_sc_hd__conb_1 tt_um_hpretl_tt06_tdc_16 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net16));
 sky130_fd_sc_hd__conb_1 tt_um_hpretl_tt06_tdc_17 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net17));
 sky130_fd_sc_hd__conb_1 tt_um_hpretl_tt06_tdc_18 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net18));
 sky130_fd_sc_hd__conb_1 tt_um_hpretl_tt06_tdc_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net19));
 sky130_fd_sc_hd__conb_1 tt_um_hpretl_tt06_tdc_20 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net20));
 sky130_fd_sc_hd__conb_1 tt_um_hpretl_tt06_tdc_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net21));
 sky130_fd_sc_hd__conb_1 tt_um_hpretl_tt06_tdc_22 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net22));
 sky130_fd_sc_hd__conb_1 tt_um_hpretl_tt06_tdc_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net7));
 sky130_fd_sc_hd__conb_1 tt_um_hpretl_tt06_tdc_8 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net8));
 sky130_fd_sc_hd__conb_1 tt_um_hpretl_tt06_tdc_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net9));
 assign uio_oe[0] = net7;
 assign uio_oe[1] = net8;
 assign uio_oe[2] = net9;
 assign uio_oe[3] = net10;
 assign uio_oe[4] = net11;
 assign uio_oe[5] = net12;
 assign uio_oe[6] = net13;
 assign uio_oe[7] = net14;
 assign uio_out[0] = net15;
 assign uio_out[1] = net16;
 assign uio_out[2] = net17;
 assign uio_out[3] = net18;
 assign uio_out[4] = net19;
 assign uio_out[5] = net20;
 assign uio_out[6] = net21;
 assign uio_out[7] = net22;
endmodule
