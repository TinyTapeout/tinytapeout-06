MACRO tt_um_algofoogle_tt06_grab_bag
  CLASS BLOCK ;
  FOREIGN tt_um_algofoogle_tt06_grab_bag ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 154.870 224.760 155.170 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 158.550 224.760 158.850 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 151.190 224.760 151.490 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.480000 ;
    PORT
      LAYER met4 ;
        RECT 156.560 0.000 157.160 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 134.480 0.000 135.080 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 112.400 0.000 113.000 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 90.320 0.000 90.920 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 68.240 0.000 68.840 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 46.160 0.000 46.760 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 24.080 0.000 24.680 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 2.000 0.000 2.600 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.800000 ;
    PORT
      LAYER met4 ;
        RECT 147.510 224.760 147.810 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 140.150 224.760 140.450 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 136.470 224.760 136.770 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 129.110 224.760 129.410 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 125.430 224.760 125.730 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.070 224.760 118.370 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 114.390 224.760 114.690 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.030 224.760 107.330 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 103.350 224.760 103.650 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 95.990 224.760 96.290 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 92.310 224.760 92.610 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 203.973389 ;
    PORT
      LAYER met4 ;
        RECT 29.750 224.760 30.050 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 203.973389 ;
    PORT
      LAYER met4 ;
        RECT 26.070 224.760 26.370 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 203.973389 ;
    PORT
      LAYER met4 ;
        RECT 22.390 224.760 22.690 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 203.973389 ;
    PORT
      LAYER met4 ;
        RECT 18.710 224.760 19.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 203.973389 ;
    PORT
      LAYER met4 ;
        RECT 15.030 224.760 15.330 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 203.973389 ;
    PORT
      LAYER met4 ;
        RECT 11.350 224.760 11.650 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 203.973389 ;
    PORT
      LAYER met4 ;
        RECT 7.670 224.760 7.970 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 203.973389 ;
    PORT
      LAYER met4 ;
        RECT 3.990 224.760 4.290 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 203.973389 ;
    PORT
      LAYER met4 ;
        RECT 59.190 224.760 59.490 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 203.973389 ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 203.973389 ;
    PORT
      LAYER met4 ;
        RECT 51.830 224.760 52.130 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 203.973389 ;
    PORT
      LAYER met4 ;
        RECT 48.150 224.760 48.450 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 203.973389 ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 203.973389 ;
    PORT
      LAYER met4 ;
        RECT 40.790 224.760 41.090 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 203.973389 ;
    PORT
      LAYER met4 ;
        RECT 37.110 224.760 37.410 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 203.973389 ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.480000 ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 203.973389 ;
    PORT
      LAYER met4 ;
        RECT 84.950 224.760 85.250 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 203.973389 ;
    PORT
      LAYER met4 ;
        RECT 81.270 224.760 81.570 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 203.973389 ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 203.973389 ;
    PORT
      LAYER met4 ;
        RECT 73.910 224.760 74.210 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 203.973389 ;
    PORT
      LAYER met4 ;
        RECT 70.230 224.760 70.530 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 203.973389 ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 203.973389 ;
    PORT
      LAYER met4 ;
        RECT 62.870 224.760 63.170 225.760 ;
    END
  END uo_out[7]
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 2.500 220.760 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 49.000 5.000 50.500 220.760 ;
    END
  END VGND
  OBS
      LAYER pwell ;
        RECT 91.830 156.850 94.180 202.570 ;
        RECT 95.830 156.850 98.180 202.570 ;
        RECT 99.830 156.850 102.180 202.570 ;
        RECT 103.830 156.850 106.180 202.570 ;
        RECT 107.830 156.850 110.180 202.570 ;
        RECT 111.830 156.850 114.180 202.570 ;
        RECT 115.830 156.850 118.180 202.570 ;
        RECT 119.830 156.850 122.180 202.570 ;
        RECT 91.830 129.200 94.180 154.570 ;
        RECT 95.830 129.200 98.180 154.570 ;
        RECT 99.830 129.200 102.180 154.570 ;
        RECT 103.830 129.200 106.180 154.570 ;
        RECT 107.830 129.200 110.180 154.570 ;
        RECT 111.830 129.200 114.180 154.570 ;
        RECT 115.830 129.200 118.180 154.570 ;
        RECT 119.830 129.200 122.180 154.570 ;
      LAYER nwell ;
        RECT 144.215 24.870 146.325 35.060 ;
      LAYER pwell ;
        RECT 147.030 26.935 149.140 33.035 ;
      LAYER li1 ;
        RECT 92.010 202.220 94.000 202.390 ;
        RECT 92.010 178.710 92.180 202.220 ;
        RECT 92.660 199.580 93.350 201.740 ;
        RECT 93.830 178.710 94.000 202.220 ;
        RECT 96.010 202.220 98.000 202.390 ;
        RECT 96.010 178.710 96.180 202.220 ;
        RECT 96.660 199.580 97.350 201.740 ;
        RECT 97.830 178.710 98.000 202.220 ;
        RECT 100.010 202.220 102.000 202.390 ;
        RECT 100.010 178.710 100.180 202.220 ;
        RECT 100.660 199.580 101.350 201.740 ;
        RECT 101.830 178.710 102.000 202.220 ;
        RECT 104.010 202.220 106.000 202.390 ;
        RECT 104.010 178.710 104.180 202.220 ;
        RECT 104.660 199.580 105.350 201.740 ;
        RECT 105.830 178.710 106.000 202.220 ;
        RECT 108.010 202.220 110.000 202.390 ;
        RECT 108.010 178.710 108.180 202.220 ;
        RECT 108.660 199.580 109.350 201.740 ;
        RECT 109.830 178.710 110.000 202.220 ;
        RECT 112.010 202.220 114.000 202.390 ;
        RECT 112.010 178.710 112.180 202.220 ;
        RECT 112.660 199.580 113.350 201.740 ;
        RECT 113.830 178.710 114.000 202.220 ;
        RECT 116.010 202.220 118.000 202.390 ;
        RECT 116.010 178.710 116.180 202.220 ;
        RECT 116.660 199.580 117.350 201.740 ;
        RECT 117.830 178.710 118.000 202.220 ;
        RECT 120.010 202.220 122.000 202.390 ;
        RECT 120.010 178.710 120.180 202.220 ;
        RECT 120.660 199.580 121.350 201.740 ;
        RECT 121.830 178.710 122.000 202.220 ;
        RECT 91.930 177.910 92.270 178.710 ;
        RECT 93.730 177.910 94.070 178.710 ;
        RECT 95.930 177.910 96.270 178.710 ;
        RECT 97.730 177.910 98.070 178.710 ;
        RECT 99.930 177.910 100.270 178.710 ;
        RECT 101.730 177.910 102.070 178.710 ;
        RECT 103.930 177.910 104.270 178.710 ;
        RECT 105.730 177.910 106.070 178.710 ;
        RECT 107.930 177.910 108.270 178.710 ;
        RECT 109.730 177.910 110.070 178.710 ;
        RECT 111.930 177.910 112.270 178.710 ;
        RECT 113.730 177.910 114.070 178.710 ;
        RECT 115.930 177.910 116.270 178.710 ;
        RECT 117.730 177.910 118.070 178.710 ;
        RECT 119.930 177.910 120.270 178.710 ;
        RECT 121.730 177.910 122.070 178.710 ;
        RECT 92.010 157.200 92.180 177.910 ;
        RECT 92.660 157.680 93.350 159.840 ;
        RECT 93.830 157.200 94.000 177.910 ;
        RECT 92.010 157.030 94.000 157.200 ;
        RECT 96.010 157.200 96.180 177.910 ;
        RECT 96.660 157.680 97.350 159.840 ;
        RECT 97.830 157.200 98.000 177.910 ;
        RECT 96.010 157.030 98.000 157.200 ;
        RECT 100.010 157.200 100.180 177.910 ;
        RECT 100.660 157.680 101.350 159.840 ;
        RECT 101.830 157.200 102.000 177.910 ;
        RECT 100.010 157.030 102.000 157.200 ;
        RECT 104.010 157.200 104.180 177.910 ;
        RECT 104.660 157.680 105.350 159.840 ;
        RECT 105.830 157.200 106.000 177.910 ;
        RECT 104.010 157.030 106.000 157.200 ;
        RECT 108.010 157.200 108.180 177.910 ;
        RECT 108.660 157.680 109.350 159.840 ;
        RECT 109.830 157.200 110.000 177.910 ;
        RECT 108.010 157.030 110.000 157.200 ;
        RECT 112.010 157.200 112.180 177.910 ;
        RECT 112.660 157.680 113.350 159.840 ;
        RECT 113.830 157.200 114.000 177.910 ;
        RECT 112.010 157.030 114.000 157.200 ;
        RECT 116.010 157.200 116.180 177.910 ;
        RECT 116.660 157.680 117.350 159.840 ;
        RECT 117.830 157.200 118.000 177.910 ;
        RECT 116.010 157.030 118.000 157.200 ;
        RECT 120.010 157.200 120.180 177.910 ;
        RECT 120.660 157.680 121.350 159.840 ;
        RECT 121.830 157.200 122.000 177.910 ;
        RECT 120.010 157.030 122.000 157.200 ;
        RECT 92.010 154.220 94.000 154.390 ;
        RECT 92.010 129.550 92.180 154.220 ;
        RECT 92.660 151.580 93.350 153.740 ;
        RECT 92.660 130.030 93.350 132.190 ;
        RECT 92.380 129.550 93.640 129.640 ;
        RECT 93.830 129.550 94.000 154.220 ;
        RECT 92.010 129.380 94.000 129.550 ;
        RECT 96.010 154.220 98.000 154.390 ;
        RECT 96.010 129.550 96.180 154.220 ;
        RECT 96.660 151.580 97.350 153.740 ;
        RECT 96.660 130.030 97.350 132.190 ;
        RECT 96.380 129.550 97.640 129.640 ;
        RECT 97.830 129.550 98.000 154.220 ;
        RECT 96.010 129.380 98.000 129.550 ;
        RECT 100.010 154.220 102.000 154.390 ;
        RECT 100.010 129.550 100.180 154.220 ;
        RECT 100.660 151.580 101.350 153.740 ;
        RECT 100.660 130.030 101.350 132.190 ;
        RECT 100.380 129.550 101.640 129.640 ;
        RECT 101.830 129.550 102.000 154.220 ;
        RECT 100.010 129.380 102.000 129.550 ;
        RECT 104.010 154.220 106.000 154.390 ;
        RECT 104.010 129.550 104.180 154.220 ;
        RECT 104.660 151.580 105.350 153.740 ;
        RECT 104.660 130.030 105.350 132.190 ;
        RECT 104.380 129.550 105.640 129.640 ;
        RECT 105.830 129.550 106.000 154.220 ;
        RECT 104.010 129.380 106.000 129.550 ;
        RECT 108.010 154.220 110.000 154.390 ;
        RECT 108.010 129.550 108.180 154.220 ;
        RECT 108.660 151.580 109.350 153.740 ;
        RECT 108.660 130.030 109.350 132.190 ;
        RECT 108.380 129.550 109.640 129.640 ;
        RECT 109.830 129.550 110.000 154.220 ;
        RECT 108.010 129.380 110.000 129.550 ;
        RECT 112.010 154.220 114.000 154.390 ;
        RECT 112.010 129.550 112.180 154.220 ;
        RECT 112.660 151.580 113.350 153.740 ;
        RECT 112.660 130.030 113.350 132.190 ;
        RECT 112.380 129.550 113.640 129.640 ;
        RECT 113.830 129.550 114.000 154.220 ;
        RECT 112.010 129.380 114.000 129.550 ;
        RECT 116.010 154.220 118.000 154.390 ;
        RECT 116.010 129.550 116.180 154.220 ;
        RECT 116.660 151.580 117.350 153.740 ;
        RECT 116.660 130.030 117.350 132.190 ;
        RECT 116.380 129.550 117.640 129.640 ;
        RECT 117.830 129.550 118.000 154.220 ;
        RECT 116.010 129.380 118.000 129.550 ;
        RECT 120.010 154.220 122.000 154.390 ;
        RECT 120.010 129.550 120.180 154.220 ;
        RECT 120.660 151.580 121.350 153.740 ;
        RECT 120.660 130.030 121.350 132.190 ;
        RECT 120.380 129.550 121.640 129.640 ;
        RECT 121.830 129.550 122.000 154.220 ;
        RECT 120.010 129.380 122.000 129.550 ;
        RECT 92.380 129.280 93.640 129.380 ;
        RECT 96.380 129.280 97.640 129.380 ;
        RECT 100.380 129.280 101.640 129.380 ;
        RECT 104.380 129.280 105.640 129.380 ;
        RECT 108.380 129.280 109.640 129.380 ;
        RECT 112.380 129.280 113.640 129.380 ;
        RECT 116.380 129.280 117.640 129.380 ;
        RECT 120.380 129.280 121.640 129.380 ;
        RECT 144.395 34.710 146.145 34.880 ;
        RECT 144.395 30.535 144.565 34.710 ;
        RECT 145.105 34.200 145.435 34.370 ;
        RECT 144.330 29.835 144.630 30.535 ;
        RECT 144.395 25.220 144.565 29.835 ;
        RECT 144.965 25.945 145.135 33.985 ;
        RECT 145.405 25.945 145.575 33.985 ;
        RECT 145.105 25.560 145.435 25.730 ;
        RECT 145.975 25.220 146.145 34.710 ;
        RECT 147.210 32.685 148.960 32.855 ;
        RECT 147.210 27.285 147.380 32.685 ;
        RECT 147.920 32.175 148.250 32.345 ;
        RECT 147.780 27.965 147.950 32.005 ;
        RECT 148.220 27.965 148.390 32.005 ;
        RECT 148.790 31.735 148.960 32.685 ;
        RECT 148.730 30.935 149.030 31.735 ;
        RECT 147.920 27.625 148.250 27.795 ;
        RECT 148.790 27.285 148.960 30.935 ;
        RECT 147.210 27.115 148.960 27.285 ;
        RECT 144.395 25.050 146.145 25.220 ;
      LAYER mcon ;
        RECT 92.740 199.665 93.270 201.650 ;
        RECT 96.740 199.665 97.270 201.650 ;
        RECT 100.740 199.665 101.270 201.650 ;
        RECT 104.740 199.665 105.270 201.650 ;
        RECT 108.740 199.665 109.270 201.650 ;
        RECT 112.740 199.665 113.270 201.650 ;
        RECT 116.740 199.665 117.270 201.650 ;
        RECT 120.740 199.665 121.270 201.650 ;
        RECT 91.930 177.910 92.270 178.710 ;
        RECT 93.730 177.910 94.070 178.710 ;
        RECT 95.930 177.910 96.270 178.710 ;
        RECT 97.730 177.910 98.070 178.710 ;
        RECT 99.930 177.910 100.270 178.710 ;
        RECT 101.730 177.910 102.070 178.710 ;
        RECT 103.930 177.910 104.270 178.710 ;
        RECT 105.730 177.910 106.070 178.710 ;
        RECT 107.930 177.910 108.270 178.710 ;
        RECT 109.730 177.910 110.070 178.710 ;
        RECT 111.930 177.910 112.270 178.710 ;
        RECT 113.730 177.910 114.070 178.710 ;
        RECT 115.930 177.910 116.270 178.710 ;
        RECT 117.730 177.910 118.070 178.710 ;
        RECT 119.930 177.910 120.270 178.710 ;
        RECT 121.730 177.910 122.070 178.710 ;
        RECT 92.740 157.770 93.270 159.755 ;
        RECT 96.740 157.770 97.270 159.755 ;
        RECT 100.740 157.770 101.270 159.755 ;
        RECT 104.740 157.770 105.270 159.755 ;
        RECT 108.740 157.770 109.270 159.755 ;
        RECT 112.740 157.770 113.270 159.755 ;
        RECT 116.740 157.770 117.270 159.755 ;
        RECT 120.740 157.770 121.270 159.755 ;
        RECT 92.740 151.665 93.270 153.650 ;
        RECT 92.740 130.120 93.270 132.105 ;
        RECT 96.740 151.665 97.270 153.650 ;
        RECT 96.740 130.120 97.270 132.105 ;
        RECT 100.740 151.665 101.270 153.650 ;
        RECT 100.740 130.120 101.270 132.105 ;
        RECT 104.740 151.665 105.270 153.650 ;
        RECT 104.740 130.120 105.270 132.105 ;
        RECT 108.740 151.665 109.270 153.650 ;
        RECT 108.740 130.120 109.270 132.105 ;
        RECT 112.740 151.665 113.270 153.650 ;
        RECT 112.740 130.120 113.270 132.105 ;
        RECT 116.740 151.665 117.270 153.650 ;
        RECT 116.740 130.120 117.270 132.105 ;
        RECT 120.740 151.665 121.270 153.650 ;
        RECT 120.740 130.120 121.270 132.105 ;
        RECT 145.185 34.200 145.355 34.370 ;
        RECT 144.330 29.835 144.630 30.535 ;
        RECT 144.965 26.025 145.135 33.905 ;
        RECT 145.405 26.025 145.575 33.905 ;
        RECT 145.185 25.560 145.355 25.730 ;
        RECT 148.000 32.175 148.170 32.345 ;
        RECT 147.780 28.045 147.950 31.925 ;
        RECT 148.220 28.045 148.390 31.925 ;
        RECT 148.730 30.935 149.030 31.735 ;
        RECT 148.000 27.625 148.170 27.795 ;
      LAYER met1 ;
        RECT 88.300 210.300 89.300 216.330 ;
        RECT 88.300 209.300 145.930 210.300 ;
        RECT 54.470 206.900 123.830 207.900 ;
        RECT 92.480 200.070 93.480 206.370 ;
        RECT 96.480 200.070 97.480 206.370 ;
        RECT 100.480 200.070 101.480 206.370 ;
        RECT 104.480 200.070 105.480 206.370 ;
        RECT 108.480 200.070 109.480 206.370 ;
        RECT 112.480 200.070 113.480 206.370 ;
        RECT 116.480 200.070 117.480 206.370 ;
        RECT 92.710 199.605 93.300 200.070 ;
        RECT 96.710 199.605 97.300 200.070 ;
        RECT 100.710 199.605 101.300 200.070 ;
        RECT 104.710 199.605 105.300 200.070 ;
        RECT 108.710 199.605 109.300 200.070 ;
        RECT 112.710 199.605 113.300 200.070 ;
        RECT 116.710 199.605 117.300 200.070 ;
        RECT 118.480 178.850 119.480 206.900 ;
        RECT 120.480 200.070 121.480 206.370 ;
        RECT 120.710 199.605 121.300 200.070 ;
        RECT 118.480 178.820 119.500 178.850 ;
        RECT 91.800 177.820 122.310 178.820 ;
        RECT 118.500 177.790 119.500 177.820 ;
        RECT 92.710 159.390 93.300 159.815 ;
        RECT 96.710 159.390 97.300 159.815 ;
        RECT 100.710 159.390 101.300 159.815 ;
        RECT 104.710 159.390 105.300 159.815 ;
        RECT 108.710 159.390 109.300 159.815 ;
        RECT 112.710 159.390 113.300 159.815 ;
        RECT 116.710 159.390 117.300 159.815 ;
        RECT 120.710 159.390 121.300 159.815 ;
        RECT 92.480 156.270 93.480 159.390 ;
        RECT 86.700 155.270 93.480 156.270 ;
        RECT 86.700 125.300 87.700 155.270 ;
        RECT 92.480 152.170 93.480 155.270 ;
        RECT 96.480 153.170 97.480 159.390 ;
        RECT 100.480 153.170 101.480 159.390 ;
        RECT 104.480 153.170 105.480 159.390 ;
        RECT 108.480 153.170 109.480 159.390 ;
        RECT 112.480 153.170 113.480 159.390 ;
        RECT 116.480 153.170 117.480 159.390 ;
        RECT 120.480 153.170 121.480 159.390 ;
        RECT 94.530 152.170 97.510 153.170 ;
        RECT 98.530 152.170 101.510 153.170 ;
        RECT 102.530 152.170 105.510 153.170 ;
        RECT 106.530 152.170 109.510 153.170 ;
        RECT 110.530 152.170 113.510 153.170 ;
        RECT 114.530 152.170 117.510 153.170 ;
        RECT 118.530 152.170 121.510 153.170 ;
        RECT 92.710 151.605 93.300 152.170 ;
        RECT 92.710 131.680 93.300 132.165 ;
        RECT 94.530 131.680 95.530 152.170 ;
        RECT 96.710 151.605 97.300 152.170 ;
        RECT 96.710 131.680 97.300 132.165 ;
        RECT 98.530 131.680 99.530 152.170 ;
        RECT 100.710 151.605 101.300 152.170 ;
        RECT 100.710 131.680 101.300 132.165 ;
        RECT 102.530 131.680 103.530 152.170 ;
        RECT 104.710 151.605 105.300 152.170 ;
        RECT 104.710 131.680 105.300 132.165 ;
        RECT 106.530 131.680 107.530 152.170 ;
        RECT 108.710 151.605 109.300 152.170 ;
        RECT 108.710 131.680 109.300 132.165 ;
        RECT 110.530 131.680 111.530 152.170 ;
        RECT 112.710 151.605 113.300 152.170 ;
        RECT 112.710 131.680 113.300 132.165 ;
        RECT 114.530 131.680 115.530 152.170 ;
        RECT 116.710 151.605 117.300 152.170 ;
        RECT 116.710 131.680 117.300 132.165 ;
        RECT 118.530 131.680 119.530 152.170 ;
        RECT 120.710 151.605 121.300 152.170 ;
        RECT 92.390 130.680 95.530 131.680 ;
        RECT 96.390 130.680 99.530 131.680 ;
        RECT 100.390 130.680 103.530 131.680 ;
        RECT 104.390 130.680 107.530 131.680 ;
        RECT 108.390 130.680 111.530 131.680 ;
        RECT 112.390 130.680 115.530 131.680 ;
        RECT 116.390 130.680 119.530 131.680 ;
        RECT 120.710 131.670 121.300 132.165 ;
        RECT 122.830 131.670 123.830 206.900 ;
        RECT 92.710 130.060 93.300 130.680 ;
        RECT 96.710 130.060 97.300 130.680 ;
        RECT 100.710 130.060 101.300 130.680 ;
        RECT 104.710 130.060 105.300 130.680 ;
        RECT 108.710 130.060 109.300 130.680 ;
        RECT 112.710 130.060 113.300 130.680 ;
        RECT 116.710 130.060 117.300 130.680 ;
        RECT 120.420 130.670 123.830 131.670 ;
        RECT 120.710 130.060 121.300 130.670 ;
        RECT 91.880 128.770 121.820 129.770 ;
        RECT 86.700 124.300 135.100 125.300 ;
        RECT 134.100 38.870 135.100 124.300 ;
        RECT 147.160 38.430 148.160 222.100 ;
        RECT 149.300 210.300 150.300 210.330 ;
        RECT 149.300 209.300 155.300 210.300 ;
        RECT 149.300 209.270 150.300 209.300 ;
        RECT 147.160 37.430 152.050 38.430 ;
        RECT 147.160 37.400 148.160 37.430 ;
        RECT 57.990 35.185 150.580 36.185 ;
        RECT 145.130 34.400 148.230 34.435 ;
        RECT 145.125 34.170 148.230 34.400 ;
        RECT 145.130 34.135 148.230 34.170 ;
        RECT 144.935 30.685 145.165 33.965 ;
        RECT 145.375 30.935 145.605 33.965 ;
        RECT 147.930 32.435 148.230 34.135 ;
        RECT 149.130 32.435 149.430 32.465 ;
        RECT 147.830 32.135 149.430 32.435 ;
        RECT 149.130 32.105 149.430 32.135 ;
        RECT 147.750 30.935 147.980 31.985 ;
        RECT 148.190 31.835 148.420 31.985 ;
        RECT 149.580 31.835 150.580 35.185 ;
        RECT 10.510 29.685 145.180 30.685 ;
        RECT 145.375 29.685 147.980 30.935 ;
        RECT 148.180 30.835 150.580 31.835 ;
        RECT 144.935 25.965 145.165 29.685 ;
        RECT 145.375 25.965 145.605 29.685 ;
        RECT 146.580 26.435 146.880 29.685 ;
        RECT 147.750 27.985 147.980 29.685 ;
        RECT 148.190 27.985 148.420 30.835 ;
        RECT 151.020 30.450 152.020 37.430 ;
        RECT 149.600 30.435 152.020 30.450 ;
        RECT 149.130 30.085 149.430 30.115 ;
        RECT 149.580 30.085 152.020 30.435 ;
        RECT 149.130 29.785 152.020 30.085 ;
        RECT 149.130 29.755 149.430 29.785 ;
        RECT 149.580 29.460 152.020 29.785 ;
        RECT 149.580 29.435 150.580 29.460 ;
        RECT 149.130 27.835 149.430 27.865 ;
        RECT 147.830 27.535 149.430 27.835 ;
        RECT 147.430 26.435 147.730 26.465 ;
        RECT 146.580 26.135 147.730 26.435 ;
        RECT 147.430 26.105 147.730 26.135 ;
        RECT 147.930 25.785 148.230 27.535 ;
        RECT 149.130 27.505 149.430 27.535 ;
        RECT 149.580 26.435 150.580 26.785 ;
        RECT 148.450 26.135 150.580 26.435 ;
        RECT 145.080 25.485 148.230 25.785 ;
        RECT 149.580 19.910 150.580 26.135 ;
        RECT 154.300 20.200 155.300 209.300 ;
        RECT 154.000 19.910 155.300 20.200 ;
        RECT 149.580 18.910 155.300 19.910 ;
        RECT 149.580 10.350 150.580 18.910 ;
        RECT 152.900 18.900 155.300 18.910 ;
        RECT 156.350 10.350 157.350 10.380 ;
        RECT 149.580 9.350 157.350 10.350 ;
        RECT 156.350 9.320 157.350 9.350 ;
      LAYER via ;
        RECT 147.510 221.750 147.810 222.050 ;
        RECT 88.300 215.300 89.300 216.300 ;
        RECT 144.900 209.300 145.900 210.300 ;
        RECT 54.500 206.900 55.500 207.900 ;
        RECT 92.480 205.340 93.480 206.340 ;
        RECT 96.480 205.340 97.480 206.340 ;
        RECT 100.480 205.340 101.480 206.340 ;
        RECT 104.480 205.340 105.480 206.340 ;
        RECT 108.480 205.340 109.480 206.340 ;
        RECT 112.480 205.340 113.480 206.340 ;
        RECT 116.480 205.340 117.480 206.340 ;
        RECT 120.480 205.340 121.480 206.340 ;
        RECT 118.500 177.820 119.500 178.820 ;
        RECT 118.500 128.770 119.500 129.770 ;
        RECT 134.100 38.900 135.100 39.900 ;
        RECT 58.020 35.185 59.020 36.185 ;
        RECT 149.130 32.135 149.430 32.435 ;
        RECT 10.540 29.685 11.540 30.685 ;
        RECT 149.130 27.535 149.430 27.835 ;
        RECT 147.430 26.135 147.730 26.435 ;
        RECT 148.480 26.135 148.780 26.435 ;
        RECT 156.350 9.350 157.350 10.350 ;
      LAYER met2 ;
        RECT 147.510 222.950 147.810 222.960 ;
        RECT 147.475 222.670 147.845 222.950 ;
        RECT 147.510 221.720 147.810 222.670 ;
        RECT 88.300 216.300 89.300 218.545 ;
        RECT 88.270 215.300 89.330 216.300 ;
        RECT 54.500 207.900 55.500 207.930 ;
        RECT 53.055 206.900 55.500 207.900 ;
        RECT 54.500 206.870 55.500 206.900 ;
        RECT 92.480 206.340 93.480 211.945 ;
        RECT 96.480 206.340 97.480 211.945 ;
        RECT 100.480 206.340 101.480 211.945 ;
        RECT 104.480 206.340 105.480 211.945 ;
        RECT 108.480 206.340 109.480 211.945 ;
        RECT 112.480 206.340 113.480 211.945 ;
        RECT 116.480 206.340 117.480 211.945 ;
        RECT 120.480 206.340 121.480 211.945 ;
        RECT 144.900 210.300 145.900 210.330 ;
        RECT 144.900 209.300 150.330 210.300 ;
        RECT 144.900 209.270 145.900 209.300 ;
        RECT 92.450 205.340 93.510 206.340 ;
        RECT 96.450 205.340 97.510 206.340 ;
        RECT 100.450 205.340 101.510 206.340 ;
        RECT 104.450 205.340 105.510 206.340 ;
        RECT 108.450 205.340 109.510 206.340 ;
        RECT 112.450 205.340 113.510 206.340 ;
        RECT 116.450 205.340 117.510 206.340 ;
        RECT 120.450 205.340 121.510 206.340 ;
        RECT 118.470 177.820 119.530 178.820 ;
        RECT 118.500 128.740 119.500 177.820 ;
        RECT 134.070 38.900 135.130 39.900 ;
        RECT 58.020 36.185 59.020 36.215 ;
        RECT 55.735 35.185 59.020 36.185 ;
        RECT 58.020 35.155 59.020 35.185 ;
        RECT 10.540 30.685 11.540 30.715 ;
        RECT 8.055 29.685 11.540 30.685 ;
        RECT 10.540 29.655 11.540 29.685 ;
        RECT 134.100 7.055 135.100 38.900 ;
        RECT 149.100 32.135 149.460 32.435 ;
        RECT 149.130 30.085 149.430 32.135 ;
        RECT 149.100 29.785 149.460 30.085 ;
        RECT 149.130 27.835 149.430 29.785 ;
        RECT 149.100 27.535 149.460 27.835 ;
        RECT 148.480 26.435 148.780 26.465 ;
        RECT 147.400 26.135 148.780 26.435 ;
        RECT 148.480 26.105 148.780 26.135 ;
        RECT 156.320 9.350 157.380 10.350 ;
        RECT 156.350 7.255 157.350 9.350 ;
      LAYER via2 ;
        RECT 147.520 222.670 147.800 222.950 ;
        RECT 88.300 217.500 89.300 218.500 ;
        RECT 92.480 210.900 93.480 211.900 ;
        RECT 53.100 206.900 54.100 207.900 ;
        RECT 96.480 210.900 97.480 211.900 ;
        RECT 100.480 210.900 101.480 211.900 ;
        RECT 104.480 210.900 105.480 211.900 ;
        RECT 108.480 210.900 109.480 211.900 ;
        RECT 112.480 210.900 113.480 211.900 ;
        RECT 116.480 210.900 117.480 211.900 ;
        RECT 120.480 210.900 121.480 211.900 ;
        RECT 55.780 35.185 56.780 36.185 ;
        RECT 8.100 29.685 9.100 30.685 ;
        RECT 134.100 7.100 135.100 8.100 ;
        RECT 156.350 7.300 157.350 8.300 ;
      LAYER met3 ;
        RECT 147.470 223.760 147.850 224.080 ;
        RECT 147.510 222.975 147.810 223.760 ;
        RECT 147.495 222.645 147.825 222.975 ;
        RECT 88.300 218.525 89.300 220.480 ;
        RECT 88.275 217.475 89.325 218.525 ;
        RECT 92.480 211.925 93.480 214.330 ;
        RECT 96.480 211.925 97.480 214.330 ;
        RECT 100.480 211.925 101.480 214.330 ;
        RECT 104.480 211.925 105.480 214.330 ;
        RECT 108.480 211.925 109.480 214.330 ;
        RECT 112.480 211.925 113.480 214.330 ;
        RECT 116.480 211.925 117.480 214.330 ;
        RECT 120.480 211.925 121.480 214.330 ;
        RECT 92.455 210.875 93.505 211.925 ;
        RECT 96.455 210.875 97.505 211.925 ;
        RECT 100.455 210.875 101.505 211.925 ;
        RECT 104.455 210.875 105.505 211.925 ;
        RECT 108.455 210.875 109.505 211.925 ;
        RECT 112.455 210.875 113.505 211.925 ;
        RECT 116.455 210.875 117.505 211.925 ;
        RECT 120.455 210.875 121.505 211.925 ;
        RECT 53.075 207.900 54.125 207.925 ;
        RECT 51.870 206.900 54.125 207.900 ;
        RECT 53.075 206.875 54.125 206.900 ;
        RECT 55.755 36.185 56.805 36.210 ;
        RECT 53.320 35.185 56.805 36.185 ;
        RECT 55.755 35.160 56.805 35.185 ;
        RECT 8.075 30.685 9.125 30.710 ;
        RECT 5.390 29.685 9.125 30.685 ;
        RECT 8.075 29.660 9.125 29.685 ;
        RECT 134.075 7.075 135.125 8.125 ;
        RECT 156.325 7.275 157.375 8.325 ;
        RECT 134.100 4.670 135.100 7.075 ;
        RECT 156.350 5.170 157.350 7.275 ;
      LAYER via3 ;
        RECT 147.500 223.760 147.820 224.080 ;
        RECT 88.300 219.450 89.300 220.450 ;
        RECT 92.480 213.300 93.480 214.300 ;
        RECT 96.480 213.300 97.480 214.300 ;
        RECT 100.480 213.300 101.480 214.300 ;
        RECT 104.480 213.300 105.480 214.300 ;
        RECT 108.480 213.300 109.480 214.300 ;
        RECT 112.480 213.300 113.480 214.300 ;
        RECT 116.480 213.300 117.480 214.300 ;
        RECT 120.480 213.300 121.480 214.300 ;
        RECT 51.900 206.900 52.900 207.900 ;
        RECT 53.350 35.185 54.350 36.185 ;
        RECT 5.420 29.685 6.420 30.685 ;
        RECT 134.100 4.700 135.100 5.700 ;
        RECT 156.350 5.200 157.350 6.200 ;
      LAYER met4 ;
        RECT 3.990 222.190 4.290 224.760 ;
        RECT 7.670 222.190 7.970 224.760 ;
        RECT 11.350 222.190 11.650 224.760 ;
        RECT 15.030 222.190 15.330 224.760 ;
        RECT 18.710 222.190 19.010 224.760 ;
        RECT 22.390 222.190 22.690 224.760 ;
        RECT 26.070 222.190 26.370 224.760 ;
        RECT 29.750 222.190 30.050 224.760 ;
        RECT 33.430 222.190 33.730 224.760 ;
        RECT 37.110 222.190 37.410 224.760 ;
        RECT 40.790 222.190 41.090 224.760 ;
        RECT 44.470 222.190 44.770 224.760 ;
        RECT 48.150 222.190 48.450 224.760 ;
        RECT 51.830 222.190 52.130 224.760 ;
        RECT 55.510 222.190 55.810 224.760 ;
        RECT 59.190 222.190 59.490 224.760 ;
        RECT 62.870 222.190 63.170 224.760 ;
        RECT 66.550 222.190 66.850 224.760 ;
        RECT 70.230 222.190 70.530 224.760 ;
        RECT 73.910 222.190 74.210 224.760 ;
        RECT 77.590 222.190 77.890 224.760 ;
        RECT 81.270 222.190 81.570 224.760 ;
        RECT 84.950 222.190 85.250 224.760 ;
        RECT 88.630 223.100 88.930 224.760 ;
        RECT 3.740 220.760 85.840 222.190 ;
        RECT 3.740 219.630 49.000 220.760 ;
        RECT 50.500 219.630 85.840 220.760 ;
        RECT 88.300 220.455 89.300 223.100 ;
        RECT 92.310 220.750 92.610 224.760 ;
        RECT 95.990 220.750 96.290 224.760 ;
        RECT 99.670 220.750 99.970 224.760 ;
        RECT 103.350 220.750 103.650 224.760 ;
        RECT 107.030 220.750 107.330 224.760 ;
        RECT 110.710 220.750 111.010 224.760 ;
        RECT 114.390 220.750 114.690 224.760 ;
        RECT 118.070 220.750 118.370 224.760 ;
        RECT 147.510 224.085 147.810 224.760 ;
        RECT 147.495 223.755 147.825 224.085 ;
        RECT 88.295 219.445 89.305 220.455 ;
        RECT 92.310 220.450 93.150 220.750 ;
        RECT 95.990 220.450 97.150 220.750 ;
        RECT 99.670 220.450 101.150 220.750 ;
        RECT 103.350 220.450 105.150 220.750 ;
        RECT 107.030 220.450 109.150 220.750 ;
        RECT 110.710 220.450 113.150 220.750 ;
        RECT 114.390 220.450 117.150 220.750 ;
        RECT 118.070 220.450 121.150 220.750 ;
        RECT 92.850 216.900 93.150 220.450 ;
        RECT 96.850 216.900 97.150 220.450 ;
        RECT 100.850 216.900 101.150 220.450 ;
        RECT 104.850 216.900 105.150 220.450 ;
        RECT 108.850 216.900 109.150 220.450 ;
        RECT 112.850 216.900 113.150 220.450 ;
        RECT 116.850 216.900 117.150 220.450 ;
        RECT 120.850 216.900 121.150 220.450 ;
        RECT 92.480 214.305 93.480 216.900 ;
        RECT 96.480 214.305 97.480 216.900 ;
        RECT 100.480 214.305 101.480 216.900 ;
        RECT 104.480 214.305 105.480 216.900 ;
        RECT 108.480 214.305 109.480 216.900 ;
        RECT 112.480 214.305 113.480 216.900 ;
        RECT 116.480 214.305 117.480 216.900 ;
        RECT 120.480 214.305 121.480 216.900 ;
        RECT 92.475 213.295 93.485 214.305 ;
        RECT 96.475 213.295 97.485 214.305 ;
        RECT 100.475 213.295 101.485 214.305 ;
        RECT 104.475 213.295 105.485 214.305 ;
        RECT 108.475 213.295 109.485 214.305 ;
        RECT 112.475 213.295 113.485 214.305 ;
        RECT 116.475 213.295 117.485 214.305 ;
        RECT 120.475 213.295 121.485 214.305 ;
        RECT 51.895 207.900 52.905 207.905 ;
        RECT 50.500 206.900 52.905 207.900 ;
        RECT 51.895 206.895 52.905 206.900 ;
        RECT 53.345 36.185 54.355 36.190 ;
        RECT 50.500 35.185 54.355 36.185 ;
        RECT 53.345 35.180 54.355 35.185 ;
        RECT 5.415 30.685 6.425 30.690 ;
        RECT 2.500 29.685 6.425 30.685 ;
        RECT 5.415 29.680 6.425 29.685 ;
        RECT 134.095 4.695 135.105 5.705 ;
        RECT 156.345 5.195 157.355 6.205 ;
        RECT 134.100 2.900 135.100 4.695 ;
        RECT 134.480 1.000 135.080 2.900 ;
        RECT 156.430 2.480 157.275 5.195 ;
        RECT 156.560 1.000 157.160 2.480 ;
  END
END tt_um_algofoogle_tt06_grab_bag
END LIBRARY

