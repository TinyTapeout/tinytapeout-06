VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_obriensp_be8
  CLASS BLOCK ;
  FOREIGN tt_um_obriensp_be8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 111.520 ;
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 146.280 2.480 147.880 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 95.080 10.000 96.680 107.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 43.880 10.000 45.480 107.700 ;
    END
  END VGND
  PIN VPWR
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 143.180 10.000 144.780 107.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 120.680 10.000 122.280 107.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 69.480 10.000 71.080 107.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 18.280 10.000 19.880 107.700 ;
    END
  END VPWR
  PIN clk
    ANTENNAGATEAREA 0.852000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 154.870 110.350 155.170 111.520 ;
    END
  END clk
  PIN ena
    PORT
      LAYER met4 ;
        RECT 158.550 110.520 158.850 111.520 ;
    END
  END ena
  PIN rst_n
    ANTENNAGATEAREA 0.585000 ;
    ANTENNADIFFAREA 1.304100 ;
    PORT
      LAYER met4 ;
        RECT 151.190 103.180 151.490 111.520 ;
    END
  END rst_n
  PIN ui_in[0]
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 147.510 110.350 147.810 111.520 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 143.830 110.350 144.130 111.520 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 140.150 102.500 140.450 111.520 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 136.470 110.350 136.770 111.520 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 132.790 94.340 133.090 111.520 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 129.110 110.520 129.410 111.520 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 125.430 110.520 125.730 111.520 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 121.750 110.350 122.050 111.520 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    PORT
      LAYER met4 ;
        RECT 118.070 110.520 118.370 111.520 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    PORT
      LAYER met4 ;
        RECT 114.390 110.520 114.690 111.520 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 110.710 92.300 111.010 111.520 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 107.030 110.350 107.330 111.520 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    PORT
      LAYER met4 ;
        RECT 103.350 110.520 103.650 111.520 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    PORT
      LAYER met4 ;
        RECT 99.670 110.520 99.970 111.520 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    PORT
      LAYER met4 ;
        RECT 95.990 110.520 96.290 111.520 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    PORT
      LAYER met4 ;
        RECT 92.310 110.520 92.610 111.520 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 29.750 96.380 30.050 111.520 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 26.070 96.380 26.370 111.520 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 22.390 78.020 22.690 111.520 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 18.710 110.350 19.010 111.520 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 15.030 52.860 15.330 111.520 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 11.350 94.340 11.650 111.520 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 7.670 90.260 7.970 111.520 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 3.990 94.340 4.290 111.520 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 59.190 103.180 59.490 111.520 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 55.510 109.980 55.810 111.520 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 51.830 110.350 52.130 111.520 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 48.150 110.350 48.450 111.520 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met4 ;
        RECT 44.470 110.520 44.770 111.520 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 40.790 109.980 41.090 111.520 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 37.110 107.940 37.410 111.520 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 33.430 95.020 33.730 111.520 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    ANTENNAGATEAREA 0.252000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met4 ;
        RECT 88.630 89.580 88.930 111.520 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    ANTENNAGATEAREA 0.252000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met4 ;
        RECT 84.950 84.820 85.250 111.520 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    ANTENNAGATEAREA 0.252000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met4 ;
        RECT 81.270 95.700 81.570 111.520 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    ANTENNAGATEAREA 0.252000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met4 ;
        RECT 77.590 91.620 77.890 111.520 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    ANTENNAGATEAREA 0.252000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met4 ;
        RECT 73.910 87.540 74.210 111.520 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    ANTENNAGATEAREA 0.252000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met4 ;
        RECT 70.230 110.350 70.530 111.520 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    ANTENNAGATEAREA 0.252000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met4 ;
        RECT 66.550 90.260 66.850 111.520 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    ANTENNAGATEAREA 0.252000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met4 ;
        RECT 62.870 100.150 63.170 111.520 ;
    END
  END uo_out[7]
  OBS
      LAYER li1 ;
        RECT 2.760 2.635 158.240 108.885 ;
      LAYER met1 ;
        RECT 0.530 0.720 160.930 111.480 ;
      LAYER met2 ;
        RECT 0.560 0.155 160.900 111.510 ;
      LAYER met3 ;
        RECT 0.985 0.175 160.730 111.340 ;
      LAYER met4 ;
        RECT 4.690 93.940 7.270 111.345 ;
        RECT 3.975 89.860 7.270 93.940 ;
        RECT 8.370 93.940 10.950 111.345 ;
        RECT 12.050 93.940 14.630 111.345 ;
        RECT 8.370 89.860 14.630 93.940 ;
        RECT 3.975 52.460 14.630 89.860 ;
        RECT 15.730 109.950 18.310 111.345 ;
        RECT 19.410 109.950 21.990 111.345 ;
        RECT 15.730 108.100 21.990 109.950 ;
        RECT 15.730 52.460 17.880 108.100 ;
        RECT 3.975 9.600 17.880 52.460 ;
        RECT 20.280 77.620 21.990 108.100 ;
        RECT 23.090 95.980 25.670 111.345 ;
        RECT 26.770 95.980 29.350 111.345 ;
        RECT 30.450 95.980 33.030 111.345 ;
        RECT 23.090 94.620 33.030 95.980 ;
        RECT 34.130 107.540 36.710 111.345 ;
        RECT 37.810 109.580 40.390 111.345 ;
        RECT 41.490 110.120 44.070 111.345 ;
        RECT 45.170 110.120 47.750 111.345 ;
        RECT 41.490 109.950 47.750 110.120 ;
        RECT 48.850 109.950 51.430 111.345 ;
        RECT 52.530 109.950 55.110 111.345 ;
        RECT 41.490 109.580 55.110 109.950 ;
        RECT 56.210 109.580 58.790 111.345 ;
        RECT 37.810 108.100 58.790 109.580 ;
        RECT 37.810 107.540 43.480 108.100 ;
        RECT 34.130 94.620 43.480 107.540 ;
        RECT 23.090 77.620 43.480 94.620 ;
        RECT 20.280 9.600 43.480 77.620 ;
        RECT 45.880 102.780 58.790 108.100 ;
        RECT 59.890 102.780 62.470 111.345 ;
        RECT 45.880 99.750 62.470 102.780 ;
        RECT 63.570 99.750 66.150 111.345 ;
        RECT 45.880 89.860 66.150 99.750 ;
        RECT 67.250 109.950 69.830 111.345 ;
        RECT 70.930 109.950 73.510 111.345 ;
        RECT 67.250 108.100 73.510 109.950 ;
        RECT 67.250 89.860 69.080 108.100 ;
        RECT 45.880 9.600 69.080 89.860 ;
        RECT 71.480 87.140 73.510 108.100 ;
        RECT 74.610 91.220 77.190 111.345 ;
        RECT 78.290 95.300 80.870 111.345 ;
        RECT 81.970 95.300 84.550 111.345 ;
        RECT 78.290 91.220 84.550 95.300 ;
        RECT 74.610 87.140 84.550 91.220 ;
        RECT 71.480 84.420 84.550 87.140 ;
        RECT 85.650 89.180 88.230 111.345 ;
        RECT 89.330 110.120 91.910 111.345 ;
        RECT 93.010 110.120 95.590 111.345 ;
        RECT 96.690 110.120 99.270 111.345 ;
        RECT 100.370 110.120 102.950 111.345 ;
        RECT 104.050 110.120 106.630 111.345 ;
        RECT 89.330 109.950 106.630 110.120 ;
        RECT 107.730 109.950 110.310 111.345 ;
        RECT 89.330 108.100 110.310 109.950 ;
        RECT 89.330 89.180 94.680 108.100 ;
        RECT 85.650 84.420 94.680 89.180 ;
        RECT 71.480 9.600 94.680 84.420 ;
        RECT 97.080 91.900 110.310 108.100 ;
        RECT 111.410 110.120 113.990 111.345 ;
        RECT 115.090 110.120 117.670 111.345 ;
        RECT 118.770 110.120 121.350 111.345 ;
        RECT 111.410 109.950 121.350 110.120 ;
        RECT 122.450 110.120 125.030 111.345 ;
        RECT 126.130 110.120 128.710 111.345 ;
        RECT 129.810 110.120 132.390 111.345 ;
        RECT 122.450 109.950 132.390 110.120 ;
        RECT 111.410 108.100 132.390 109.950 ;
        RECT 111.410 91.900 120.280 108.100 ;
        RECT 97.080 9.600 120.280 91.900 ;
        RECT 122.680 93.940 132.390 108.100 ;
        RECT 133.490 109.950 136.070 111.345 ;
        RECT 137.170 109.950 139.750 111.345 ;
        RECT 133.490 102.100 139.750 109.950 ;
        RECT 140.850 109.950 143.430 111.345 ;
        RECT 144.530 109.950 147.110 111.345 ;
        RECT 148.210 109.950 150.790 111.345 ;
        RECT 140.850 109.440 150.790 109.950 ;
        RECT 140.850 108.100 145.880 109.440 ;
        RECT 140.850 102.100 142.780 108.100 ;
        RECT 133.490 93.940 142.780 102.100 ;
        RECT 122.680 9.600 142.780 93.940 ;
        RECT 145.180 9.600 145.880 108.100 ;
        RECT 3.975 2.080 145.880 9.600 ;
        RECT 148.280 102.780 150.790 109.440 ;
        RECT 151.890 109.950 154.470 111.345 ;
        RECT 155.570 110.120 158.150 111.345 ;
        RECT 159.250 110.120 160.705 111.345 ;
        RECT 155.570 109.950 160.705 110.120 ;
        RECT 151.890 102.780 160.705 109.950 ;
        RECT 148.280 2.080 160.705 102.780 ;
        RECT 3.975 0.855 160.705 2.080 ;
  END
END tt_um_obriensp_be8
END LIBRARY

