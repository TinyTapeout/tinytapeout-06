VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_dsatizabal_opamp
  CLASS BLOCK ;
  FOREIGN tt_um_dsatizabal_opamp ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 154.870 224.760 155.170 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 158.550 224.760 158.850 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 151.190 224.760 151.490 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.740000 ;
    PORT
      LAYER met4 ;
        RECT 156.560 0.000 157.160 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.600000 ;
    PORT
      LAYER met4 ;
        RECT 134.480 0.000 135.080 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.600000 ;
    PORT
      LAYER met4 ;
        RECT 112.400 0.000 113.000 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.480000 ;
    PORT
      LAYER met4 ;
        RECT 90.320 0.000 90.920 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 68.240 0.000 68.840 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 46.160 0.000 46.760 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 24.080 0.000 24.680 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 2.000 0.000 2.600 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 147.510 224.760 147.810 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 140.150 224.760 140.450 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 136.470 224.760 136.770 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 129.110 224.760 129.410 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 125.430 224.760 125.730 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.070 224.760 118.370 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 114.390 224.760 114.690 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.030 224.760 107.330 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 103.350 224.760 103.650 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 95.990 224.760 96.290 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 92.310 224.760 92.610 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 10.800000 ;
    ANTENNADIFFAREA 16.202000 ;
    PORT
      LAYER met4 ;
        RECT 29.750 224.760 30.050 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 10.800000 ;
    ANTENNADIFFAREA 16.202000 ;
    PORT
      LAYER met4 ;
        RECT 26.070 224.760 26.370 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 10.800000 ;
    ANTENNADIFFAREA 16.202000 ;
    PORT
      LAYER met4 ;
        RECT 22.390 224.760 22.690 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 10.800000 ;
    ANTENNADIFFAREA 16.202000 ;
    PORT
      LAYER met4 ;
        RECT 18.710 224.760 19.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 10.800000 ;
    ANTENNADIFFAREA 16.202000 ;
    PORT
      LAYER met4 ;
        RECT 15.030 224.760 15.330 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 10.800000 ;
    ANTENNADIFFAREA 16.202000 ;
    PORT
      LAYER met4 ;
        RECT 11.350 224.760 11.650 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 10.800000 ;
    ANTENNADIFFAREA 16.202000 ;
    PORT
      LAYER met4 ;
        RECT 7.670 224.760 7.970 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 10.800000 ;
    ANTENNADIFFAREA 16.202000 ;
    PORT
      LAYER met4 ;
        RECT 3.990 224.760 4.290 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 10.800000 ;
    ANTENNADIFFAREA 16.202000 ;
    PORT
      LAYER met4 ;
        RECT 59.190 224.760 59.490 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 10.800000 ;
    ANTENNADIFFAREA 16.202000 ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 10.800000 ;
    ANTENNADIFFAREA 16.202000 ;
    PORT
      LAYER met4 ;
        RECT 51.830 224.760 52.130 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 10.800000 ;
    ANTENNADIFFAREA 16.202000 ;
    PORT
      LAYER met4 ;
        RECT 48.150 224.760 48.450 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 10.800000 ;
    ANTENNADIFFAREA 16.202000 ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 10.800000 ;
    ANTENNADIFFAREA 16.202000 ;
    PORT
      LAYER met4 ;
        RECT 40.790 224.760 41.090 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 10.800000 ;
    ANTENNADIFFAREA 16.202000 ;
    PORT
      LAYER met4 ;
        RECT 37.110 224.760 37.410 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 10.800000 ;
    ANTENNADIFFAREA 16.202000 ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 10.800000 ;
    ANTENNADIFFAREA 16.202000 ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 10.800000 ;
    ANTENNADIFFAREA 16.202000 ;
    PORT
      LAYER met4 ;
        RECT 84.950 224.760 85.250 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 10.800000 ;
    ANTENNADIFFAREA 16.202000 ;
    PORT
      LAYER met4 ;
        RECT 81.270 224.760 81.570 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 10.800000 ;
    ANTENNADIFFAREA 16.202000 ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 10.800000 ;
    ANTENNADIFFAREA 16.202000 ;
    PORT
      LAYER met4 ;
        RECT 73.910 224.760 74.210 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 10.800000 ;
    ANTENNADIFFAREA 16.202000 ;
    PORT
      LAYER met4 ;
        RECT 70.230 224.760 70.530 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 10.800000 ;
    ANTENNADIFFAREA 16.202000 ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 10.800000 ;
    ANTENNADIFFAREA 16.202000 ;
    PORT
      LAYER met4 ;
        RECT 62.870 224.760 63.170 225.760 ;
    END
  END uo_out[7]
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 2.500 220.760 ;
    END
  END VPWR
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 49.000 14.360 50.500 224.120 ;
    END
  END VGND
  OBS
      LAYER pwell ;
        RECT 110.270 21.950 118.370 24.270 ;
        RECT 110.270 21.710 120.890 21.950 ;
        RECT 118.330 18.850 120.890 21.710 ;
        RECT 121.130 20.420 136.800 22.980 ;
      LAYER nwell ;
        RECT 121.010 17.840 136.860 20.400 ;
        RECT 110.180 14.580 118.370 17.140 ;
        RECT 121.010 13.930 136.860 16.490 ;
      LAYER li1 ;
        RECT 136.960 25.175 137.960 25.460 ;
        RECT 110.450 23.920 118.190 24.090 ;
        RECT 110.450 22.060 110.620 23.920 ;
        RECT 111.300 23.350 117.340 23.520 ;
        RECT 110.960 22.690 111.130 23.290 ;
        RECT 117.510 22.690 117.680 23.290 ;
        RECT 111.300 22.460 117.340 22.630 ;
        RECT 118.020 22.060 118.190 23.920 ;
        RECT 110.450 21.890 118.190 22.060 ;
        RECT 121.310 22.630 136.620 22.800 ;
        RECT 118.510 21.600 120.710 21.770 ;
        RECT 118.510 19.200 118.680 21.600 ;
        RECT 119.310 21.090 119.910 21.260 ;
        RECT 119.080 19.880 119.250 20.920 ;
        RECT 119.970 19.880 120.140 20.920 ;
        RECT 119.310 19.540 119.910 19.710 ;
        RECT 120.540 19.200 120.710 21.600 ;
        RECT 121.310 20.770 121.480 22.630 ;
        RECT 122.160 22.060 128.200 22.230 ;
        RECT 121.820 21.400 121.990 22.000 ;
        RECT 128.370 21.400 128.540 22.000 ;
        RECT 122.160 21.170 128.200 21.340 ;
        RECT 128.880 20.770 129.050 22.630 ;
        RECT 129.730 22.060 135.770 22.230 ;
        RECT 129.390 21.400 129.560 22.000 ;
        RECT 135.940 21.400 136.110 22.000 ;
        RECT 129.730 21.170 135.770 21.340 ;
        RECT 136.450 20.770 136.620 22.630 ;
        RECT 121.310 20.600 136.620 20.770 ;
        RECT 118.510 19.030 120.710 19.200 ;
        RECT 121.190 20.050 136.680 20.220 ;
        RECT 121.190 18.190 121.360 20.050 ;
        RECT 122.085 19.480 128.125 19.650 ;
        RECT 121.700 18.820 121.870 19.420 ;
        RECT 128.340 18.820 128.510 19.420 ;
        RECT 122.085 18.590 128.125 18.760 ;
        RECT 128.850 18.190 129.020 20.050 ;
        RECT 129.745 19.480 135.785 19.650 ;
        RECT 129.360 18.820 129.530 19.420 ;
        RECT 136.000 18.820 136.170 19.420 ;
        RECT 129.745 18.590 135.785 18.760 ;
        RECT 136.510 18.190 136.680 20.050 ;
        RECT 136.960 20.170 137.960 20.175 ;
        RECT 139.170 20.170 140.070 22.080 ;
        RECT 136.960 20.020 140.070 20.170 ;
        RECT 136.960 19.890 140.080 20.020 ;
        RECT 136.960 19.885 137.960 19.890 ;
        RECT 121.190 18.020 136.680 18.190 ;
        RECT 110.360 16.790 118.190 16.960 ;
        RECT 110.360 14.930 110.530 16.790 ;
        RECT 111.255 16.220 117.295 16.390 ;
        RECT 110.870 15.560 111.040 16.160 ;
        RECT 117.510 15.560 117.680 16.160 ;
        RECT 111.255 15.330 117.295 15.500 ;
        RECT 118.020 14.930 118.190 16.790 ;
        RECT 110.360 14.760 118.190 14.930 ;
        RECT 121.190 16.140 136.680 16.310 ;
        RECT 121.190 14.280 121.360 16.140 ;
        RECT 122.085 15.570 128.125 15.740 ;
        RECT 121.700 14.910 121.870 15.510 ;
        RECT 128.340 14.910 128.510 15.510 ;
        RECT 122.085 14.680 128.125 14.850 ;
        RECT 128.850 14.280 129.020 16.140 ;
        RECT 129.745 15.570 135.785 15.740 ;
        RECT 129.360 14.910 129.530 15.510 ;
        RECT 136.000 14.910 136.170 15.510 ;
        RECT 129.745 14.680 135.785 14.850 ;
        RECT 136.510 14.280 136.680 16.140 ;
        RECT 139.170 15.590 140.080 19.890 ;
        RECT 136.960 14.600 137.960 14.885 ;
        RECT 121.190 14.110 136.680 14.280 ;
      LAYER mcon ;
        RECT 137.030 25.230 137.900 25.400 ;
        RECT 113.140 23.920 115.700 24.090 ;
        RECT 111.380 23.350 117.260 23.520 ;
        RECT 110.960 22.770 111.130 23.210 ;
        RECT 117.510 22.770 117.680 23.210 ;
        RECT 111.380 22.460 117.260 22.630 ;
        RECT 124.520 22.630 125.570 22.800 ;
        RECT 132.050 22.630 133.600 22.800 ;
        RECT 119.380 21.600 119.850 21.770 ;
        RECT 119.390 21.090 119.830 21.260 ;
        RECT 119.080 19.960 119.250 20.840 ;
        RECT 119.970 19.960 120.140 20.840 ;
        RECT 119.390 19.540 119.830 19.710 ;
        RECT 122.240 22.060 128.120 22.230 ;
        RECT 121.820 21.480 121.990 21.920 ;
        RECT 128.370 21.480 128.540 21.920 ;
        RECT 122.240 21.170 128.120 21.340 ;
        RECT 129.810 22.060 135.690 22.230 ;
        RECT 129.390 21.480 129.560 21.920 ;
        RECT 135.940 21.480 136.110 21.920 ;
        RECT 129.810 21.170 135.690 21.340 ;
        RECT 139.340 21.280 139.890 21.880 ;
        RECT 122.165 19.480 128.045 19.650 ;
        RECT 121.700 18.900 121.870 19.340 ;
        RECT 128.340 18.900 128.510 19.340 ;
        RECT 122.165 18.590 128.045 18.760 ;
        RECT 129.825 19.480 135.705 19.650 ;
        RECT 129.360 18.900 129.530 19.340 ;
        RECT 136.000 18.900 136.170 19.340 ;
        RECT 129.825 18.590 135.705 18.760 ;
        RECT 124.620 18.020 125.500 18.190 ;
        RECT 131.890 18.020 133.920 18.190 ;
        RECT 111.335 16.220 117.215 16.390 ;
        RECT 110.870 15.640 111.040 16.080 ;
        RECT 117.510 15.640 117.680 16.080 ;
        RECT 111.335 15.330 117.215 15.500 ;
        RECT 113.190 14.760 115.570 14.930 ;
        RECT 122.165 15.570 128.045 15.740 ;
        RECT 121.700 14.990 121.870 15.430 ;
        RECT 128.340 14.990 128.510 15.430 ;
        RECT 122.165 14.680 128.045 14.850 ;
        RECT 129.825 15.570 135.705 15.740 ;
        RECT 129.360 14.990 129.530 15.430 ;
        RECT 136.000 14.990 136.170 15.430 ;
        RECT 129.825 14.680 135.705 14.850 ;
        RECT 139.230 15.660 140.010 15.940 ;
        RECT 137.030 14.650 137.850 14.830 ;
        RECT 124.220 14.110 126.150 14.280 ;
        RECT 131.890 14.110 133.910 14.280 ;
      LAYER met1 ;
        RECT 136.970 27.730 137.970 27.740 ;
        RECT 53.580 26.710 137.970 27.730 ;
        RECT 136.970 25.480 137.970 26.710 ;
        RECT 116.130 25.470 118.140 25.480 ;
        RECT 136.970 25.470 138.780 25.480 ;
        RECT 116.130 25.460 138.780 25.470 ;
        RECT 112.650 25.180 138.780 25.460 ;
        RECT 112.650 25.170 119.910 25.180 ;
        RECT 90.320 19.520 104.720 19.730 ;
        RECT 105.950 19.520 106.970 25.090 ;
        RECT 112.650 23.550 116.160 25.170 ;
        RECT 111.320 23.320 117.320 23.550 ;
        RECT 110.930 23.070 111.160 23.270 ;
        RECT 117.480 23.070 117.710 23.270 ;
        RECT 118.460 23.070 119.000 23.160 ;
        RECT 110.930 22.860 119.000 23.070 ;
        RECT 110.930 22.710 111.160 22.860 ;
        RECT 117.440 22.850 119.000 22.860 ;
        RECT 117.480 22.710 117.710 22.850 ;
        RECT 118.460 22.740 119.000 22.850 ;
        RECT 111.320 22.430 117.320 22.660 ;
        RECT 113.230 19.520 115.240 22.430 ;
        RECT 119.270 21.820 119.910 25.170 ;
        RECT 120.700 22.770 121.130 23.170 ;
        RECT 119.260 21.560 119.910 21.820 ;
        RECT 119.330 21.060 119.890 21.290 ;
        RECT 119.050 20.750 119.280 20.900 ;
        RECT 116.350 20.080 119.280 20.750 ;
        RECT 119.050 19.900 119.280 20.080 ;
        RECT 119.450 19.740 119.730 21.060 ;
        RECT 119.940 20.590 120.170 20.900 ;
        RECT 120.890 20.590 121.130 22.770 ;
        RECT 124.420 22.260 125.670 25.180 ;
        RECT 131.660 22.260 134.160 25.180 ;
        RECT 136.970 25.170 138.780 25.180 ;
        RECT 138.310 25.070 138.780 25.170 ;
        RECT 122.180 22.030 128.180 22.260 ;
        RECT 129.750 22.030 135.750 22.260 ;
        RECT 121.790 21.850 122.020 21.980 ;
        RECT 128.340 21.850 128.570 21.980 ;
        RECT 129.360 21.850 129.590 21.980 ;
        RECT 135.910 21.850 136.140 21.980 ;
        RECT 121.790 21.600 136.140 21.850 ;
        RECT 121.790 21.420 122.020 21.600 ;
        RECT 128.340 21.420 128.570 21.600 ;
        RECT 129.360 21.420 129.590 21.600 ;
        RECT 131.660 21.370 134.160 21.600 ;
        RECT 135.910 21.420 136.140 21.600 ;
        RECT 139.170 21.740 140.090 22.080 ;
        RECT 142.470 21.740 157.150 22.080 ;
        RECT 139.170 21.420 157.150 21.740 ;
        RECT 122.180 21.140 128.180 21.370 ;
        RECT 129.750 21.140 135.750 21.370 ;
        RECT 124.420 20.590 125.660 21.140 ;
        RECT 119.940 20.220 125.660 20.590 ;
        RECT 119.940 19.900 120.170 20.220 ;
        RECT 90.320 18.960 115.240 19.520 ;
        RECT 119.330 19.510 119.890 19.740 ;
        RECT 124.420 19.680 125.660 20.220 ;
        RECT 131.660 19.680 134.160 21.140 ;
        RECT 139.170 21.080 140.090 21.420 ;
        RECT 142.470 21.080 157.150 21.420 ;
        RECT 90.320 18.730 104.720 18.960 ;
        RECT 90.320 18.290 91.850 18.730 ;
        RECT 113.230 16.420 115.240 18.960 ;
        RECT 111.275 16.190 117.275 16.420 ;
        RECT 110.840 15.980 111.070 16.140 ;
        RECT 117.480 15.980 117.710 16.140 ;
        RECT 110.840 15.750 118.940 15.980 ;
        RECT 110.840 15.580 111.070 15.750 ;
        RECT 117.480 15.580 117.710 15.750 ;
        RECT 111.275 15.300 117.275 15.530 ;
        RECT 118.760 15.390 118.940 15.750 ;
        RECT 112.600 13.860 116.080 15.300 ;
        RECT 118.580 15.020 119.070 15.390 ;
        RECT 119.450 13.860 119.730 19.510 ;
        RECT 122.105 19.450 128.105 19.680 ;
        RECT 129.765 19.450 135.765 19.680 ;
        RECT 121.680 19.400 121.880 19.420 ;
        RECT 121.670 19.240 121.900 19.400 ;
        RECT 128.310 19.240 128.540 19.400 ;
        RECT 121.670 19.030 128.540 19.240 ;
        RECT 121.670 18.840 121.900 19.030 ;
        RECT 128.310 18.840 128.540 19.030 ;
        RECT 129.330 19.310 129.560 19.400 ;
        RECT 135.970 19.310 136.200 19.400 ;
        RECT 129.330 19.300 136.200 19.310 ;
        RECT 142.460 19.300 154.190 19.590 ;
        RECT 129.330 18.930 154.190 19.300 ;
        RECT 129.330 18.840 129.560 18.930 ;
        RECT 135.970 18.840 136.200 18.930 ;
        RECT 121.680 17.080 121.880 18.840 ;
        RECT 122.105 18.560 128.105 18.790 ;
        RECT 129.765 18.560 135.765 18.790 ;
        RECT 142.460 18.590 154.190 18.930 ;
        RECT 124.430 17.840 125.650 18.560 ;
        RECT 131.680 17.840 134.160 18.560 ;
        RECT 124.430 17.520 134.160 17.840 ;
        RECT 121.680 16.740 122.090 17.080 ;
        RECT 124.430 15.770 125.650 17.520 ;
        RECT 142.480 17.080 149.020 17.400 ;
        RECT 126.820 16.740 149.020 17.080 ;
        RECT 142.480 16.400 149.020 16.740 ;
        RECT 139.170 15.900 140.080 16.020 ;
        RECT 129.820 15.770 140.080 15.900 ;
        RECT 122.105 15.540 128.105 15.770 ;
        RECT 129.765 15.740 140.080 15.770 ;
        RECT 129.765 15.540 135.765 15.740 ;
        RECT 139.170 15.590 140.080 15.740 ;
        RECT 120.040 15.300 120.620 15.390 ;
        RECT 121.670 15.300 121.900 15.490 ;
        RECT 128.310 15.300 128.540 15.490 ;
        RECT 129.330 15.300 129.560 15.490 ;
        RECT 135.970 15.300 136.200 15.490 ;
        RECT 138.310 15.300 138.780 15.420 ;
        RECT 120.040 15.090 138.780 15.300 ;
        RECT 120.040 15.080 121.910 15.090 ;
        RECT 120.040 15.010 120.620 15.080 ;
        RECT 121.670 14.930 121.900 15.080 ;
        RECT 128.310 14.930 128.540 15.090 ;
        RECT 129.330 14.930 129.560 15.090 ;
        RECT 135.970 14.930 136.200 15.090 ;
        RECT 122.105 14.650 128.105 14.880 ;
        RECT 129.765 14.650 135.765 14.880 ;
        RECT 122.130 13.900 128.090 14.650 ;
        RECT 122.120 13.860 128.090 13.900 ;
        RECT 129.800 13.860 135.730 14.650 ;
        RECT 136.960 13.860 137.970 14.890 ;
        RECT 112.600 13.430 137.970 13.860 ;
        RECT 115.930 13.420 137.970 13.430 ;
        RECT 136.960 13.000 137.970 13.420 ;
        RECT 95.380 11.980 137.970 13.000 ;
        RECT 148.260 8.120 149.020 16.400 ;
        RECT 112.390 7.310 149.020 8.120 ;
        RECT 153.280 5.240 154.190 18.590 ;
        RECT 134.480 4.460 154.190 5.240 ;
      LAYER via ;
        RECT 53.690 26.830 55.260 27.580 ;
        RECT 106.020 23.360 106.880 25.000 ;
        RECT 90.460 18.420 91.720 19.590 ;
        RECT 118.520 22.800 118.950 23.100 ;
        RECT 120.740 22.820 121.080 23.120 ;
        RECT 116.410 20.140 117.500 20.670 ;
        RECT 138.340 25.110 138.740 25.430 ;
        RECT 155.920 21.190 157.050 21.950 ;
        RECT 118.610 15.070 119.030 15.340 ;
        RECT 121.710 16.780 122.050 17.050 ;
        RECT 126.860 16.760 127.520 17.060 ;
        RECT 120.080 15.050 120.580 15.340 ;
        RECT 138.340 15.120 138.740 15.380 ;
        RECT 95.550 12.150 96.810 12.810 ;
        RECT 112.530 7.410 113.970 8.030 ;
        RECT 134.600 4.590 135.510 5.130 ;
      LAYER met2 ;
        RECT 53.570 26.700 55.390 27.740 ;
        RECT 105.930 23.250 106.970 25.090 ;
        RECT 118.460 23.080 119.000 23.160 ;
        RECT 120.700 23.080 121.130 23.170 ;
        RECT 118.460 22.850 121.130 23.080 ;
        RECT 118.460 22.740 119.000 22.850 ;
        RECT 120.700 22.770 121.130 22.850 ;
        RECT 116.350 20.080 117.580 20.750 ;
        RECT 90.320 18.280 91.860 19.740 ;
        RECT 121.680 16.740 127.590 17.080 ;
        RECT 118.580 15.300 119.070 15.390 ;
        RECT 120.040 15.300 120.620 15.390 ;
        RECT 118.580 15.080 120.620 15.300 ;
        RECT 138.310 15.090 138.780 25.480 ;
        RECT 155.770 21.080 157.160 22.080 ;
        RECT 118.580 15.020 119.070 15.080 ;
        RECT 120.040 15.010 120.620 15.080 ;
        RECT 5.810 13.000 56.270 13.040 ;
        RECT 5.810 11.970 96.990 13.000 ;
        RECT 55.460 11.960 96.990 11.970 ;
        RECT 112.390 7.310 114.080 8.120 ;
        RECT 134.480 4.460 135.610 5.240 ;
      LAYER via2 ;
        RECT 53.690 26.830 55.260 27.580 ;
        RECT 106.020 23.360 106.880 25.000 ;
        RECT 116.410 20.140 117.500 20.670 ;
        RECT 90.460 18.420 91.720 19.590 ;
        RECT 155.920 21.190 157.050 21.950 ;
        RECT 5.920 12.070 7.290 12.910 ;
        RECT 112.530 7.410 113.970 8.030 ;
        RECT 134.600 4.590 135.510 5.130 ;
      LAYER met3 ;
        RECT 53.570 26.700 55.390 27.740 ;
        RECT 114.440 26.240 133.850 41.640 ;
        RECT 105.930 23.250 106.970 25.090 ;
        RECT 155.770 21.080 157.160 22.080 ;
        RECT 116.350 20.080 117.580 20.750 ;
        RECT 90.320 18.280 91.860 19.740 ;
        RECT 5.810 11.970 7.390 13.040 ;
        RECT 112.390 7.310 114.080 8.120 ;
        RECT 134.480 4.460 135.610 5.240 ;
      LAYER via3 ;
        RECT 53.690 26.830 55.260 27.580 ;
        RECT 114.540 26.380 114.860 41.500 ;
        RECT 106.020 23.360 106.880 25.000 ;
        RECT 155.920 21.190 157.050 21.950 ;
        RECT 116.410 20.140 117.500 20.670 ;
        RECT 90.460 18.420 91.720 19.590 ;
        RECT 5.920 12.070 7.290 12.910 ;
        RECT 112.530 7.410 113.970 8.030 ;
        RECT 134.600 4.590 135.510 5.130 ;
      LAYER met4 ;
        RECT 3.990 224.120 4.290 224.760 ;
        RECT 7.670 224.120 7.970 224.760 ;
        RECT 11.350 224.120 11.650 224.760 ;
        RECT 15.030 224.120 15.330 224.760 ;
        RECT 18.710 224.120 19.010 224.760 ;
        RECT 22.390 224.120 22.690 224.760 ;
        RECT 26.070 224.120 26.370 224.760 ;
        RECT 29.750 224.120 30.050 224.760 ;
        RECT 33.430 224.120 33.730 224.760 ;
        RECT 37.110 224.120 37.410 224.760 ;
        RECT 40.790 224.120 41.090 224.760 ;
        RECT 44.470 224.120 44.770 224.760 ;
        RECT 48.150 224.120 48.450 224.760 ;
        RECT 51.830 224.120 52.130 224.760 ;
        RECT 55.510 224.120 55.810 224.760 ;
        RECT 59.190 224.120 59.490 224.760 ;
        RECT 62.870 224.120 63.170 224.760 ;
        RECT 66.550 224.120 66.850 224.760 ;
        RECT 70.230 224.120 70.530 224.760 ;
        RECT 73.910 224.120 74.210 224.760 ;
        RECT 77.590 224.120 77.890 224.760 ;
        RECT 81.270 224.120 81.570 224.760 ;
        RECT 84.950 224.120 85.250 224.760 ;
        RECT 88.630 224.120 88.930 224.760 ;
        RECT 92.310 224.510 92.610 224.760 ;
        RECT 95.990 224.510 96.290 224.760 ;
        RECT 99.670 224.510 99.970 224.760 ;
        RECT 103.350 224.510 103.650 224.760 ;
        RECT 107.030 224.510 107.330 224.760 ;
        RECT 110.710 224.510 111.010 224.760 ;
        RECT 114.390 224.510 114.690 224.760 ;
        RECT 118.070 224.510 118.370 224.760 ;
        RECT 121.750 224.510 122.050 224.760 ;
        RECT 125.430 224.510 125.730 224.760 ;
        RECT 129.110 224.510 129.410 224.760 ;
        RECT 132.790 224.510 133.090 224.760 ;
        RECT 136.470 224.510 136.770 224.760 ;
        RECT 140.150 224.510 140.450 224.760 ;
        RECT 143.830 224.510 144.130 224.760 ;
        RECT 147.510 224.510 147.810 224.760 ;
        RECT 151.190 224.510 151.490 224.760 ;
        RECT 154.870 224.510 155.170 224.760 ;
        RECT 158.550 224.510 158.850 224.760 ;
        RECT 3.990 223.090 49.000 224.120 ;
        RECT 50.500 223.090 88.940 224.120 ;
        RECT 114.460 35.460 114.940 41.580 ;
        RECT 105.940 32.900 114.950 35.460 ;
        RECT 105.950 28.770 106.970 32.900 ;
        RECT 105.940 28.530 106.970 28.770 ;
        RECT 50.500 26.710 55.390 27.740 ;
        RECT 105.940 23.260 106.950 28.530 ;
        RECT 114.460 26.300 114.940 32.900 ;
        RECT 116.295 26.635 133.455 41.245 ;
        RECT 116.300 25.680 118.140 26.635 ;
        RECT 109.360 24.940 118.140 25.680 ;
        RECT 109.360 20.760 110.070 24.940 ;
        RECT 155.770 21.080 157.160 22.080 ;
        RECT 109.360 20.090 117.580 20.760 ;
        RECT 90.320 18.290 91.850 19.730 ;
        RECT 2.500 11.970 7.390 13.040 ;
        RECT 2.500 11.960 2.510 11.970 ;
        RECT 49.000 10.630 50.490 14.360 ;
        RECT 90.320 12.040 90.920 18.290 ;
        RECT 90.310 10.820 90.920 12.040 ;
        RECT 49.000 5.000 50.500 10.630 ;
        RECT 90.320 1.000 90.920 10.820 ;
        RECT 112.390 7.310 114.080 8.120 ;
        RECT 112.390 1.000 113.010 7.310 ;
        RECT 134.480 4.460 135.610 5.240 ;
        RECT 134.480 1.000 135.080 4.460 ;
        RECT 156.550 1.000 157.150 21.080 ;
        RECT 112.390 0.890 112.400 1.000 ;
        RECT 113.000 0.890 113.010 1.000 ;
        RECT 156.550 0.880 156.560 1.000 ;
  END
END tt_um_dsatizabal_opamp
END LIBRARY

