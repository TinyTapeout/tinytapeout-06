VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_mattvenn_r2r_dac
  CLASS BLOCK ;
  FOREIGN tt_um_mattvenn_r2r_dac ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met4 ;
        RECT 154.870 224.760 155.170 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 158.550 224.760 158.850 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 151.190 224.760 151.490 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 156.560 0.000 157.160 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 134.480 0.000 135.080 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 112.400 0.000 113.000 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 90.320 0.000 90.920 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 68.240 0.000 68.840 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 46.160 0.000 46.760 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 24.080 0.000 24.680 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 2.000 0.000 2.600 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 147.510 224.760 147.810 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 140.150 224.760 140.450 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 136.470 224.760 136.770 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 129.110 224.760 129.410 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 125.430 224.760 125.730 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met4 ;
        RECT 118.070 224.760 118.370 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met4 ;
        RECT 114.390 224.760 114.690 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.030 224.760 107.330 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 103.350 224.760 103.650 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 95.990 224.760 96.290 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 92.310 224.760 92.610 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 770.732971 ;
    ANTENNADIFFAREA 198.969498 ;
    PORT
      LAYER met4 ;
        RECT 29.750 224.760 30.050 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 770.732971 ;
    ANTENNADIFFAREA 198.969498 ;
    PORT
      LAYER met4 ;
        RECT 26.070 224.760 26.370 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 770.732971 ;
    ANTENNADIFFAREA 198.969498 ;
    PORT
      LAYER met4 ;
        RECT 22.390 224.760 22.690 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 770.732971 ;
    ANTENNADIFFAREA 198.969498 ;
    PORT
      LAYER met4 ;
        RECT 18.710 224.760 19.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 770.732971 ;
    ANTENNADIFFAREA 198.969498 ;
    PORT
      LAYER met4 ;
        RECT 15.030 224.760 15.330 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 770.732971 ;
    ANTENNADIFFAREA 198.969498 ;
    PORT
      LAYER met4 ;
        RECT 11.350 224.760 11.650 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 770.732971 ;
    ANTENNADIFFAREA 198.969498 ;
    PORT
      LAYER met4 ;
        RECT 7.670 224.760 7.970 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 770.732971 ;
    ANTENNADIFFAREA 198.969498 ;
    PORT
      LAYER met4 ;
        RECT 3.990 224.760 4.290 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 770.732971 ;
    ANTENNADIFFAREA 198.969498 ;
    PORT
      LAYER met4 ;
        RECT 59.190 224.760 59.490 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 770.732971 ;
    ANTENNADIFFAREA 198.969498 ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 770.732971 ;
    ANTENNADIFFAREA 198.969498 ;
    PORT
      LAYER met4 ;
        RECT 51.830 224.760 52.130 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 770.732971 ;
    ANTENNADIFFAREA 198.969498 ;
    PORT
      LAYER met4 ;
        RECT 48.150 224.760 48.450 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 770.732971 ;
    ANTENNADIFFAREA 198.969498 ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 770.732971 ;
    ANTENNADIFFAREA 198.969498 ;
    PORT
      LAYER met4 ;
        RECT 40.790 224.760 41.090 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 770.732971 ;
    ANTENNADIFFAREA 198.969498 ;
    PORT
      LAYER met4 ;
        RECT 37.110 224.760 37.410 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 770.732971 ;
    ANTENNADIFFAREA 198.969498 ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 770.732971 ;
    ANTENNADIFFAREA 198.969498 ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 770.732971 ;
    ANTENNADIFFAREA 198.969498 ;
    PORT
      LAYER met4 ;
        RECT 84.950 224.760 85.250 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 770.732971 ;
    ANTENNADIFFAREA 198.969498 ;
    PORT
      LAYER met4 ;
        RECT 81.270 224.760 81.570 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 770.732971 ;
    ANTENNADIFFAREA 198.969498 ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 770.732971 ;
    ANTENNADIFFAREA 198.969498 ;
    PORT
      LAYER met4 ;
        RECT 73.910 224.760 74.210 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 770.732971 ;
    ANTENNADIFFAREA 198.969498 ;
    PORT
      LAYER met4 ;
        RECT 70.230 224.760 70.530 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 770.732971 ;
    ANTENNADIFFAREA 198.969498 ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 770.732971 ;
    ANTENNADIFFAREA 198.969498 ;
    PORT
      LAYER met4 ;
        RECT 62.870 224.760 63.170 225.760 ;
    END
  END uo_out[7]
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 2.500 220.760 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 8.440 5.520 9.940 221.280 ;
    END
  END VGND
  OBS
      LAYER nwell ;
        RECT 18.090 204.925 92.530 206.530 ;
      LAYER pwell ;
        RECT 18.285 203.725 19.655 204.535 ;
        RECT 20.125 203.725 21.955 204.405 ;
        RECT 21.965 203.725 25.635 204.535 ;
        RECT 26.565 203.725 28.395 204.405 ;
        RECT 28.405 203.725 31.155 204.535 ;
        RECT 31.175 203.810 31.605 204.595 ;
        RECT 31.625 203.725 32.995 204.535 ;
        RECT 33.005 203.725 34.375 204.505 ;
        RECT 34.385 203.725 38.055 204.535 ;
        RECT 38.525 204.435 39.470 204.635 ;
        RECT 40.805 204.435 41.735 204.635 ;
        RECT 38.525 203.955 41.735 204.435 ;
        RECT 38.525 203.755 41.595 203.955 ;
        RECT 38.525 203.725 39.470 203.755 ;
        RECT 18.425 203.515 18.595 203.725 ;
        RECT 19.805 203.675 19.975 203.705 ;
        RECT 19.800 203.565 19.975 203.675 ;
        RECT 19.805 203.515 19.975 203.565 ;
        RECT 20.265 203.535 20.435 203.725 ;
        RECT 22.105 203.535 22.275 203.725 ;
        RECT 25.325 203.515 25.495 203.705 ;
        RECT 25.795 203.570 25.955 203.680 ;
        RECT 26.705 203.535 26.875 203.725 ;
        RECT 28.545 203.535 28.715 203.725 ;
        RECT 30.845 203.515 31.015 203.705 ;
        RECT 31.765 203.535 31.935 203.725 ;
        RECT 33.155 203.535 33.325 203.725 ;
        RECT 33.600 203.565 33.720 203.675 ;
        RECT 34.525 203.535 34.695 203.725 ;
        RECT 38.200 203.565 38.320 203.675 ;
        RECT 40.965 203.515 41.135 203.705 ;
        RECT 41.425 203.535 41.595 203.755 ;
        RECT 41.745 203.725 43.115 204.505 ;
        RECT 44.055 203.810 44.485 204.595 ;
        RECT 44.505 203.725 45.875 204.535 ;
        RECT 45.885 203.725 47.255 204.505 ;
        RECT 47.265 203.725 50.935 204.535 ;
        RECT 50.945 203.725 52.315 204.535 ;
        RECT 52.325 203.725 53.695 204.505 ;
        RECT 53.705 203.725 56.455 204.535 ;
        RECT 56.935 203.810 57.365 204.595 ;
        RECT 57.385 204.435 58.330 204.635 ;
        RECT 59.665 204.435 60.595 204.635 ;
        RECT 57.385 203.955 60.595 204.435 ;
        RECT 57.385 203.755 60.455 203.955 ;
        RECT 57.385 203.725 58.330 203.755 ;
        RECT 41.895 203.535 42.065 203.725 ;
        RECT 42.805 203.515 42.975 203.705 ;
        RECT 43.275 203.560 43.435 203.680 ;
        RECT 44.645 203.535 44.815 203.725 ;
        RECT 46.035 203.535 46.205 203.725 ;
        RECT 47.405 203.535 47.575 203.725 ;
        RECT 51.085 203.535 51.255 203.725 ;
        RECT 51.545 203.515 51.715 203.705 ;
        RECT 52.475 203.535 52.645 203.725 ;
        RECT 53.845 203.535 54.015 203.725 ;
        RECT 18.285 202.705 19.655 203.515 ;
        RECT 19.665 202.705 25.175 203.515 ;
        RECT 25.185 202.705 30.695 203.515 ;
        RECT 30.705 202.705 33.455 203.515 ;
        RECT 33.965 202.835 41.275 203.515 ;
        RECT 41.285 202.835 43.115 203.515 ;
        RECT 33.965 202.605 35.315 202.835 ;
        RECT 36.850 202.615 37.760 202.835 ;
        RECT 41.285 202.605 42.630 202.835 ;
        RECT 44.055 202.645 44.485 203.430 ;
        RECT 44.545 202.835 51.855 203.515 ;
        RECT 51.865 203.485 52.810 203.515 ;
        RECT 54.765 203.485 54.935 203.705 ;
        RECT 55.235 203.560 55.395 203.670 ;
        RECT 56.600 203.565 56.720 203.675 ;
        RECT 60.285 203.535 60.455 203.755 ;
        RECT 60.605 203.725 61.975 204.505 ;
        RECT 61.985 203.725 64.735 204.535 ;
        RECT 65.205 203.725 66.575 204.505 ;
        RECT 66.585 203.725 69.335 204.535 ;
        RECT 69.815 203.810 70.245 204.595 ;
        RECT 70.265 203.725 71.635 204.535 ;
        RECT 71.645 203.725 73.015 204.505 ;
        RECT 73.025 203.725 76.695 204.535 ;
        RECT 76.705 203.725 78.075 204.535 ;
        RECT 78.085 203.725 79.455 204.505 ;
        RECT 80.845 203.725 82.675 204.535 ;
        RECT 82.695 203.810 83.125 204.595 ;
        RECT 83.145 203.725 84.515 204.535 ;
        RECT 84.525 203.725 85.895 204.505 ;
        RECT 85.905 203.725 89.575 204.535 ;
        RECT 89.585 203.725 90.955 204.535 ;
        RECT 90.965 203.725 92.335 204.535 ;
        RECT 60.755 203.535 60.925 203.725 ;
        RECT 62.125 203.535 62.295 203.725 ;
        RECT 63.045 203.515 63.215 203.705 ;
        RECT 63.505 203.515 63.675 203.705 ;
        RECT 64.880 203.565 65.000 203.675 ;
        RECT 65.355 203.535 65.525 203.725 ;
        RECT 66.265 203.535 66.435 203.705 ;
        RECT 66.725 203.535 66.895 203.725 ;
        RECT 69.480 203.565 69.600 203.675 ;
        RECT 70.405 203.535 70.575 203.725 ;
        RECT 71.795 203.535 71.965 203.725 ;
        RECT 73.165 203.535 73.335 203.725 ;
        RECT 76.845 203.535 77.015 203.725 ;
        RECT 66.265 203.515 66.465 203.535 ;
        RECT 77.305 203.515 77.475 203.705 ;
        RECT 77.765 203.515 77.935 203.705 ;
        RECT 79.135 203.535 79.305 203.725 ;
        RECT 79.605 203.535 79.775 203.705 ;
        RECT 80.985 203.535 81.155 203.725 ;
        RECT 83.285 203.535 83.455 203.725 ;
        RECT 84.665 203.535 84.835 203.725 ;
        RECT 86.045 203.535 86.215 203.725 ;
        RECT 87.425 203.515 87.595 203.705 ;
        RECT 88.805 203.515 88.975 203.705 ;
        RECT 89.725 203.535 89.895 203.725 ;
        RECT 90.640 203.565 90.760 203.675 ;
        RECT 92.025 203.515 92.195 203.725 ;
        RECT 51.865 203.285 54.935 203.485 ;
        RECT 44.545 202.605 45.895 202.835 ;
        RECT 47.430 202.615 48.340 202.835 ;
        RECT 51.865 202.805 55.075 203.285 ;
        RECT 51.865 202.605 52.810 202.805 ;
        RECT 54.145 202.605 55.075 202.805 ;
        RECT 56.045 202.835 63.355 203.515 ;
        RECT 56.045 202.605 57.395 202.835 ;
        RECT 58.930 202.615 59.840 202.835 ;
        RECT 63.365 202.705 66.115 203.515 ;
        RECT 66.265 202.835 69.795 203.515 ;
        RECT 66.970 202.605 69.795 202.835 ;
        RECT 69.815 202.645 70.245 203.430 ;
        RECT 70.305 202.835 77.615 203.515 ;
        RECT 77.625 202.835 87.235 203.515 ;
        RECT 70.305 202.605 71.655 202.835 ;
        RECT 73.190 202.615 74.100 202.835 ;
        RECT 82.135 202.615 83.065 202.835 ;
        RECT 85.895 202.605 87.235 202.835 ;
        RECT 87.295 202.605 88.645 203.515 ;
        RECT 88.665 202.705 90.495 203.515 ;
        RECT 90.965 202.705 92.335 203.515 ;
      LAYER nwell ;
        RECT 18.090 199.485 92.530 202.315 ;
      LAYER pwell ;
        RECT 18.285 198.285 19.655 199.095 ;
        RECT 19.665 198.285 25.175 199.095 ;
        RECT 25.185 198.285 30.695 199.095 ;
        RECT 31.175 198.370 31.605 199.155 ;
        RECT 31.625 198.285 37.135 199.095 ;
        RECT 37.990 198.965 40.815 199.195 ;
        RECT 37.285 198.285 40.815 198.965 ;
        RECT 40.825 198.285 46.335 199.095 ;
        RECT 48.110 198.965 50.935 199.195 ;
        RECT 47.405 198.285 50.935 198.965 ;
        RECT 50.945 198.285 56.455 199.095 ;
        RECT 56.935 198.370 57.365 199.155 ;
        RECT 59.150 198.965 61.975 199.195 ;
        RECT 58.445 198.285 61.975 198.965 ;
        RECT 61.985 198.285 67.495 199.095 ;
        RECT 67.505 198.995 68.450 199.195 ;
        RECT 69.785 198.995 70.715 199.195 ;
        RECT 67.505 198.515 70.715 198.995 ;
        RECT 67.505 198.315 70.575 198.515 ;
        RECT 67.505 198.285 68.450 198.315 ;
        RECT 18.425 198.075 18.595 198.285 ;
        RECT 19.805 198.075 19.975 198.285 ;
        RECT 25.325 198.075 25.495 198.285 ;
        RECT 30.845 198.235 31.015 198.265 ;
        RECT 30.840 198.125 31.015 198.235 ;
        RECT 30.845 198.075 31.015 198.125 ;
        RECT 31.765 198.095 31.935 198.285 ;
        RECT 37.285 198.265 37.485 198.285 ;
        RECT 34.520 198.125 34.640 198.235 ;
        RECT 34.985 198.095 35.155 198.265 ;
        RECT 37.285 198.095 37.455 198.265 ;
        RECT 34.985 198.075 35.185 198.095 ;
        RECT 38.665 198.075 38.835 198.265 ;
        RECT 40.965 198.095 41.135 198.285 ;
        RECT 47.405 198.265 47.605 198.285 ;
        RECT 46.495 198.130 46.655 198.240 ;
        RECT 47.405 198.095 47.575 198.265 ;
        RECT 47.865 198.095 48.035 198.265 ;
        RECT 47.835 198.075 48.035 198.095 ;
        RECT 48.325 198.075 48.495 198.265 ;
        RECT 51.085 198.235 51.255 198.285 ;
        RECT 58.445 198.265 58.645 198.285 ;
        RECT 51.080 198.125 51.255 198.235 ;
        RECT 56.600 198.125 56.720 198.235 ;
        RECT 57.535 198.130 57.695 198.240 ;
        RECT 51.085 198.095 51.255 198.125 ;
        RECT 58.445 198.075 58.615 198.265 ;
        RECT 58.905 198.075 59.075 198.265 ;
        RECT 60.745 198.075 60.915 198.265 ;
        RECT 62.125 198.095 62.295 198.285 ;
        RECT 68.105 198.075 68.275 198.265 ;
        RECT 70.405 198.075 70.575 198.315 ;
        RECT 71.195 198.285 73.935 198.965 ;
        RECT 74.885 198.285 76.235 199.195 ;
        RECT 76.265 198.285 77.615 199.195 ;
        RECT 78.545 198.285 80.360 199.195 ;
        RECT 80.385 198.285 82.215 199.095 ;
        RECT 82.695 198.370 83.125 199.155 ;
        RECT 83.145 198.285 84.515 199.095 ;
        RECT 84.620 198.965 85.540 199.195 ;
        RECT 84.620 198.285 88.085 198.965 ;
        RECT 88.215 198.285 89.565 199.195 ;
        RECT 89.585 198.285 90.955 199.095 ;
        RECT 90.965 198.285 92.335 199.095 ;
        RECT 70.860 198.125 70.980 198.235 ;
        RECT 73.625 198.095 73.795 198.285 ;
        RECT 74.095 198.130 74.255 198.240 ;
        RECT 75.000 198.095 75.170 198.285 ;
        RECT 76.380 198.075 76.550 198.265 ;
        RECT 76.855 198.120 77.015 198.230 ;
        RECT 77.300 198.095 77.470 198.285 ;
        RECT 77.770 198.075 77.940 198.265 ;
        RECT 79.605 198.075 79.775 198.265 ;
        RECT 80.065 198.095 80.235 198.285 ;
        RECT 80.525 198.095 80.695 198.285 ;
        RECT 82.365 198.235 82.535 198.265 ;
        RECT 82.360 198.125 82.535 198.235 ;
        RECT 82.365 198.075 82.535 198.125 ;
        RECT 83.285 198.095 83.455 198.285 ;
        RECT 87.885 198.095 88.055 198.285 ;
        RECT 88.345 198.095 88.515 198.285 ;
        RECT 89.725 198.095 89.895 198.285 ;
        RECT 92.025 198.075 92.195 198.285 ;
        RECT 18.285 197.265 19.655 198.075 ;
        RECT 19.665 197.265 25.175 198.075 ;
        RECT 25.185 197.265 30.695 198.075 ;
        RECT 30.705 197.265 34.375 198.075 ;
        RECT 34.985 197.395 38.515 198.075 ;
        RECT 35.690 197.165 38.515 197.395 ;
        RECT 38.525 197.265 44.035 198.075 ;
        RECT 44.055 197.205 44.485 197.990 ;
        RECT 44.505 197.395 48.035 198.075 ;
        RECT 44.505 197.165 47.330 197.395 ;
        RECT 48.185 197.265 50.935 198.075 ;
        RECT 51.445 197.395 58.755 198.075 ;
        RECT 51.445 197.165 52.795 197.395 ;
        RECT 54.330 197.175 55.240 197.395 ;
        RECT 58.765 197.265 60.595 198.075 ;
        RECT 60.605 197.395 67.915 198.075 ;
        RECT 64.120 197.175 65.030 197.395 ;
        RECT 66.565 197.165 67.915 197.395 ;
        RECT 67.965 197.265 69.795 198.075 ;
        RECT 69.815 197.205 70.245 197.990 ;
        RECT 70.265 197.265 73.015 198.075 ;
        RECT 73.025 197.165 76.695 198.075 ;
        RECT 77.625 197.165 79.455 198.075 ;
        RECT 79.465 197.265 82.215 198.075 ;
        RECT 82.225 197.395 90.925 198.075 ;
        RECT 85.770 197.175 86.680 197.395 ;
        RECT 88.220 197.165 90.925 197.395 ;
        RECT 90.965 197.265 92.335 198.075 ;
      LAYER nwell ;
        RECT 18.090 194.045 92.530 196.875 ;
      LAYER pwell ;
        RECT 18.285 192.845 19.655 193.655 ;
        RECT 19.665 192.845 25.175 193.655 ;
        RECT 25.185 192.845 30.695 193.655 ;
        RECT 31.175 192.930 31.605 193.715 ;
        RECT 31.665 193.525 33.015 193.755 ;
        RECT 34.550 193.525 35.460 193.745 ;
        RECT 31.665 192.845 38.975 193.525 ;
        RECT 38.985 192.845 41.735 193.655 ;
        RECT 45.260 193.525 46.170 193.745 ;
        RECT 47.705 193.525 49.055 193.755 ;
        RECT 41.745 192.845 49.055 193.525 ;
        RECT 49.105 193.555 50.060 193.755 ;
        RECT 49.105 192.875 51.385 193.555 ;
        RECT 49.105 192.845 50.060 192.875 ;
        RECT 18.425 192.635 18.595 192.845 ;
        RECT 19.805 192.635 19.975 192.845 ;
        RECT 25.325 192.635 25.495 192.845 ;
        RECT 30.845 192.795 31.015 192.825 ;
        RECT 30.840 192.685 31.015 192.795 ;
        RECT 36.360 192.685 36.480 192.795 ;
        RECT 30.845 192.635 31.015 192.685 ;
        RECT 38.665 192.655 38.835 192.845 ;
        RECT 39.125 192.655 39.295 192.845 ;
        RECT 18.285 191.825 19.655 192.635 ;
        RECT 19.665 191.825 25.175 192.635 ;
        RECT 25.185 191.825 30.695 192.635 ;
        RECT 30.705 191.825 36.215 192.635 ;
        RECT 36.685 192.605 37.630 192.635 ;
        RECT 39.585 192.605 39.755 192.825 ;
        RECT 40.045 192.635 40.215 192.825 ;
        RECT 41.885 192.655 42.055 192.845 ;
        RECT 43.720 192.685 43.840 192.795 ;
        RECT 44.645 192.635 44.815 192.825 ;
        RECT 50.165 192.635 50.335 192.825 ;
        RECT 51.090 192.655 51.260 192.875 ;
        RECT 51.415 192.845 52.765 193.755 ;
        RECT 53.705 193.555 54.635 193.755 ;
        RECT 55.970 193.555 56.915 193.755 ;
        RECT 53.705 193.075 56.915 193.555 ;
        RECT 53.845 192.875 56.915 193.075 ;
        RECT 56.935 192.930 57.365 193.715 ;
        RECT 58.230 193.525 61.055 193.755 ;
        RECT 51.545 192.655 51.715 192.845 ;
        RECT 52.935 192.690 53.095 192.800 ;
        RECT 53.845 192.655 54.015 192.875 ;
        RECT 55.970 192.845 56.915 192.875 ;
        RECT 57.525 192.845 61.055 193.525 ;
        RECT 61.065 192.845 64.735 193.655 ;
        RECT 65.205 193.525 68.030 193.755 ;
        RECT 68.885 193.555 69.830 193.755 ;
        RECT 71.165 193.555 72.095 193.755 ;
        RECT 73.245 193.665 74.195 193.755 ;
        RECT 65.205 192.845 68.735 193.525 ;
        RECT 68.885 193.075 72.095 193.555 ;
        RECT 68.885 192.875 71.955 193.075 ;
        RECT 68.885 192.845 69.830 192.875 ;
        RECT 57.525 192.825 57.725 192.845 ;
        RECT 57.525 192.635 57.695 192.825 ;
        RECT 57.985 192.635 58.155 192.825 ;
        RECT 60.745 192.635 60.915 192.825 ;
        RECT 61.205 192.655 61.375 192.845 ;
        RECT 68.535 192.825 68.735 192.845 ;
        RECT 62.580 192.685 62.700 192.795 ;
        RECT 63.045 192.635 63.215 192.825 ;
        RECT 64.880 192.685 65.000 192.795 ;
        RECT 65.805 192.635 65.975 192.825 ;
        RECT 68.565 192.655 68.735 192.825 ;
        RECT 69.480 192.685 69.600 192.795 ;
        RECT 70.405 192.635 70.575 192.825 ;
        RECT 71.785 192.655 71.955 192.875 ;
        RECT 72.265 192.845 74.195 193.665 ;
        RECT 74.405 192.845 75.755 193.755 ;
        RECT 75.785 192.845 79.455 193.755 ;
        RECT 80.515 193.525 81.445 193.755 ;
        RECT 79.610 192.845 81.445 193.525 ;
        RECT 82.695 192.930 83.125 193.715 ;
        RECT 83.145 192.845 86.620 193.755 ;
        RECT 86.825 192.845 90.495 193.655 ;
        RECT 90.965 192.845 92.335 193.655 ;
        RECT 72.265 192.825 72.415 192.845 ;
        RECT 72.245 192.655 72.415 192.825 ;
        RECT 75.470 192.655 75.640 192.845 ;
        RECT 75.935 192.680 76.095 192.790 ;
        RECT 76.845 192.655 77.015 192.825 ;
        RECT 76.865 192.635 77.015 192.655 ;
        RECT 79.145 192.635 79.315 192.845 ;
        RECT 79.610 192.825 79.775 192.845 ;
        RECT 79.605 192.655 79.775 192.825 ;
        RECT 81.915 192.795 82.075 192.800 ;
        RECT 81.900 192.690 82.075 192.795 ;
        RECT 81.900 192.685 82.020 192.690 ;
        RECT 82.365 192.635 82.535 192.825 ;
        RECT 83.290 192.655 83.460 192.845 ;
        RECT 86.965 192.655 87.135 192.845 ;
        RECT 90.640 192.685 90.760 192.795 ;
        RECT 92.025 192.635 92.195 192.845 ;
        RECT 36.685 192.405 39.755 192.605 ;
        RECT 36.685 191.925 39.895 192.405 ;
        RECT 36.685 191.725 37.630 191.925 ;
        RECT 38.965 191.725 39.895 191.925 ;
        RECT 39.905 191.825 43.575 192.635 ;
        RECT 44.055 191.765 44.485 192.550 ;
        RECT 44.505 191.825 50.015 192.635 ;
        RECT 50.025 191.825 53.695 192.635 ;
        RECT 54.625 191.725 57.835 192.635 ;
        RECT 57.845 191.955 60.595 192.635 ;
        RECT 59.665 191.725 60.595 191.955 ;
        RECT 60.605 191.825 62.435 192.635 ;
        RECT 62.905 191.955 65.655 192.635 ;
        RECT 64.725 191.725 65.655 191.955 ;
        RECT 65.665 191.825 69.335 192.635 ;
        RECT 69.815 191.765 70.245 192.550 ;
        RECT 70.265 191.825 75.775 192.635 ;
        RECT 76.865 191.815 78.795 192.635 ;
        RECT 79.005 191.825 81.755 192.635 ;
        RECT 82.225 191.955 90.925 192.635 ;
        RECT 77.845 191.725 78.795 191.815 ;
        RECT 85.770 191.735 86.680 191.955 ;
        RECT 88.220 191.725 90.925 191.955 ;
        RECT 90.965 191.825 92.335 192.635 ;
      LAYER nwell ;
        RECT 18.090 188.605 92.530 191.435 ;
      LAYER pwell ;
        RECT 18.285 187.405 19.655 188.215 ;
        RECT 19.665 187.405 25.175 188.215 ;
        RECT 25.185 187.405 30.695 188.215 ;
        RECT 31.175 187.490 31.605 188.275 ;
        RECT 31.625 187.405 34.375 188.215 ;
        RECT 34.425 187.405 37.595 188.315 ;
        RECT 37.605 187.405 40.355 188.215 ;
        RECT 41.020 187.405 44.495 188.315 ;
        RECT 44.505 187.405 46.335 188.215 ;
        RECT 48.625 188.085 49.555 188.315 ;
        RECT 46.805 187.405 49.555 188.085 ;
        RECT 49.565 187.405 53.220 188.315 ;
        RECT 53.245 188.085 54.165 188.315 ;
        RECT 53.245 187.405 56.830 188.085 ;
        RECT 56.935 187.490 57.365 188.275 ;
        RECT 58.320 187.405 61.975 188.315 ;
        RECT 61.985 187.405 63.815 188.215 ;
        RECT 67.340 188.085 68.250 188.305 ;
        RECT 69.785 188.085 71.135 188.315 ;
        RECT 63.825 187.405 71.135 188.085 ;
        RECT 71.280 188.085 72.200 188.315 ;
        RECT 71.280 187.405 74.745 188.085 ;
        RECT 75.805 187.405 77.155 188.315 ;
        RECT 77.165 187.405 78.995 188.215 ;
        RECT 79.005 188.085 79.925 188.315 ;
        RECT 79.005 187.405 81.295 188.085 ;
        RECT 81.305 187.405 82.675 188.215 ;
        RECT 82.695 187.490 83.125 188.275 ;
        RECT 83.145 187.405 86.620 188.315 ;
        RECT 86.825 187.405 90.495 188.215 ;
        RECT 90.965 187.405 92.335 188.215 ;
        RECT 18.425 187.195 18.595 187.405 ;
        RECT 19.805 187.195 19.975 187.405 ;
        RECT 25.325 187.195 25.495 187.405 ;
        RECT 30.845 187.355 31.015 187.385 ;
        RECT 30.840 187.245 31.015 187.355 ;
        RECT 30.845 187.195 31.015 187.245 ;
        RECT 31.765 187.215 31.935 187.405 ;
        RECT 34.525 187.385 34.695 187.405 ;
        RECT 34.525 187.215 34.700 187.385 ;
        RECT 18.285 186.385 19.655 187.195 ;
        RECT 19.665 186.385 25.175 187.195 ;
        RECT 25.185 186.385 30.695 187.195 ;
        RECT 30.705 186.385 34.375 187.195 ;
        RECT 34.530 187.165 34.700 187.215 ;
        RECT 36.190 187.165 37.135 187.195 ;
        RECT 37.290 187.165 37.460 187.385 ;
        RECT 37.745 187.215 37.915 187.405 ;
        RECT 38.950 187.165 39.895 187.195 ;
        RECT 34.385 186.485 37.135 187.165 ;
        RECT 37.145 186.485 39.895 187.165 ;
        RECT 40.045 187.165 40.215 187.385 ;
        RECT 40.500 187.245 40.620 187.355 ;
        RECT 43.275 187.240 43.435 187.350 ;
        RECT 44.180 187.215 44.350 187.405 ;
        RECT 44.645 187.215 44.815 187.405 ;
        RECT 46.480 187.245 46.600 187.355 ;
        RECT 46.945 187.215 47.115 187.405 ;
        RECT 47.405 187.195 47.575 187.385 ;
        RECT 47.865 187.195 48.035 187.385 ;
        RECT 49.710 187.215 49.880 187.405 ;
        RECT 51.085 187.195 51.255 187.385 ;
        RECT 52.925 187.195 53.095 187.385 ;
        RECT 53.390 187.215 53.560 187.405 ;
        RECT 55.225 187.195 55.395 187.385 ;
        RECT 57.535 187.250 57.695 187.360 ;
        RECT 42.170 187.165 43.115 187.195 ;
        RECT 40.045 186.965 43.115 187.165 ;
        RECT 36.190 186.285 37.135 186.485 ;
        RECT 38.950 186.285 39.895 186.485 ;
        RECT 39.905 186.485 43.115 186.965 ;
        RECT 39.905 186.285 40.835 186.485 ;
        RECT 42.170 186.285 43.115 186.485 ;
        RECT 44.055 186.325 44.485 187.110 ;
        RECT 44.635 186.285 47.635 187.195 ;
        RECT 47.725 186.285 50.935 187.195 ;
        RECT 50.945 186.285 55.065 187.195 ;
        RECT 55.085 186.385 57.835 187.195 ;
        RECT 57.990 187.165 58.160 187.385 ;
        RECT 60.745 187.195 60.915 187.385 ;
        RECT 61.660 187.215 61.830 187.405 ;
        RECT 62.125 187.215 62.295 187.405 ;
        RECT 63.965 187.385 64.135 187.405 ;
        RECT 63.500 187.245 63.620 187.355 ;
        RECT 63.960 187.215 64.135 187.385 ;
        RECT 63.960 187.195 64.130 187.215 ;
        RECT 68.565 187.195 68.735 187.385 ;
        RECT 69.035 187.240 69.195 187.350 ;
        RECT 70.405 187.195 70.575 187.385 ;
        RECT 74.545 187.215 74.715 187.405 ;
        RECT 75.015 187.250 75.175 187.360 ;
        RECT 76.570 187.195 76.740 187.385 ;
        RECT 76.840 187.215 77.010 187.405 ;
        RECT 77.305 187.385 77.475 187.405 ;
        RECT 77.305 187.215 77.480 187.385 ;
        RECT 77.310 187.195 77.480 187.215 ;
        RECT 80.985 187.195 81.155 187.405 ;
        RECT 81.445 187.215 81.615 187.405 ;
        RECT 82.365 187.195 82.535 187.385 ;
        RECT 83.290 187.215 83.460 187.405 ;
        RECT 86.965 187.215 87.135 187.405 ;
        RECT 90.640 187.245 90.760 187.355 ;
        RECT 92.025 187.195 92.195 187.405 ;
        RECT 59.650 187.165 60.595 187.195 ;
        RECT 57.845 186.485 60.595 187.165 ;
        RECT 59.650 186.285 60.595 186.485 ;
        RECT 60.605 186.385 63.355 187.195 ;
        RECT 63.835 186.285 67.495 187.195 ;
        RECT 67.515 186.285 68.865 187.195 ;
        RECT 69.815 186.325 70.245 187.110 ;
        RECT 70.265 186.385 73.015 187.195 ;
        RECT 73.255 186.515 77.155 187.195 ;
        RECT 76.225 186.285 77.155 186.515 ;
        RECT 77.165 186.285 80.820 187.195 ;
        RECT 80.845 186.385 82.215 187.195 ;
        RECT 82.225 186.515 90.925 187.195 ;
        RECT 85.770 186.295 86.680 186.515 ;
        RECT 88.220 186.285 90.925 186.515 ;
        RECT 90.965 186.385 92.335 187.195 ;
      LAYER nwell ;
        RECT 18.090 183.165 92.530 185.995 ;
      LAYER pwell ;
        RECT 18.285 181.965 19.655 182.775 ;
        RECT 19.665 181.965 25.175 182.775 ;
        RECT 25.185 181.965 30.695 182.775 ;
        RECT 31.175 182.050 31.605 182.835 ;
        RECT 31.625 181.965 37.135 182.775 ;
        RECT 39.885 182.645 40.815 182.875 ;
        RECT 38.065 181.965 40.815 182.645 ;
        RECT 41.830 181.965 50.935 182.645 ;
        RECT 50.945 181.965 56.455 182.775 ;
        RECT 56.935 182.050 57.365 182.835 ;
        RECT 57.385 181.965 62.895 182.775 ;
        RECT 62.905 181.965 64.275 182.775 ;
        RECT 64.575 181.965 67.495 182.875 ;
        RECT 67.505 181.965 76.610 182.645 ;
        RECT 76.705 181.965 78.535 182.775 ;
        RECT 78.555 181.965 81.285 182.875 ;
        RECT 81.305 181.965 82.655 182.875 ;
        RECT 82.695 182.050 83.125 182.835 ;
        RECT 83.145 181.965 88.655 182.775 ;
        RECT 88.665 181.965 90.495 182.775 ;
        RECT 90.965 181.965 92.335 182.775 ;
        RECT 18.425 181.755 18.595 181.965 ;
        RECT 19.805 181.755 19.975 181.965 ;
        RECT 25.325 181.755 25.495 181.965 ;
        RECT 30.845 181.915 31.015 181.945 ;
        RECT 30.840 181.805 31.015 181.915 ;
        RECT 30.845 181.755 31.015 181.805 ;
        RECT 31.765 181.775 31.935 181.965 ;
        RECT 36.365 181.755 36.535 181.945 ;
        RECT 37.295 181.810 37.455 181.920 ;
        RECT 38.205 181.775 38.375 181.965 ;
        RECT 40.045 181.755 40.215 181.945 ;
        RECT 40.975 181.810 41.135 181.920 ;
        RECT 42.340 181.755 42.510 181.945 ;
        RECT 42.805 181.755 42.975 181.945 ;
        RECT 44.645 181.755 44.815 181.945 ;
        RECT 48.325 181.755 48.495 181.945 ;
        RECT 48.785 181.755 48.955 181.945 ;
        RECT 50.625 181.775 50.795 181.965 ;
        RECT 51.085 181.775 51.255 181.965 ;
        RECT 51.540 181.805 51.660 181.915 ;
        RECT 52.925 181.755 53.095 181.945 ;
        RECT 54.305 181.755 54.475 181.945 ;
        RECT 54.765 181.755 54.935 181.945 ;
        RECT 57.525 181.915 57.695 181.965 ;
        RECT 56.600 181.805 56.720 181.915 ;
        RECT 57.520 181.805 57.695 181.915 ;
        RECT 57.525 181.775 57.695 181.805 ;
        RECT 60.285 181.755 60.455 181.945 ;
        RECT 63.045 181.775 63.215 181.965 ;
        RECT 63.960 181.755 64.130 181.945 ;
        RECT 65.805 181.755 65.975 181.945 ;
        RECT 66.265 181.755 66.435 181.945 ;
        RECT 67.180 181.775 67.350 181.965 ;
        RECT 67.645 181.775 67.815 181.965 ;
        RECT 70.405 181.755 70.575 181.945 ;
        RECT 71.785 181.755 71.955 181.945 ;
        RECT 74.545 181.755 74.715 181.945 ;
        RECT 76.380 181.805 76.500 181.915 ;
        RECT 76.845 181.775 77.015 181.965 ;
        RECT 78.685 181.775 78.855 181.965 ;
        RECT 82.370 181.945 82.540 181.965 ;
        RECT 76.855 181.755 77.015 181.775 ;
        RECT 81.900 181.755 82.070 181.945 ;
        RECT 82.365 181.775 82.540 181.945 ;
        RECT 83.285 181.775 83.455 181.965 ;
        RECT 88.805 181.775 88.975 181.965 ;
        RECT 90.640 181.805 90.760 181.915 ;
        RECT 82.365 181.755 82.535 181.775 ;
        RECT 92.025 181.755 92.195 181.965 ;
        RECT 18.285 180.945 19.655 181.755 ;
        RECT 19.665 180.945 25.175 181.755 ;
        RECT 25.185 180.945 30.695 181.755 ;
        RECT 30.705 180.945 36.215 181.755 ;
        RECT 36.225 180.945 39.895 181.755 ;
        RECT 39.905 180.945 41.275 181.755 ;
        RECT 41.305 180.845 42.655 181.755 ;
        RECT 42.665 180.945 44.035 181.755 ;
        RECT 44.055 180.885 44.485 181.670 ;
        RECT 44.505 181.075 47.245 181.755 ;
        RECT 47.275 180.845 48.625 181.755 ;
        RECT 48.645 180.945 51.395 181.755 ;
        RECT 51.875 180.845 53.225 181.755 ;
        RECT 53.255 180.845 54.605 181.755 ;
        RECT 54.625 180.945 57.375 181.755 ;
        RECT 57.855 180.845 60.585 181.755 ;
        RECT 60.800 180.845 64.275 181.755 ;
        RECT 64.285 180.845 66.100 181.755 ;
        RECT 66.125 180.945 69.795 181.755 ;
        RECT 69.815 180.885 70.245 181.670 ;
        RECT 70.265 180.945 71.635 181.755 ;
        RECT 71.645 181.075 74.385 181.755 ;
        RECT 74.405 180.945 76.235 181.755 ;
        RECT 76.855 180.845 80.510 181.755 ;
        RECT 80.865 180.845 82.215 181.755 ;
        RECT 82.225 181.075 90.925 181.755 ;
        RECT 85.770 180.855 86.680 181.075 ;
        RECT 88.220 180.845 90.925 181.075 ;
        RECT 90.965 180.945 92.335 181.755 ;
      LAYER nwell ;
        RECT 18.090 177.725 92.530 180.555 ;
      LAYER pwell ;
        RECT 18.285 176.525 19.655 177.335 ;
        RECT 19.665 176.525 25.175 177.335 ;
        RECT 25.185 176.525 30.695 177.335 ;
        RECT 31.175 176.610 31.605 177.395 ;
        RECT 31.625 176.525 37.135 177.335 ;
        RECT 37.145 176.525 39.895 177.335 ;
        RECT 43.420 177.205 44.330 177.425 ;
        RECT 45.865 177.205 47.215 177.435 ;
        RECT 39.905 176.525 47.215 177.205 ;
        RECT 47.265 176.525 49.095 177.335 ;
        RECT 49.275 176.525 52.775 177.435 ;
        RECT 53.245 177.205 54.165 177.435 ;
        RECT 53.245 176.525 55.535 177.205 ;
        RECT 55.545 176.525 56.915 177.335 ;
        RECT 56.935 176.610 57.365 177.395 ;
        RECT 58.755 177.205 59.675 177.435 ;
        RECT 57.385 176.525 59.675 177.205 ;
        RECT 59.685 176.525 61.515 177.335 ;
        RECT 62.025 177.205 63.375 177.435 ;
        RECT 64.910 177.205 65.820 177.425 ;
        RECT 62.025 176.525 69.335 177.205 ;
        RECT 69.365 176.525 70.715 177.435 ;
        RECT 71.670 177.205 73.015 177.435 ;
        RECT 71.185 176.525 73.015 177.205 ;
        RECT 73.025 176.525 76.695 177.335 ;
        RECT 77.625 176.525 81.280 177.435 ;
        RECT 81.325 176.525 82.675 177.435 ;
        RECT 82.695 176.610 83.125 177.395 ;
        RECT 83.145 176.525 86.620 177.435 ;
        RECT 86.825 176.525 90.495 177.335 ;
        RECT 90.965 176.525 92.335 177.335 ;
        RECT 18.425 176.315 18.595 176.525 ;
        RECT 19.805 176.315 19.975 176.525 ;
        RECT 25.325 176.315 25.495 176.525 ;
        RECT 30.845 176.475 31.015 176.505 ;
        RECT 30.840 176.365 31.015 176.475 ;
        RECT 30.845 176.315 31.015 176.365 ;
        RECT 31.765 176.335 31.935 176.525 ;
        RECT 37.285 176.335 37.455 176.525 ;
        RECT 40.045 176.335 40.215 176.525 ;
        RECT 41.425 176.315 41.595 176.505 ;
        RECT 42.800 176.315 42.970 176.505 ;
        RECT 43.275 176.360 43.435 176.470 ;
        RECT 44.655 176.360 44.815 176.470 ;
        RECT 45.560 176.335 45.730 176.505 ;
        RECT 47.405 176.335 47.575 176.525 ;
        RECT 49.275 176.505 49.410 176.525 ;
        RECT 49.240 176.335 49.415 176.505 ;
        RECT 50.620 176.365 50.740 176.475 ;
        RECT 45.595 176.315 45.730 176.335 ;
        RECT 49.245 176.315 49.415 176.335 ;
        RECT 51.085 176.315 51.255 176.505 ;
        RECT 52.920 176.365 53.040 176.475 ;
        RECT 53.385 176.315 53.555 176.505 ;
        RECT 54.765 176.315 54.935 176.505 ;
        RECT 55.225 176.335 55.395 176.525 ;
        RECT 55.685 176.335 55.855 176.525 ;
        RECT 57.525 176.475 57.695 176.525 ;
        RECT 57.520 176.365 57.695 176.475 ;
        RECT 57.525 176.335 57.695 176.365 ;
        RECT 59.825 176.335 59.995 176.525 ;
        RECT 61.660 176.365 61.780 176.475 ;
        RECT 66.725 176.315 66.895 176.505 ;
        RECT 67.185 176.315 67.355 176.505 ;
        RECT 69.025 176.335 69.195 176.525 ;
        RECT 69.480 176.335 69.650 176.525 ;
        RECT 70.860 176.365 70.980 176.475 ;
        RECT 71.325 176.335 71.495 176.525 ;
        RECT 73.165 176.505 73.335 176.525 ;
        RECT 73.160 176.335 73.335 176.505 ;
        RECT 73.160 176.315 73.330 176.335 ;
        RECT 18.285 175.505 19.655 176.315 ;
        RECT 19.665 175.505 25.175 176.315 ;
        RECT 25.185 175.505 30.695 176.315 ;
        RECT 30.705 175.505 34.375 176.315 ;
        RECT 34.425 175.635 41.735 176.315 ;
        RECT 34.425 175.405 35.775 175.635 ;
        RECT 37.310 175.415 38.220 175.635 ;
        RECT 41.765 175.405 43.115 176.315 ;
        RECT 44.055 175.445 44.485 176.230 ;
        RECT 45.595 175.405 49.095 176.315 ;
        RECT 49.115 175.405 50.465 176.315 ;
        RECT 50.960 175.405 52.775 176.315 ;
        RECT 53.255 175.405 54.605 176.315 ;
        RECT 54.625 175.505 57.375 176.315 ;
        RECT 57.930 175.635 67.035 176.315 ;
        RECT 67.045 175.505 69.795 176.315 ;
        RECT 69.815 175.445 70.245 176.230 ;
        RECT 70.555 175.405 73.475 176.315 ;
        RECT 73.485 176.285 74.440 176.315 ;
        RECT 75.470 176.285 75.640 176.505 ;
        RECT 75.925 176.315 76.095 176.505 ;
        RECT 76.855 176.370 77.015 176.480 ;
        RECT 77.305 176.335 77.475 176.505 ;
        RECT 77.770 176.335 77.940 176.525 ;
        RECT 82.360 176.505 82.530 176.525 ;
        RECT 77.310 176.315 77.475 176.335 ;
        RECT 79.605 176.315 79.775 176.505 ;
        RECT 82.360 176.335 82.535 176.505 ;
        RECT 83.290 176.335 83.460 176.525 ;
        RECT 86.965 176.335 87.135 176.525 ;
        RECT 90.640 176.365 90.760 176.475 ;
        RECT 82.365 176.315 82.535 176.335 ;
        RECT 92.025 176.315 92.195 176.525 ;
        RECT 73.485 175.605 75.765 176.285 ;
        RECT 73.485 175.405 74.440 175.605 ;
        RECT 75.785 175.505 77.155 176.315 ;
        RECT 77.310 175.635 79.145 176.315 ;
        RECT 78.215 175.405 79.145 175.635 ;
        RECT 79.465 175.505 82.215 176.315 ;
        RECT 82.225 175.635 90.925 176.315 ;
        RECT 85.770 175.415 86.680 175.635 ;
        RECT 88.220 175.405 90.925 175.635 ;
        RECT 90.965 175.505 92.335 176.315 ;
      LAYER nwell ;
        RECT 18.090 172.285 92.530 175.115 ;
      LAYER pwell ;
        RECT 18.285 171.085 19.655 171.895 ;
        RECT 19.665 171.085 25.175 171.895 ;
        RECT 25.185 171.085 30.695 171.895 ;
        RECT 31.175 171.170 31.605 171.955 ;
        RECT 31.625 171.085 37.135 171.895 ;
        RECT 40.720 171.765 41.640 171.995 ;
        RECT 38.175 171.085 41.640 171.765 ;
        RECT 41.745 171.085 44.495 171.895 ;
        RECT 44.965 171.085 46.780 171.995 ;
        RECT 46.805 171.085 50.475 171.895 ;
        RECT 50.965 171.085 52.315 171.995 ;
        RECT 53.465 171.905 54.415 171.995 ;
        RECT 52.485 171.085 54.415 171.905 ;
        RECT 55.675 171.765 56.605 171.995 ;
        RECT 54.770 171.085 56.605 171.765 ;
        RECT 56.935 171.170 57.365 171.955 ;
        RECT 57.385 171.085 61.055 171.995 ;
        RECT 61.085 171.085 62.435 171.995 ;
        RECT 62.485 171.765 63.835 171.995 ;
        RECT 65.370 171.765 66.280 171.985 ;
        RECT 62.485 171.085 69.795 171.765 ;
        RECT 69.805 171.085 72.555 171.895 ;
        RECT 73.025 171.085 74.840 171.995 ;
        RECT 75.325 171.765 76.245 171.995 ;
        RECT 75.325 171.085 77.615 171.765 ;
        RECT 77.625 171.085 78.995 171.895 ;
        RECT 81.080 171.765 82.215 171.995 ;
        RECT 79.005 171.085 82.215 171.765 ;
        RECT 82.695 171.170 83.125 171.955 ;
        RECT 83.225 171.085 86.675 171.995 ;
        RECT 87.380 171.765 88.300 171.995 ;
        RECT 87.380 171.085 90.845 171.765 ;
        RECT 90.965 171.085 92.335 171.895 ;
        RECT 18.425 170.875 18.595 171.085 ;
        RECT 19.805 170.875 19.975 171.085 ;
        RECT 25.325 170.875 25.495 171.085 ;
        RECT 30.845 171.035 31.015 171.065 ;
        RECT 30.840 170.925 31.015 171.035 ;
        RECT 30.845 170.875 31.015 170.925 ;
        RECT 31.765 170.895 31.935 171.085 ;
        RECT 32.680 170.925 32.800 171.035 ;
        RECT 37.295 170.930 37.455 171.040 ;
        RECT 38.205 170.895 38.375 171.085 ;
        RECT 40.045 170.875 40.215 171.065 ;
        RECT 40.505 170.875 40.675 171.065 ;
        RECT 41.885 170.895 42.055 171.085 ;
        RECT 42.340 170.875 42.510 171.065 ;
        RECT 43.720 170.925 43.840 171.035 ;
        RECT 44.635 170.875 44.805 171.065 ;
        RECT 46.485 170.895 46.655 171.085 ;
        RECT 46.945 170.895 47.115 171.085 ;
        RECT 47.870 170.875 48.040 171.065 ;
        RECT 49.245 170.875 49.415 171.065 ;
        RECT 50.620 170.925 50.740 171.035 ;
        RECT 51.080 170.895 51.250 171.085 ;
        RECT 52.485 171.065 52.635 171.085 ;
        RECT 54.770 171.065 54.935 171.085 ;
        RECT 60.740 171.065 60.910 171.085 ;
        RECT 52.465 170.875 52.635 171.065 ;
        RECT 54.765 170.895 54.935 171.065 ;
        RECT 57.985 170.875 58.155 171.065 ;
        RECT 60.740 170.895 60.915 171.065 ;
        RECT 61.200 170.895 61.370 171.085 ;
        RECT 60.765 170.875 60.915 170.895 ;
        RECT 63.045 170.875 63.215 171.065 ;
        RECT 64.425 170.875 64.595 171.065 ;
        RECT 69.485 170.895 69.655 171.085 ;
        RECT 69.945 170.895 70.115 171.085 ;
        RECT 70.405 170.875 70.575 171.065 ;
        RECT 72.705 171.035 72.875 171.065 ;
        RECT 72.240 170.925 72.360 171.035 ;
        RECT 72.700 170.925 72.875 171.035 ;
        RECT 72.705 170.875 72.875 170.925 ;
        RECT 74.545 170.895 74.715 171.085 ;
        RECT 75.000 170.925 75.120 171.035 ;
        RECT 75.930 170.875 76.100 171.065 ;
        RECT 77.305 170.875 77.475 171.085 ;
        RECT 77.765 170.895 77.935 171.085 ;
        RECT 79.145 170.895 79.315 171.085 ;
        RECT 80.985 170.875 81.155 171.065 ;
        RECT 82.365 171.035 82.535 171.065 ;
        RECT 82.360 170.925 82.535 171.035 ;
        RECT 82.365 170.875 82.535 170.925 ;
        RECT 83.285 170.895 83.455 171.085 ;
        RECT 86.960 170.925 87.080 171.035 ;
        RECT 90.645 170.895 90.815 171.085 ;
        RECT 92.025 170.875 92.195 171.085 ;
        RECT 18.285 170.065 19.655 170.875 ;
        RECT 19.665 170.065 25.175 170.875 ;
        RECT 25.185 170.065 30.695 170.875 ;
        RECT 30.705 170.065 32.535 170.875 ;
        RECT 33.045 170.195 40.355 170.875 ;
        RECT 33.045 169.965 34.395 170.195 ;
        RECT 35.930 169.975 36.840 170.195 ;
        RECT 40.380 169.965 42.195 170.875 ;
        RECT 42.225 169.965 43.575 170.875 ;
        RECT 44.055 170.005 44.485 170.790 ;
        RECT 44.505 169.965 47.715 170.875 ;
        RECT 47.725 169.965 49.075 170.875 ;
        RECT 49.105 170.195 52.315 170.875 ;
        RECT 51.180 169.965 52.315 170.195 ;
        RECT 52.325 170.065 57.835 170.875 ;
        RECT 57.845 170.065 60.595 170.875 ;
        RECT 60.765 170.055 62.695 170.875 ;
        RECT 62.905 170.095 64.275 170.875 ;
        RECT 64.285 170.065 69.795 170.875 ;
        RECT 61.745 169.965 62.695 170.055 ;
        RECT 69.815 170.005 70.245 170.790 ;
        RECT 70.265 170.065 72.095 170.875 ;
        RECT 72.565 169.965 75.775 170.875 ;
        RECT 75.785 169.965 77.135 170.875 ;
        RECT 77.165 170.065 80.835 170.875 ;
        RECT 80.845 170.065 82.215 170.875 ;
        RECT 82.225 170.195 90.925 170.875 ;
        RECT 85.770 169.975 86.680 170.195 ;
        RECT 88.220 169.965 90.925 170.195 ;
        RECT 90.965 170.065 92.335 170.875 ;
      LAYER nwell ;
        RECT 18.090 166.845 92.530 169.675 ;
      LAYER pwell ;
        RECT 18.285 165.645 19.655 166.455 ;
        RECT 19.665 165.645 25.175 166.455 ;
        RECT 25.185 165.645 30.695 166.455 ;
        RECT 31.175 165.730 31.605 166.515 ;
        RECT 54.385 166.465 55.335 166.555 ;
        RECT 31.625 165.645 37.135 166.455 ;
        RECT 37.145 165.645 42.655 166.455 ;
        RECT 42.665 165.645 48.175 166.455 ;
        RECT 48.185 165.645 51.855 166.455 ;
        RECT 51.865 165.645 53.235 166.455 ;
        RECT 53.405 165.645 55.335 166.465 ;
        RECT 55.545 165.645 56.915 166.455 ;
        RECT 56.935 165.730 57.365 166.515 ;
        RECT 57.385 165.645 61.055 166.555 ;
        RECT 61.065 165.645 63.805 166.325 ;
        RECT 63.825 165.645 69.335 166.455 ;
        RECT 69.345 165.645 72.095 166.455 ;
        RECT 72.200 166.325 73.120 166.555 ;
        RECT 72.200 165.645 75.665 166.325 ;
        RECT 76.245 165.645 78.060 166.555 ;
        RECT 78.085 165.645 79.435 166.555 ;
        RECT 79.465 165.645 82.215 166.455 ;
        RECT 82.695 165.730 83.125 166.515 ;
        RECT 83.145 165.645 88.655 166.455 ;
        RECT 88.665 165.645 90.495 166.455 ;
        RECT 90.965 165.645 92.335 166.455 ;
        RECT 18.425 165.435 18.595 165.645 ;
        RECT 19.805 165.435 19.975 165.645 ;
        RECT 25.325 165.435 25.495 165.645 ;
        RECT 30.845 165.595 31.015 165.625 ;
        RECT 30.840 165.485 31.015 165.595 ;
        RECT 30.845 165.435 31.015 165.485 ;
        RECT 31.765 165.455 31.935 165.645 ;
        RECT 36.365 165.435 36.535 165.625 ;
        RECT 37.285 165.455 37.455 165.645 ;
        RECT 38.200 165.485 38.320 165.595 ;
        RECT 38.670 165.435 38.840 165.625 ;
        RECT 40.045 165.435 40.215 165.625 ;
        RECT 42.805 165.455 42.975 165.645 ;
        RECT 43.720 165.485 43.840 165.595 ;
        RECT 44.640 165.455 44.810 165.625 ;
        RECT 48.325 165.455 48.495 165.645 ;
        RECT 44.675 165.435 44.810 165.455 ;
        RECT 50.165 165.435 50.335 165.625 ;
        RECT 52.005 165.455 52.175 165.645 ;
        RECT 53.405 165.625 53.555 165.645 ;
        RECT 52.465 165.455 52.635 165.625 ;
        RECT 53.385 165.455 53.555 165.625 ;
        RECT 52.465 165.435 52.615 165.455 ;
        RECT 53.850 165.435 54.020 165.625 ;
        RECT 54.305 165.455 54.475 165.625 ;
        RECT 55.685 165.455 55.855 165.645 ;
        RECT 56.605 165.455 56.775 165.625 ;
        RECT 57.530 165.455 57.700 165.645 ;
        RECT 61.205 165.455 61.375 165.645 ;
        RECT 63.965 165.455 64.135 165.645 ;
        RECT 54.310 165.435 54.475 165.455 ;
        RECT 56.625 165.435 56.775 165.455 ;
        RECT 65.805 165.435 65.975 165.625 ;
        RECT 66.275 165.480 66.435 165.590 ;
        RECT 69.485 165.435 69.655 165.645 ;
        RECT 70.405 165.435 70.575 165.625 ;
        RECT 75.465 165.455 75.635 165.645 ;
        RECT 75.920 165.485 76.040 165.595 ;
        RECT 77.765 165.455 77.935 165.645 ;
        RECT 78.230 165.455 78.400 165.645 ;
        RECT 79.140 165.435 79.310 165.625 ;
        RECT 79.605 165.455 79.775 165.645 ;
        RECT 80.530 165.435 80.700 165.625 ;
        RECT 82.365 165.595 82.535 165.625 ;
        RECT 82.360 165.485 82.535 165.595 ;
        RECT 82.365 165.435 82.535 165.485 ;
        RECT 83.285 165.455 83.455 165.645 ;
        RECT 88.805 165.455 88.975 165.645 ;
        RECT 90.640 165.485 90.760 165.595 ;
        RECT 92.025 165.435 92.195 165.645 ;
        RECT 18.285 164.625 19.655 165.435 ;
        RECT 19.665 164.625 25.175 165.435 ;
        RECT 25.185 164.625 30.695 165.435 ;
        RECT 30.705 164.625 36.215 165.435 ;
        RECT 36.225 164.625 38.055 165.435 ;
        RECT 38.525 164.525 39.875 165.435 ;
        RECT 39.905 164.625 43.575 165.435 ;
        RECT 44.055 164.565 44.485 165.350 ;
        RECT 44.675 164.525 48.175 165.435 ;
        RECT 48.185 164.755 50.475 165.435 ;
        RECT 48.185 164.525 49.105 164.755 ;
        RECT 50.685 164.615 52.615 165.435 ;
        RECT 50.685 164.525 51.635 164.615 ;
        RECT 52.785 164.525 54.135 165.435 ;
        RECT 54.310 164.755 56.145 165.435 ;
        RECT 55.215 164.525 56.145 164.755 ;
        RECT 56.625 164.615 58.555 165.435 ;
        RECT 57.605 164.525 58.555 164.615 ;
        RECT 58.805 164.755 66.115 165.435 ;
        RECT 58.805 164.525 60.155 164.755 ;
        RECT 61.690 164.535 62.600 164.755 ;
        RECT 67.045 164.525 69.795 165.435 ;
        RECT 69.815 164.565 70.245 165.350 ;
        RECT 70.265 164.755 77.575 165.435 ;
        RECT 73.780 164.535 74.690 164.755 ;
        RECT 76.225 164.525 77.575 164.755 ;
        RECT 77.625 164.525 79.455 165.435 ;
        RECT 80.385 164.525 82.215 165.435 ;
        RECT 82.225 164.755 90.925 165.435 ;
        RECT 85.770 164.535 86.680 164.755 ;
        RECT 88.220 164.525 90.925 164.755 ;
        RECT 90.965 164.625 92.335 165.435 ;
      LAYER nwell ;
        RECT 18.090 161.405 92.530 164.235 ;
      LAYER pwell ;
        RECT 18.285 160.205 19.655 161.015 ;
        RECT 19.665 160.205 25.175 161.015 ;
        RECT 25.185 160.205 30.695 161.015 ;
        RECT 31.175 160.290 31.605 161.075 ;
        RECT 31.625 160.205 35.295 161.015 ;
        RECT 39.740 160.885 40.650 161.105 ;
        RECT 42.185 160.885 43.535 161.115 ;
        RECT 36.225 160.205 43.535 160.885 ;
        RECT 43.585 160.205 46.335 161.015 ;
        RECT 46.815 160.205 48.165 161.115 ;
        RECT 48.185 160.205 50.935 161.015 ;
        RECT 51.405 160.885 52.325 161.115 ;
        RECT 51.405 160.205 53.695 160.885 ;
        RECT 53.705 160.205 55.055 161.115 ;
        RECT 55.085 160.205 56.915 161.015 ;
        RECT 56.935 160.290 57.365 161.075 ;
        RECT 57.385 160.205 60.125 160.885 ;
        RECT 60.145 160.205 61.515 160.985 ;
        RECT 61.525 160.205 67.035 161.015 ;
        RECT 67.045 160.205 68.415 161.015 ;
        RECT 68.440 160.205 70.255 161.115 ;
        RECT 70.265 160.205 75.775 161.015 ;
        RECT 76.265 160.205 77.615 161.115 ;
        RECT 77.625 160.205 79.440 161.115 ;
        RECT 79.465 160.205 82.215 161.015 ;
        RECT 82.695 160.290 83.125 161.075 ;
        RECT 83.160 160.205 84.975 161.115 ;
        RECT 84.985 160.205 90.495 161.015 ;
        RECT 90.965 160.205 92.335 161.015 ;
        RECT 18.425 159.995 18.595 160.205 ;
        RECT 19.805 159.995 19.975 160.205 ;
        RECT 25.325 159.995 25.495 160.205 ;
        RECT 30.845 160.155 31.015 160.185 ;
        RECT 30.840 160.045 31.015 160.155 ;
        RECT 30.845 159.995 31.015 160.045 ;
        RECT 31.765 160.015 31.935 160.205 ;
        RECT 35.455 160.050 35.615 160.160 ;
        RECT 36.365 160.155 36.535 160.205 ;
        RECT 36.360 160.045 36.535 160.155 ;
        RECT 36.365 160.015 36.535 160.045 ;
        RECT 36.825 159.995 36.995 160.185 ;
        RECT 43.725 160.015 43.895 160.205 ;
        RECT 46.480 160.045 46.600 160.155 ;
        RECT 46.945 160.015 47.115 160.205 ;
        RECT 48.325 160.015 48.495 160.205 ;
        RECT 51.080 160.045 51.200 160.155 ;
        RECT 53.385 159.995 53.555 160.205 ;
        RECT 53.850 160.015 54.020 160.205 ;
        RECT 54.765 159.995 54.935 160.185 ;
        RECT 55.225 160.015 55.395 160.205 ;
        RECT 56.605 159.995 56.775 160.185 ;
        RECT 57.525 160.015 57.695 160.205 ;
        RECT 60.285 160.015 60.455 160.205 ;
        RECT 61.665 160.015 61.835 160.205 ;
        RECT 62.125 159.995 62.295 160.185 ;
        RECT 67.185 160.015 67.355 160.205 ;
        RECT 67.645 159.995 67.815 160.185 ;
        RECT 68.565 160.015 68.735 160.205 ;
        RECT 69.480 160.045 69.600 160.155 ;
        RECT 70.405 159.995 70.575 160.205 ;
        RECT 75.920 160.045 76.040 160.155 ;
        RECT 76.380 160.015 76.550 160.205 ;
        RECT 79.145 160.015 79.315 160.205 ;
        RECT 79.605 159.995 79.775 160.205 ;
        RECT 82.360 160.045 82.480 160.155 ;
        RECT 83.285 160.015 83.455 160.205 ;
        RECT 85.125 160.015 85.295 160.205 ;
        RECT 88.345 159.995 88.515 160.185 ;
        RECT 90.640 160.045 90.760 160.155 ;
        RECT 92.025 159.995 92.195 160.205 ;
        RECT 18.285 159.185 19.655 159.995 ;
        RECT 19.665 159.185 25.175 159.995 ;
        RECT 25.185 159.185 30.695 159.995 ;
        RECT 30.705 159.185 36.215 159.995 ;
        RECT 36.685 159.315 43.995 159.995 ;
        RECT 40.200 159.095 41.110 159.315 ;
        RECT 42.645 159.085 43.995 159.315 ;
        RECT 44.055 159.125 44.485 159.910 ;
        RECT 44.590 159.315 53.695 159.995 ;
        RECT 54.625 159.315 56.455 159.995 ;
        RECT 55.110 159.085 56.455 159.315 ;
        RECT 56.465 159.185 61.975 159.995 ;
        RECT 61.985 159.185 67.495 159.995 ;
        RECT 67.505 159.185 69.335 159.995 ;
        RECT 69.815 159.125 70.245 159.910 ;
        RECT 70.265 159.315 79.370 159.995 ;
        RECT 79.465 159.315 88.165 159.995 ;
        RECT 83.010 159.095 83.920 159.315 ;
        RECT 85.460 159.085 88.165 159.315 ;
        RECT 88.205 159.185 90.955 159.995 ;
        RECT 90.965 159.185 92.335 159.995 ;
      LAYER nwell ;
        RECT 18.090 155.965 92.530 158.795 ;
      LAYER pwell ;
        RECT 18.285 154.765 19.655 155.575 ;
        RECT 19.665 154.765 25.175 155.575 ;
        RECT 25.185 154.765 30.695 155.575 ;
        RECT 31.175 154.850 31.605 155.635 ;
        RECT 31.625 154.765 37.135 155.575 ;
        RECT 37.145 154.765 42.655 155.575 ;
        RECT 42.665 154.765 44.495 155.575 ;
        RECT 44.525 154.765 45.875 155.675 ;
        RECT 45.895 154.765 47.245 155.675 ;
        RECT 47.360 155.445 48.280 155.675 ;
        RECT 53.940 155.445 55.075 155.675 ;
        RECT 47.360 154.765 50.825 155.445 ;
        RECT 51.865 154.765 55.075 155.445 ;
        RECT 55.085 154.765 56.915 155.575 ;
        RECT 56.935 154.850 57.365 155.635 ;
        RECT 57.405 154.765 58.755 155.675 ;
        RECT 62.280 155.445 63.190 155.665 ;
        RECT 64.725 155.445 66.075 155.675 ;
        RECT 58.765 154.765 66.075 155.445 ;
        RECT 66.295 154.765 69.795 155.675 ;
        RECT 72.460 155.445 73.380 155.675 ;
        RECT 69.915 154.765 73.380 155.445 ;
        RECT 73.655 154.765 77.155 155.675 ;
        RECT 79.820 155.445 80.740 155.675 ;
        RECT 77.275 154.765 80.740 155.445 ;
        RECT 80.845 154.765 82.660 155.675 ;
        RECT 82.695 154.850 83.125 155.635 ;
        RECT 83.155 154.765 84.505 155.675 ;
        RECT 84.525 154.765 90.035 155.575 ;
        RECT 90.965 154.765 92.335 155.575 ;
        RECT 18.425 154.555 18.595 154.765 ;
        RECT 19.805 154.555 19.975 154.765 ;
        RECT 25.325 154.555 25.495 154.765 ;
        RECT 30.845 154.715 31.015 154.745 ;
        RECT 30.840 154.605 31.015 154.715 ;
        RECT 30.845 154.555 31.015 154.605 ;
        RECT 31.765 154.575 31.935 154.765 ;
        RECT 36.365 154.555 36.535 154.745 ;
        RECT 37.285 154.575 37.455 154.765 ;
        RECT 41.885 154.555 42.055 154.745 ;
        RECT 42.805 154.575 42.975 154.765 ;
        RECT 43.720 154.605 43.840 154.715 ;
        RECT 44.645 154.555 44.815 154.745 ;
        RECT 45.560 154.575 45.730 154.765 ;
        RECT 46.480 154.575 46.650 154.745 ;
        RECT 46.945 154.575 47.115 154.765 ;
        RECT 50.625 154.575 50.795 154.765 ;
        RECT 51.095 154.610 51.255 154.720 ;
        RECT 52.005 154.575 52.175 154.765 ;
        RECT 46.515 154.555 46.650 154.575 ;
        RECT 18.285 153.745 19.655 154.555 ;
        RECT 19.665 153.745 25.175 154.555 ;
        RECT 25.185 153.745 30.695 154.555 ;
        RECT 30.705 153.745 36.215 154.555 ;
        RECT 36.225 153.745 41.735 154.555 ;
        RECT 41.760 153.645 43.575 154.555 ;
        RECT 44.055 153.685 44.485 154.470 ;
        RECT 44.505 153.745 46.335 154.555 ;
        RECT 46.515 153.645 50.015 154.555 ;
        RECT 50.025 154.525 50.970 154.555 ;
        RECT 52.925 154.525 53.095 154.745 ;
        RECT 55.225 154.575 55.395 154.765 ;
        RECT 58.440 154.745 58.610 154.765 ;
        RECT 56.145 154.555 56.315 154.745 ;
        RECT 58.440 154.575 58.615 154.745 ;
        RECT 58.445 154.555 58.595 154.575 ;
        RECT 58.905 154.555 59.075 154.765 ;
        RECT 66.295 154.745 66.430 154.765 ;
        RECT 64.425 154.555 64.595 154.745 ;
        RECT 66.260 154.575 66.430 154.745 ;
        RECT 67.180 154.555 67.350 154.745 ;
        RECT 69.485 154.555 69.655 154.745 ;
        RECT 69.945 154.575 70.115 154.765 ;
        RECT 73.655 154.745 73.790 154.765 ;
        RECT 70.410 154.555 70.580 154.745 ;
        RECT 73.620 154.575 73.790 154.745 ;
        RECT 74.085 154.555 74.255 154.745 ;
        RECT 75.465 154.555 75.635 154.745 ;
        RECT 77.305 154.575 77.475 154.765 ;
        RECT 82.365 154.575 82.535 154.765 ;
        RECT 82.825 154.555 82.995 154.745 ;
        RECT 83.285 154.575 83.455 154.765 ;
        RECT 84.665 154.575 84.835 154.765 ;
        RECT 88.345 154.555 88.515 154.745 ;
        RECT 90.195 154.610 90.355 154.720 ;
        RECT 92.025 154.555 92.195 154.765 ;
        RECT 50.025 154.325 53.095 154.525 ;
        RECT 50.025 153.845 53.235 154.325 ;
        RECT 50.025 153.645 50.970 153.845 ;
        RECT 52.305 153.645 53.235 153.845 ;
        RECT 53.245 153.875 56.455 154.555 ;
        RECT 53.245 153.645 54.380 153.875 ;
        RECT 56.665 153.735 58.595 154.555 ;
        RECT 58.765 153.745 64.275 154.555 ;
        RECT 64.285 153.745 66.115 154.555 ;
        RECT 56.665 153.645 57.615 153.735 ;
        RECT 66.145 153.645 67.495 154.555 ;
        RECT 67.505 153.875 69.795 154.555 ;
        RECT 67.505 153.645 68.425 153.875 ;
        RECT 69.815 153.685 70.245 154.470 ;
        RECT 70.265 153.875 73.935 154.555 ;
        RECT 72.345 153.645 73.935 153.875 ;
        RECT 73.955 153.645 75.305 154.555 ;
        RECT 75.325 153.875 82.635 154.555 ;
        RECT 78.840 153.655 79.750 153.875 ;
        RECT 81.285 153.645 82.635 153.875 ;
        RECT 82.685 153.745 88.195 154.555 ;
        RECT 88.205 153.745 90.955 154.555 ;
        RECT 90.965 153.745 92.335 154.555 ;
      LAYER nwell ;
        RECT 18.090 150.525 92.530 153.355 ;
      LAYER pwell ;
        RECT 18.285 149.325 19.655 150.135 ;
        RECT 19.665 149.325 25.175 150.135 ;
        RECT 25.185 149.325 30.695 150.135 ;
        RECT 31.175 149.410 31.605 150.195 ;
        RECT 31.625 149.325 35.295 150.135 ;
        RECT 35.305 149.325 36.675 150.135 ;
        RECT 40.200 150.005 41.110 150.225 ;
        RECT 42.645 150.005 43.995 150.235 ;
        RECT 47.160 150.005 48.080 150.235 ;
        RECT 36.685 149.325 43.995 150.005 ;
        RECT 44.615 149.325 48.080 150.005 ;
        RECT 48.205 149.325 49.555 150.235 ;
        RECT 50.025 149.325 52.945 150.235 ;
        RECT 53.245 149.325 56.915 150.135 ;
        RECT 56.935 149.410 57.365 150.195 ;
        RECT 57.385 149.325 60.135 150.135 ;
        RECT 60.160 149.325 61.975 150.235 ;
        RECT 62.005 149.325 63.355 150.235 ;
        RECT 63.365 149.325 68.875 150.135 ;
        RECT 69.445 149.325 72.555 150.235 ;
        RECT 72.565 149.325 73.935 150.135 ;
        RECT 73.945 149.325 75.295 150.235 ;
        RECT 75.325 149.325 80.835 150.135 ;
        RECT 80.845 149.325 82.675 150.135 ;
        RECT 82.695 149.410 83.125 150.195 ;
        RECT 83.145 149.325 88.655 150.135 ;
        RECT 88.665 149.325 90.495 150.135 ;
        RECT 90.965 149.325 92.335 150.135 ;
        RECT 18.425 149.115 18.595 149.325 ;
        RECT 19.805 149.115 19.975 149.325 ;
        RECT 25.325 149.115 25.495 149.325 ;
        RECT 30.845 149.275 31.015 149.305 ;
        RECT 30.840 149.165 31.015 149.275 ;
        RECT 30.845 149.115 31.015 149.165 ;
        RECT 31.765 149.135 31.935 149.325 ;
        RECT 35.445 149.135 35.615 149.325 ;
        RECT 36.365 149.115 36.535 149.305 ;
        RECT 36.825 149.135 36.995 149.325 ;
        RECT 41.885 149.115 42.055 149.305 ;
        RECT 43.720 149.165 43.840 149.275 ;
        RECT 44.180 149.165 44.300 149.275 ;
        RECT 44.645 149.115 44.815 149.325 ;
        RECT 48.320 149.135 48.490 149.325 ;
        RECT 50.170 149.305 50.340 149.325 ;
        RECT 49.700 149.165 49.820 149.275 ;
        RECT 50.165 149.135 50.340 149.305 ;
        RECT 53.385 149.135 53.555 149.325 ;
        RECT 50.165 149.115 50.335 149.135 ;
        RECT 53.840 149.115 54.010 149.305 ;
        RECT 55.220 149.165 55.340 149.275 ;
        RECT 56.610 149.115 56.780 149.305 ;
        RECT 57.525 149.135 57.695 149.325 ;
        RECT 60.285 149.115 60.455 149.325 ;
        RECT 18.285 148.305 19.655 149.115 ;
        RECT 19.665 148.305 25.175 149.115 ;
        RECT 25.185 148.305 30.695 149.115 ;
        RECT 30.705 148.305 36.215 149.115 ;
        RECT 36.225 148.305 41.735 149.115 ;
        RECT 41.745 148.305 43.575 149.115 ;
        RECT 44.055 148.245 44.485 149.030 ;
        RECT 44.505 148.305 50.015 149.115 ;
        RECT 50.025 148.305 53.695 149.115 ;
        RECT 53.725 148.205 55.075 149.115 ;
        RECT 55.545 148.205 56.895 149.115 ;
        RECT 57.020 148.435 60.485 149.115 ;
        RECT 60.745 149.085 60.915 149.305 ;
        RECT 63.040 149.135 63.210 149.325 ;
        RECT 63.505 149.135 63.675 149.325 ;
        RECT 66.265 149.115 66.435 149.305 ;
        RECT 66.725 149.115 66.895 149.305 ;
        RECT 69.485 149.275 69.655 149.325 ;
        RECT 69.020 149.165 69.140 149.275 ;
        RECT 69.480 149.165 69.655 149.275 ;
        RECT 69.485 149.135 69.655 149.165 ;
        RECT 70.410 149.115 70.580 149.305 ;
        RECT 72.705 149.135 72.875 149.325 ;
        RECT 74.090 149.305 74.260 149.325 ;
        RECT 74.085 149.135 74.260 149.305 ;
        RECT 75.465 149.135 75.635 149.325 ;
        RECT 74.085 149.115 74.255 149.135 ;
        RECT 79.605 149.115 79.775 149.305 ;
        RECT 80.985 149.135 81.155 149.325 ;
        RECT 83.285 149.135 83.455 149.325 ;
        RECT 85.125 149.115 85.295 149.305 ;
        RECT 88.805 149.135 88.975 149.325 ;
        RECT 90.640 149.165 90.760 149.275 ;
        RECT 92.025 149.115 92.195 149.325 ;
        RECT 62.870 149.085 63.815 149.115 ;
        RECT 60.745 148.885 63.815 149.085 ;
        RECT 57.020 148.205 57.940 148.435 ;
        RECT 60.605 148.405 63.815 148.885 ;
        RECT 63.835 148.435 66.575 149.115 ;
        RECT 60.605 148.205 61.535 148.405 ;
        RECT 62.870 148.205 63.815 148.405 ;
        RECT 66.585 148.305 69.335 149.115 ;
        RECT 69.815 148.245 70.245 149.030 ;
        RECT 70.265 148.435 73.935 149.115 ;
        RECT 70.265 148.205 71.190 148.435 ;
        RECT 73.945 148.305 79.455 149.115 ;
        RECT 79.465 148.305 84.975 149.115 ;
        RECT 84.985 148.305 90.495 149.115 ;
        RECT 90.965 148.305 92.335 149.115 ;
      LAYER nwell ;
        RECT 18.090 145.085 92.530 147.915 ;
      LAYER pwell ;
        RECT 18.285 143.885 19.655 144.695 ;
        RECT 19.665 143.885 25.175 144.695 ;
        RECT 25.185 143.885 30.695 144.695 ;
        RECT 31.175 143.970 31.605 144.755 ;
        RECT 31.625 143.885 37.135 144.695 ;
        RECT 37.145 143.885 42.655 144.695 ;
        RECT 46.180 144.565 47.090 144.785 ;
        RECT 48.625 144.565 49.975 144.795 ;
        RECT 42.665 143.885 49.975 144.565 ;
        RECT 50.025 144.565 50.950 144.795 ;
        RECT 50.025 143.885 53.695 144.565 ;
        RECT 53.705 143.885 56.875 144.795 ;
        RECT 56.935 143.970 57.365 144.755 ;
        RECT 57.425 144.565 58.775 144.795 ;
        RECT 60.310 144.565 61.220 144.785 ;
        RECT 68.720 144.565 69.630 144.785 ;
        RECT 71.165 144.565 72.515 144.795 ;
        RECT 57.425 143.885 64.735 144.565 ;
        RECT 65.205 143.885 72.515 144.565 ;
        RECT 72.565 143.885 78.075 144.695 ;
        RECT 78.085 143.885 81.755 144.695 ;
        RECT 82.695 143.970 83.125 144.755 ;
        RECT 83.145 143.885 88.655 144.695 ;
        RECT 88.665 143.885 90.495 144.695 ;
        RECT 90.965 143.885 92.335 144.695 ;
        RECT 18.425 143.675 18.595 143.885 ;
        RECT 19.805 143.675 19.975 143.885 ;
        RECT 25.325 143.675 25.495 143.885 ;
        RECT 30.845 143.835 31.015 143.865 ;
        RECT 30.840 143.725 31.015 143.835 ;
        RECT 30.845 143.675 31.015 143.725 ;
        RECT 31.765 143.695 31.935 143.885 ;
        RECT 36.365 143.675 36.535 143.865 ;
        RECT 37.285 143.695 37.455 143.885 ;
        RECT 41.885 143.675 42.055 143.865 ;
        RECT 42.805 143.695 42.975 143.885 ;
        RECT 43.720 143.725 43.840 143.835 ;
        RECT 45.560 143.675 45.730 143.865 ;
        RECT 46.025 143.675 46.195 143.865 ;
        RECT 50.170 143.695 50.340 143.885 ;
        RECT 51.545 143.675 51.715 143.865 ;
        RECT 56.605 143.695 56.775 143.885 ;
        RECT 57.065 143.675 57.235 143.865 ;
        RECT 62.585 143.675 62.755 143.865 ;
        RECT 64.425 143.695 64.595 143.885 ;
        RECT 64.880 143.725 65.000 143.835 ;
        RECT 65.345 143.695 65.515 143.885 ;
        RECT 66.260 143.725 66.380 143.835 ;
        RECT 67.640 143.675 67.810 143.865 ;
        RECT 68.105 143.675 68.275 143.865 ;
        RECT 70.405 143.675 70.575 143.865 ;
        RECT 72.705 143.695 72.875 143.885 ;
        RECT 75.925 143.675 76.095 143.865 ;
        RECT 78.225 143.695 78.395 143.885 ;
        RECT 81.445 143.675 81.615 143.865 ;
        RECT 81.915 143.730 82.075 143.840 ;
        RECT 83.285 143.695 83.455 143.885 ;
        RECT 86.965 143.675 87.135 143.865 ;
        RECT 88.805 143.695 88.975 143.885 ;
        RECT 90.640 143.725 90.760 143.835 ;
        RECT 92.025 143.675 92.195 143.885 ;
        RECT 18.285 142.865 19.655 143.675 ;
        RECT 19.665 142.865 25.175 143.675 ;
        RECT 25.185 142.865 30.695 143.675 ;
        RECT 30.705 142.865 36.215 143.675 ;
        RECT 36.225 142.865 41.735 143.675 ;
        RECT 41.745 142.865 43.575 143.675 ;
        RECT 44.055 142.805 44.485 143.590 ;
        RECT 44.525 142.765 45.875 143.675 ;
        RECT 45.885 142.865 51.395 143.675 ;
        RECT 51.405 142.865 56.915 143.675 ;
        RECT 56.925 142.865 62.435 143.675 ;
        RECT 62.445 142.865 66.115 143.675 ;
        RECT 66.605 142.765 67.955 143.675 ;
        RECT 67.965 142.865 69.795 143.675 ;
        RECT 69.815 142.805 70.245 143.590 ;
        RECT 70.265 142.865 75.775 143.675 ;
        RECT 75.785 142.865 81.295 143.675 ;
        RECT 81.305 142.865 86.815 143.675 ;
        RECT 86.825 142.865 90.495 143.675 ;
        RECT 90.965 142.865 92.335 143.675 ;
      LAYER nwell ;
        RECT 18.090 139.645 92.530 142.475 ;
      LAYER pwell ;
        RECT 18.285 138.445 19.655 139.255 ;
        RECT 19.665 138.445 25.175 139.255 ;
        RECT 25.185 138.445 30.695 139.255 ;
        RECT 31.175 138.530 31.605 139.315 ;
        RECT 31.625 138.445 37.135 139.255 ;
        RECT 37.145 138.445 42.655 139.255 ;
        RECT 42.665 138.445 48.175 139.255 ;
        RECT 48.185 138.445 53.695 139.255 ;
        RECT 53.705 138.445 56.455 139.255 ;
        RECT 56.935 138.530 57.365 139.315 ;
        RECT 57.385 138.445 62.895 139.255 ;
        RECT 62.905 138.445 68.415 139.255 ;
        RECT 68.425 138.445 73.935 139.255 ;
        RECT 73.945 138.445 79.455 139.255 ;
        RECT 79.465 138.445 82.215 139.255 ;
        RECT 82.695 138.530 83.125 139.315 ;
        RECT 83.145 138.445 88.655 139.255 ;
        RECT 88.665 138.445 90.495 139.255 ;
        RECT 90.965 138.445 92.335 139.255 ;
        RECT 18.425 138.235 18.595 138.445 ;
        RECT 19.805 138.235 19.975 138.445 ;
        RECT 25.325 138.235 25.495 138.445 ;
        RECT 30.845 138.395 31.015 138.425 ;
        RECT 30.840 138.285 31.015 138.395 ;
        RECT 30.845 138.235 31.015 138.285 ;
        RECT 31.765 138.255 31.935 138.445 ;
        RECT 36.365 138.235 36.535 138.425 ;
        RECT 37.285 138.255 37.455 138.445 ;
        RECT 41.885 138.235 42.055 138.425 ;
        RECT 42.805 138.255 42.975 138.445 ;
        RECT 43.720 138.285 43.840 138.395 ;
        RECT 44.645 138.235 44.815 138.425 ;
        RECT 48.325 138.255 48.495 138.445 ;
        RECT 50.165 138.235 50.335 138.425 ;
        RECT 53.845 138.255 54.015 138.445 ;
        RECT 55.685 138.235 55.855 138.425 ;
        RECT 56.600 138.285 56.720 138.395 ;
        RECT 57.525 138.255 57.695 138.445 ;
        RECT 61.205 138.235 61.375 138.425 ;
        RECT 63.045 138.255 63.215 138.445 ;
        RECT 66.725 138.235 66.895 138.425 ;
        RECT 68.565 138.255 68.735 138.445 ;
        RECT 69.480 138.285 69.600 138.395 ;
        RECT 70.405 138.235 70.575 138.425 ;
        RECT 74.085 138.255 74.255 138.445 ;
        RECT 75.925 138.235 76.095 138.425 ;
        RECT 79.605 138.255 79.775 138.445 ;
        RECT 81.445 138.235 81.615 138.425 ;
        RECT 82.360 138.285 82.480 138.395 ;
        RECT 83.285 138.255 83.455 138.445 ;
        RECT 86.965 138.235 87.135 138.425 ;
        RECT 88.805 138.255 88.975 138.445 ;
        RECT 90.640 138.285 90.760 138.395 ;
        RECT 92.025 138.235 92.195 138.445 ;
        RECT 18.285 137.425 19.655 138.235 ;
        RECT 19.665 137.425 25.175 138.235 ;
        RECT 25.185 137.425 30.695 138.235 ;
        RECT 30.705 137.425 36.215 138.235 ;
        RECT 36.225 137.425 41.735 138.235 ;
        RECT 41.745 137.425 43.575 138.235 ;
        RECT 44.055 137.365 44.485 138.150 ;
        RECT 44.505 137.425 50.015 138.235 ;
        RECT 50.025 137.425 55.535 138.235 ;
        RECT 55.545 137.425 61.055 138.235 ;
        RECT 61.065 137.425 66.575 138.235 ;
        RECT 66.585 137.425 69.335 138.235 ;
        RECT 69.815 137.365 70.245 138.150 ;
        RECT 70.265 137.425 75.775 138.235 ;
        RECT 75.785 137.425 81.295 138.235 ;
        RECT 81.305 137.425 86.815 138.235 ;
        RECT 86.825 137.425 90.495 138.235 ;
        RECT 90.965 137.425 92.335 138.235 ;
      LAYER nwell ;
        RECT 18.090 134.205 92.530 137.035 ;
      LAYER pwell ;
        RECT 18.285 133.005 19.655 133.815 ;
        RECT 19.665 133.005 25.175 133.815 ;
        RECT 25.185 133.005 30.695 133.815 ;
        RECT 31.175 133.090 31.605 133.875 ;
        RECT 31.625 133.005 37.135 133.815 ;
        RECT 37.145 133.005 42.655 133.815 ;
        RECT 42.665 133.005 44.035 133.815 ;
        RECT 44.055 133.090 44.485 133.875 ;
        RECT 44.505 133.005 50.015 133.815 ;
        RECT 50.025 133.005 55.535 133.815 ;
        RECT 55.545 133.005 56.915 133.815 ;
        RECT 56.935 133.090 57.365 133.875 ;
        RECT 57.385 133.005 62.895 133.815 ;
        RECT 62.905 133.005 68.415 133.815 ;
        RECT 68.425 133.005 69.795 133.815 ;
        RECT 69.815 133.090 70.245 133.875 ;
        RECT 70.265 133.005 75.775 133.815 ;
        RECT 75.785 133.005 81.295 133.815 ;
        RECT 81.305 133.005 82.675 133.815 ;
        RECT 82.695 133.090 83.125 133.875 ;
        RECT 83.145 133.005 88.655 133.815 ;
        RECT 88.665 133.005 90.495 133.815 ;
        RECT 90.965 133.005 92.335 133.815 ;
        RECT 18.425 132.815 18.595 133.005 ;
        RECT 19.805 132.815 19.975 133.005 ;
        RECT 25.325 132.815 25.495 133.005 ;
        RECT 30.840 132.845 30.960 132.955 ;
        RECT 31.765 132.815 31.935 133.005 ;
        RECT 37.285 132.815 37.455 133.005 ;
        RECT 42.805 132.815 42.975 133.005 ;
        RECT 44.645 132.815 44.815 133.005 ;
        RECT 50.165 132.815 50.335 133.005 ;
        RECT 55.685 132.815 55.855 133.005 ;
        RECT 57.525 132.815 57.695 133.005 ;
        RECT 63.045 132.815 63.215 133.005 ;
        RECT 68.565 132.815 68.735 133.005 ;
        RECT 70.405 132.815 70.575 133.005 ;
        RECT 75.925 132.815 76.095 133.005 ;
        RECT 81.445 132.815 81.615 133.005 ;
        RECT 83.285 132.815 83.455 133.005 ;
        RECT 88.805 132.815 88.975 133.005 ;
        RECT 90.640 132.845 90.760 132.955 ;
        RECT 92.025 132.815 92.195 133.005 ;
        RECT 106.000 70.700 108.010 114.980 ;
        RECT 110.000 96.000 112.010 141.980 ;
        RECT 113.000 96.000 115.010 141.980 ;
        RECT 116.000 96.000 118.010 141.980 ;
        RECT 119.000 96.000 121.010 141.980 ;
        RECT 122.000 96.000 124.010 141.980 ;
        RECT 125.000 96.000 127.010 141.980 ;
        RECT 128.000 96.000 130.010 141.980 ;
        RECT 131.000 96.000 133.010 141.980 ;
        RECT 103.600 70.300 108.010 70.700 ;
        RECT 106.000 69.000 108.010 70.300 ;
        RECT 110.000 69.000 112.010 94.980 ;
        RECT 113.000 69.000 115.010 94.980 ;
        RECT 116.000 69.000 118.010 94.980 ;
        RECT 119.000 69.000 121.010 94.980 ;
        RECT 122.000 69.000 124.010 94.980 ;
        RECT 125.000 69.000 127.010 94.980 ;
        RECT 128.000 69.000 130.010 94.980 ;
      LAYER li1 ;
        RECT 18.280 206.255 92.340 206.425 ;
        RECT 18.365 205.165 19.575 206.255 ;
        RECT 18.365 204.455 18.885 204.995 ;
        RECT 19.055 204.625 19.575 205.165 ;
        RECT 20.205 205.285 20.475 206.055 ;
        RECT 20.645 205.475 20.975 206.255 ;
        RECT 21.180 205.650 21.365 206.055 ;
        RECT 21.535 205.830 21.870 206.255 ;
        RECT 21.180 205.475 21.845 205.650 ;
        RECT 20.205 205.115 21.335 205.285 ;
        RECT 18.365 203.705 19.575 204.455 ;
        RECT 20.205 204.205 20.375 205.115 ;
        RECT 20.545 204.365 20.905 204.945 ;
        RECT 21.085 204.615 21.335 205.115 ;
        RECT 21.505 204.445 21.845 205.475 ;
        RECT 22.045 205.165 25.555 206.255 ;
        RECT 21.160 204.275 21.845 204.445 ;
        RECT 22.045 204.475 23.695 204.995 ;
        RECT 23.865 204.645 25.555 205.165 ;
        RECT 26.645 205.285 26.915 206.055 ;
        RECT 27.085 205.475 27.415 206.255 ;
        RECT 27.620 205.650 27.805 206.055 ;
        RECT 27.975 205.830 28.310 206.255 ;
        RECT 27.620 205.475 28.285 205.650 ;
        RECT 26.645 205.115 27.775 205.285 ;
        RECT 20.205 203.875 20.465 204.205 ;
        RECT 20.675 203.705 20.950 204.185 ;
        RECT 21.160 203.875 21.365 204.275 ;
        RECT 21.535 203.705 21.870 204.105 ;
        RECT 22.045 203.705 25.555 204.475 ;
        RECT 26.645 204.205 26.815 205.115 ;
        RECT 26.985 204.365 27.345 204.945 ;
        RECT 27.525 204.615 27.775 205.115 ;
        RECT 27.945 204.445 28.285 205.475 ;
        RECT 28.485 205.165 31.075 206.255 ;
        RECT 27.600 204.275 28.285 204.445 ;
        RECT 28.485 204.475 29.695 204.995 ;
        RECT 29.865 204.645 31.075 205.165 ;
        RECT 31.245 205.090 31.535 206.255 ;
        RECT 31.705 205.165 32.915 206.255 ;
        RECT 26.645 203.875 26.905 204.205 ;
        RECT 27.115 203.705 27.390 204.185 ;
        RECT 27.600 203.875 27.805 204.275 ;
        RECT 27.975 203.705 28.310 204.105 ;
        RECT 28.485 203.705 31.075 204.475 ;
        RECT 31.705 204.455 32.225 204.995 ;
        RECT 32.395 204.625 32.915 205.165 ;
        RECT 33.165 205.325 33.345 206.085 ;
        RECT 33.525 205.495 33.855 206.255 ;
        RECT 33.165 205.155 33.840 205.325 ;
        RECT 34.025 205.180 34.295 206.085 ;
        RECT 33.670 205.010 33.840 205.155 ;
        RECT 33.105 204.605 33.445 204.975 ;
        RECT 33.670 204.680 33.945 205.010 ;
        RECT 31.245 203.705 31.535 204.430 ;
        RECT 31.705 203.705 32.915 204.455 ;
        RECT 33.670 204.425 33.840 204.680 ;
        RECT 33.175 204.255 33.840 204.425 ;
        RECT 34.115 204.380 34.295 205.180 ;
        RECT 34.465 205.165 37.975 206.255 ;
        RECT 33.175 203.875 33.345 204.255 ;
        RECT 33.525 203.705 33.855 204.085 ;
        RECT 34.035 203.875 34.295 204.380 ;
        RECT 34.465 204.475 36.115 204.995 ;
        RECT 36.285 204.645 37.975 205.165 ;
        RECT 38.605 205.115 38.880 206.085 ;
        RECT 39.090 205.455 39.370 206.255 ;
        RECT 39.540 205.745 41.155 206.075 ;
        RECT 39.540 205.405 40.715 205.575 ;
        RECT 39.540 205.285 39.710 205.405 ;
        RECT 39.050 205.115 39.710 205.285 ;
        RECT 34.465 203.705 37.975 204.475 ;
        RECT 38.605 204.380 38.775 205.115 ;
        RECT 39.050 204.945 39.220 205.115 ;
        RECT 39.970 204.945 40.215 205.235 ;
        RECT 40.385 205.115 40.715 205.405 ;
        RECT 40.975 204.945 41.145 205.505 ;
        RECT 41.395 205.115 41.655 206.255 ;
        RECT 41.905 205.325 42.085 206.085 ;
        RECT 42.265 205.495 42.595 206.255 ;
        RECT 41.905 205.155 42.580 205.325 ;
        RECT 42.765 205.180 43.035 206.085 ;
        RECT 42.410 205.010 42.580 205.155 ;
        RECT 38.945 204.615 39.220 204.945 ;
        RECT 39.390 204.615 40.215 204.945 ;
        RECT 40.430 204.615 41.145 204.945 ;
        RECT 41.315 204.695 41.650 204.945 ;
        RECT 39.050 204.445 39.220 204.615 ;
        RECT 40.895 204.525 41.145 204.615 ;
        RECT 41.845 204.605 42.185 204.975 ;
        RECT 42.410 204.680 42.685 205.010 ;
        RECT 38.605 204.035 38.880 204.380 ;
        RECT 39.050 204.275 40.715 204.445 ;
        RECT 39.070 203.705 39.445 204.105 ;
        RECT 39.615 203.925 39.785 204.275 ;
        RECT 39.955 203.705 40.285 204.105 ;
        RECT 40.455 203.875 40.715 204.275 ;
        RECT 40.895 204.105 41.225 204.525 ;
        RECT 41.395 203.705 41.655 204.525 ;
        RECT 42.410 204.425 42.580 204.680 ;
        RECT 41.915 204.255 42.580 204.425 ;
        RECT 42.855 204.380 43.035 205.180 ;
        RECT 44.125 205.090 44.415 206.255 ;
        RECT 44.585 205.165 45.795 206.255 ;
        RECT 44.585 204.455 45.105 204.995 ;
        RECT 45.275 204.625 45.795 205.165 ;
        RECT 46.045 205.325 46.225 206.085 ;
        RECT 46.405 205.495 46.735 206.255 ;
        RECT 46.045 205.155 46.720 205.325 ;
        RECT 46.905 205.180 47.175 206.085 ;
        RECT 46.550 205.010 46.720 205.155 ;
        RECT 45.985 204.605 46.325 204.975 ;
        RECT 46.550 204.680 46.825 205.010 ;
        RECT 41.915 203.875 42.085 204.255 ;
        RECT 42.265 203.705 42.595 204.085 ;
        RECT 42.775 203.875 43.035 204.380 ;
        RECT 44.125 203.705 44.415 204.430 ;
        RECT 44.585 203.705 45.795 204.455 ;
        RECT 46.550 204.425 46.720 204.680 ;
        RECT 46.055 204.255 46.720 204.425 ;
        RECT 46.995 204.380 47.175 205.180 ;
        RECT 47.345 205.165 50.855 206.255 ;
        RECT 51.025 205.165 52.235 206.255 ;
        RECT 46.055 203.875 46.225 204.255 ;
        RECT 46.405 203.705 46.735 204.085 ;
        RECT 46.915 203.875 47.175 204.380 ;
        RECT 47.345 204.475 48.995 204.995 ;
        RECT 49.165 204.645 50.855 205.165 ;
        RECT 47.345 203.705 50.855 204.475 ;
        RECT 51.025 204.455 51.545 204.995 ;
        RECT 51.715 204.625 52.235 205.165 ;
        RECT 52.485 205.325 52.665 206.085 ;
        RECT 52.845 205.495 53.175 206.255 ;
        RECT 52.485 205.155 53.160 205.325 ;
        RECT 53.345 205.180 53.615 206.085 ;
        RECT 52.990 205.010 53.160 205.155 ;
        RECT 52.425 204.605 52.765 204.975 ;
        RECT 52.990 204.680 53.265 205.010 ;
        RECT 51.025 203.705 52.235 204.455 ;
        RECT 52.990 204.425 53.160 204.680 ;
        RECT 52.495 204.255 53.160 204.425 ;
        RECT 53.435 204.380 53.615 205.180 ;
        RECT 53.785 205.165 56.375 206.255 ;
        RECT 52.495 203.875 52.665 204.255 ;
        RECT 52.845 203.705 53.175 204.085 ;
        RECT 53.355 203.875 53.615 204.380 ;
        RECT 53.785 204.475 54.995 204.995 ;
        RECT 55.165 204.645 56.375 205.165 ;
        RECT 57.005 205.090 57.295 206.255 ;
        RECT 57.465 205.115 57.740 206.085 ;
        RECT 57.950 205.455 58.230 206.255 ;
        RECT 58.400 205.745 60.015 206.075 ;
        RECT 58.400 205.405 59.575 205.575 ;
        RECT 58.400 205.285 58.570 205.405 ;
        RECT 57.910 205.115 58.570 205.285 ;
        RECT 53.785 203.705 56.375 204.475 ;
        RECT 57.005 203.705 57.295 204.430 ;
        RECT 57.465 204.380 57.635 205.115 ;
        RECT 57.910 204.945 58.080 205.115 ;
        RECT 58.830 204.945 59.075 205.235 ;
        RECT 59.245 205.115 59.575 205.405 ;
        RECT 59.835 204.945 60.005 205.505 ;
        RECT 60.255 205.115 60.515 206.255 ;
        RECT 60.765 205.325 60.945 206.085 ;
        RECT 61.125 205.495 61.455 206.255 ;
        RECT 60.765 205.155 61.440 205.325 ;
        RECT 61.625 205.180 61.895 206.085 ;
        RECT 61.270 205.010 61.440 205.155 ;
        RECT 57.805 204.615 58.080 204.945 ;
        RECT 58.250 204.615 59.075 204.945 ;
        RECT 59.290 204.615 60.005 204.945 ;
        RECT 60.175 204.695 60.510 204.945 ;
        RECT 57.910 204.445 58.080 204.615 ;
        RECT 59.755 204.525 60.005 204.615 ;
        RECT 60.705 204.605 61.045 204.975 ;
        RECT 61.270 204.680 61.545 205.010 ;
        RECT 57.465 204.035 57.740 204.380 ;
        RECT 57.910 204.275 59.575 204.445 ;
        RECT 57.930 203.705 58.305 204.105 ;
        RECT 58.475 203.925 58.645 204.275 ;
        RECT 58.815 203.705 59.145 204.105 ;
        RECT 59.315 203.875 59.575 204.275 ;
        RECT 59.755 204.105 60.085 204.525 ;
        RECT 60.255 203.705 60.515 204.525 ;
        RECT 61.270 204.425 61.440 204.680 ;
        RECT 60.775 204.255 61.440 204.425 ;
        RECT 61.715 204.380 61.895 205.180 ;
        RECT 62.065 205.165 64.655 206.255 ;
        RECT 60.775 203.875 60.945 204.255 ;
        RECT 61.125 203.705 61.455 204.085 ;
        RECT 61.635 203.875 61.895 204.380 ;
        RECT 62.065 204.475 63.275 204.995 ;
        RECT 63.445 204.645 64.655 205.165 ;
        RECT 65.365 205.325 65.545 206.085 ;
        RECT 65.725 205.495 66.055 206.255 ;
        RECT 65.365 205.155 66.040 205.325 ;
        RECT 66.225 205.180 66.495 206.085 ;
        RECT 65.870 205.010 66.040 205.155 ;
        RECT 65.305 204.605 65.645 204.975 ;
        RECT 65.870 204.680 66.145 205.010 ;
        RECT 62.065 203.705 64.655 204.475 ;
        RECT 65.870 204.425 66.040 204.680 ;
        RECT 65.375 204.255 66.040 204.425 ;
        RECT 66.315 204.380 66.495 205.180 ;
        RECT 66.665 205.165 69.255 206.255 ;
        RECT 65.375 203.875 65.545 204.255 ;
        RECT 65.725 203.705 66.055 204.085 ;
        RECT 66.235 203.875 66.495 204.380 ;
        RECT 66.665 204.475 67.875 204.995 ;
        RECT 68.045 204.645 69.255 205.165 ;
        RECT 69.885 205.090 70.175 206.255 ;
        RECT 70.345 205.165 71.555 206.255 ;
        RECT 66.665 203.705 69.255 204.475 ;
        RECT 70.345 204.455 70.865 204.995 ;
        RECT 71.035 204.625 71.555 205.165 ;
        RECT 71.805 205.325 71.985 206.085 ;
        RECT 72.165 205.495 72.495 206.255 ;
        RECT 71.805 205.155 72.480 205.325 ;
        RECT 72.665 205.180 72.935 206.085 ;
        RECT 72.310 205.010 72.480 205.155 ;
        RECT 71.745 204.605 72.085 204.975 ;
        RECT 72.310 204.680 72.585 205.010 ;
        RECT 69.885 203.705 70.175 204.430 ;
        RECT 70.345 203.705 71.555 204.455 ;
        RECT 72.310 204.425 72.480 204.680 ;
        RECT 71.815 204.255 72.480 204.425 ;
        RECT 72.755 204.380 72.935 205.180 ;
        RECT 73.105 205.165 76.615 206.255 ;
        RECT 76.785 205.165 77.995 206.255 ;
        RECT 71.815 203.875 71.985 204.255 ;
        RECT 72.165 203.705 72.495 204.085 ;
        RECT 72.675 203.875 72.935 204.380 ;
        RECT 73.105 204.475 74.755 204.995 ;
        RECT 74.925 204.645 76.615 205.165 ;
        RECT 73.105 203.705 76.615 204.475 ;
        RECT 76.785 204.455 77.305 204.995 ;
        RECT 77.475 204.625 77.995 205.165 ;
        RECT 78.165 205.180 78.435 206.085 ;
        RECT 78.605 205.495 78.935 206.255 ;
        RECT 79.115 205.325 79.295 206.085 ;
        RECT 79.735 205.530 80.065 206.255 ;
        RECT 76.785 203.705 77.995 204.455 ;
        RECT 78.165 204.380 78.345 205.180 ;
        RECT 78.620 205.155 79.295 205.325 ;
        RECT 78.620 205.010 78.790 205.155 ;
        RECT 78.515 204.680 78.790 205.010 ;
        RECT 78.620 204.425 78.790 204.680 ;
        RECT 79.015 204.605 79.355 204.975 ;
        RECT 78.165 203.875 78.425 204.380 ;
        RECT 78.620 204.255 79.285 204.425 ;
        RECT 78.605 203.705 78.935 204.085 ;
        RECT 79.115 203.875 79.285 204.255 ;
        RECT 79.545 203.875 80.065 205.360 ;
        RECT 80.235 204.535 80.755 206.085 ;
        RECT 80.925 205.165 82.595 206.255 ;
        RECT 80.925 204.475 81.675 204.995 ;
        RECT 81.845 204.645 82.595 205.165 ;
        RECT 82.765 205.090 83.055 206.255 ;
        RECT 83.225 205.165 84.435 206.255 ;
        RECT 80.235 203.705 80.575 204.365 ;
        RECT 80.925 203.705 82.595 204.475 ;
        RECT 83.225 204.455 83.745 204.995 ;
        RECT 83.915 204.625 84.435 205.165 ;
        RECT 84.695 205.325 84.865 206.085 ;
        RECT 85.045 205.495 85.375 206.255 ;
        RECT 84.695 205.155 85.360 205.325 ;
        RECT 85.545 205.180 85.815 206.085 ;
        RECT 85.190 205.010 85.360 205.155 ;
        RECT 84.625 204.605 84.955 204.975 ;
        RECT 85.190 204.680 85.475 205.010 ;
        RECT 82.765 203.705 83.055 204.430 ;
        RECT 83.225 203.705 84.435 204.455 ;
        RECT 85.190 204.425 85.360 204.680 ;
        RECT 84.695 204.255 85.360 204.425 ;
        RECT 85.645 204.380 85.815 205.180 ;
        RECT 85.985 205.165 89.495 206.255 ;
        RECT 89.665 205.165 90.875 206.255 ;
        RECT 84.695 203.875 84.865 204.255 ;
        RECT 85.045 203.705 85.375 204.085 ;
        RECT 85.555 203.875 85.815 204.380 ;
        RECT 85.985 204.475 87.635 204.995 ;
        RECT 87.805 204.645 89.495 205.165 ;
        RECT 85.985 203.705 89.495 204.475 ;
        RECT 89.665 204.455 90.185 204.995 ;
        RECT 90.355 204.625 90.875 205.165 ;
        RECT 91.045 205.165 92.255 206.255 ;
        RECT 91.045 204.625 91.565 205.165 ;
        RECT 91.735 204.455 92.255 204.995 ;
        RECT 89.665 203.705 90.875 204.455 ;
        RECT 91.045 203.705 92.255 204.455 ;
        RECT 18.280 203.535 92.340 203.705 ;
        RECT 18.365 202.785 19.575 203.535 ;
        RECT 19.745 202.990 25.090 203.535 ;
        RECT 25.265 202.990 30.610 203.535 ;
        RECT 18.365 202.245 18.885 202.785 ;
        RECT 19.055 202.075 19.575 202.615 ;
        RECT 21.330 202.160 21.670 202.990 ;
        RECT 18.365 200.985 19.575 202.075 ;
        RECT 23.150 201.420 23.500 202.670 ;
        RECT 26.850 202.160 27.190 202.990 ;
        RECT 30.785 202.765 33.375 203.535 ;
        RECT 34.055 202.880 34.385 203.315 ;
        RECT 34.555 202.925 34.725 203.535 ;
        RECT 34.005 202.795 34.385 202.880 ;
        RECT 34.895 202.795 35.225 203.320 ;
        RECT 35.485 203.005 35.695 203.535 ;
        RECT 35.970 203.085 36.755 203.255 ;
        RECT 36.925 203.085 37.330 203.255 ;
        RECT 28.670 201.420 29.020 202.670 ;
        RECT 30.785 202.245 31.995 202.765 ;
        RECT 34.005 202.755 34.230 202.795 ;
        RECT 32.165 202.075 33.375 202.595 ;
        RECT 19.745 200.985 25.090 201.420 ;
        RECT 25.265 200.985 30.610 201.420 ;
        RECT 30.785 200.985 33.375 202.075 ;
        RECT 34.005 202.175 34.175 202.755 ;
        RECT 34.895 202.625 35.095 202.795 ;
        RECT 35.970 202.625 36.140 203.085 ;
        RECT 34.345 202.295 35.095 202.625 ;
        RECT 35.265 202.295 36.140 202.625 ;
        RECT 34.005 202.125 34.220 202.175 ;
        RECT 34.005 202.045 34.395 202.125 ;
        RECT 34.065 201.200 34.395 202.045 ;
        RECT 34.905 202.090 35.095 202.295 ;
        RECT 34.565 200.985 34.735 201.995 ;
        RECT 34.905 201.715 35.800 202.090 ;
        RECT 34.905 201.155 35.245 201.715 ;
        RECT 35.475 200.985 35.790 201.485 ;
        RECT 35.970 201.455 36.140 202.295 ;
        RECT 36.310 202.585 36.775 202.915 ;
        RECT 37.160 202.855 37.330 203.085 ;
        RECT 37.510 203.035 37.880 203.535 ;
        RECT 38.200 203.085 38.875 203.255 ;
        RECT 39.070 203.085 39.405 203.255 ;
        RECT 36.310 201.625 36.630 202.585 ;
        RECT 37.160 202.555 37.990 202.855 ;
        RECT 36.800 201.655 36.990 202.375 ;
        RECT 37.160 201.485 37.330 202.555 ;
        RECT 37.790 202.525 37.990 202.555 ;
        RECT 37.500 202.305 37.670 202.375 ;
        RECT 38.200 202.305 38.370 203.085 ;
        RECT 39.235 202.945 39.405 203.085 ;
        RECT 39.575 203.075 39.825 203.535 ;
        RECT 37.500 202.135 38.370 202.305 ;
        RECT 38.540 202.665 39.065 202.885 ;
        RECT 39.235 202.815 39.460 202.945 ;
        RECT 37.500 202.045 38.010 202.135 ;
        RECT 35.970 201.285 36.855 201.455 ;
        RECT 37.080 201.155 37.330 201.485 ;
        RECT 37.500 200.985 37.670 201.785 ;
        RECT 37.840 201.430 38.010 202.045 ;
        RECT 38.540 201.965 38.710 202.665 ;
        RECT 38.180 201.600 38.710 201.965 ;
        RECT 38.880 201.900 39.120 202.495 ;
        RECT 39.290 201.710 39.460 202.815 ;
        RECT 39.630 201.955 39.910 202.905 ;
        RECT 39.155 201.580 39.460 201.710 ;
        RECT 37.840 201.260 38.945 201.430 ;
        RECT 39.155 201.155 39.405 201.580 ;
        RECT 39.575 200.985 39.840 201.445 ;
        RECT 40.080 201.155 40.265 203.275 ;
        RECT 40.435 203.155 40.765 203.535 ;
        RECT 40.935 202.985 41.105 203.275 ;
        RECT 40.440 202.815 41.105 202.985 ;
        RECT 40.440 201.825 40.670 202.815 ;
        RECT 41.370 202.695 41.630 203.535 ;
        RECT 41.805 202.790 42.060 203.365 ;
        RECT 42.230 203.155 42.560 203.535 ;
        RECT 42.775 202.985 42.945 203.365 ;
        RECT 42.230 202.815 42.945 202.985 ;
        RECT 40.840 201.995 41.190 202.645 ;
        RECT 40.440 201.655 41.105 201.825 ;
        RECT 40.435 200.985 40.765 201.485 ;
        RECT 40.935 201.155 41.105 201.655 ;
        RECT 41.370 200.985 41.630 202.135 ;
        RECT 41.805 202.060 41.975 202.790 ;
        RECT 42.230 202.625 42.400 202.815 ;
        RECT 44.125 202.810 44.415 203.535 ;
        RECT 44.635 202.880 44.965 203.315 ;
        RECT 45.135 202.925 45.305 203.535 ;
        RECT 44.585 202.795 44.965 202.880 ;
        RECT 45.475 202.795 45.805 203.320 ;
        RECT 46.065 203.005 46.275 203.535 ;
        RECT 46.550 203.085 47.335 203.255 ;
        RECT 47.505 203.085 47.910 203.255 ;
        RECT 44.585 202.755 44.810 202.795 ;
        RECT 42.145 202.295 42.400 202.625 ;
        RECT 42.230 202.085 42.400 202.295 ;
        RECT 42.680 202.265 43.035 202.635 ;
        RECT 44.585 202.175 44.755 202.755 ;
        RECT 45.475 202.625 45.675 202.795 ;
        RECT 46.550 202.625 46.720 203.085 ;
        RECT 44.925 202.295 45.675 202.625 ;
        RECT 45.845 202.295 46.720 202.625 ;
        RECT 41.805 201.155 42.060 202.060 ;
        RECT 42.230 201.915 42.945 202.085 ;
        RECT 42.230 200.985 42.560 201.745 ;
        RECT 42.775 201.155 42.945 201.915 ;
        RECT 44.125 200.985 44.415 202.150 ;
        RECT 44.585 202.125 44.800 202.175 ;
        RECT 44.585 202.045 44.975 202.125 ;
        RECT 44.645 201.200 44.975 202.045 ;
        RECT 45.485 202.090 45.675 202.295 ;
        RECT 45.145 200.985 45.315 201.995 ;
        RECT 45.485 201.715 46.380 202.090 ;
        RECT 45.485 201.155 45.825 201.715 ;
        RECT 46.055 200.985 46.370 201.485 ;
        RECT 46.550 201.455 46.720 202.295 ;
        RECT 46.890 202.585 47.355 202.915 ;
        RECT 47.740 202.855 47.910 203.085 ;
        RECT 48.090 203.035 48.460 203.535 ;
        RECT 48.780 203.085 49.455 203.255 ;
        RECT 49.650 203.085 49.985 203.255 ;
        RECT 46.890 201.625 47.210 202.585 ;
        RECT 47.740 202.555 48.570 202.855 ;
        RECT 47.380 201.655 47.570 202.375 ;
        RECT 47.740 201.485 47.910 202.555 ;
        RECT 48.370 202.525 48.570 202.555 ;
        RECT 48.080 202.305 48.250 202.375 ;
        RECT 48.780 202.305 48.950 203.085 ;
        RECT 49.815 202.945 49.985 203.085 ;
        RECT 50.155 203.075 50.405 203.535 ;
        RECT 48.080 202.135 48.950 202.305 ;
        RECT 49.120 202.665 49.645 202.885 ;
        RECT 49.815 202.815 50.040 202.945 ;
        RECT 48.080 202.045 48.590 202.135 ;
        RECT 46.550 201.285 47.435 201.455 ;
        RECT 47.660 201.155 47.910 201.485 ;
        RECT 48.080 200.985 48.250 201.785 ;
        RECT 48.420 201.430 48.590 202.045 ;
        RECT 49.120 201.965 49.290 202.665 ;
        RECT 48.760 201.600 49.290 201.965 ;
        RECT 49.460 201.900 49.700 202.495 ;
        RECT 49.870 201.710 50.040 202.815 ;
        RECT 50.210 201.955 50.490 202.905 ;
        RECT 49.735 201.580 50.040 201.710 ;
        RECT 48.420 201.260 49.525 201.430 ;
        RECT 49.735 201.155 49.985 201.580 ;
        RECT 50.155 200.985 50.420 201.445 ;
        RECT 50.660 201.155 50.845 203.275 ;
        RECT 51.015 203.155 51.345 203.535 ;
        RECT 51.515 202.985 51.685 203.275 ;
        RECT 51.020 202.815 51.685 202.985 ;
        RECT 51.945 202.860 52.220 203.205 ;
        RECT 52.410 203.135 52.785 203.535 ;
        RECT 52.955 202.965 53.125 203.315 ;
        RECT 53.295 203.135 53.625 203.535 ;
        RECT 53.795 202.965 54.055 203.365 ;
        RECT 51.020 201.825 51.250 202.815 ;
        RECT 51.420 201.995 51.770 202.645 ;
        RECT 51.945 202.125 52.115 202.860 ;
        RECT 52.390 202.795 54.055 202.965 ;
        RECT 52.390 202.625 52.560 202.795 ;
        RECT 54.235 202.715 54.565 203.135 ;
        RECT 54.735 202.715 54.995 203.535 ;
        RECT 56.135 202.880 56.465 203.315 ;
        RECT 56.635 202.925 56.805 203.535 ;
        RECT 56.085 202.795 56.465 202.880 ;
        RECT 56.975 202.795 57.305 203.320 ;
        RECT 57.565 203.005 57.775 203.535 ;
        RECT 58.050 203.085 58.835 203.255 ;
        RECT 59.005 203.085 59.410 203.255 ;
        RECT 56.085 202.755 56.310 202.795 ;
        RECT 54.235 202.625 54.485 202.715 ;
        RECT 52.285 202.295 52.560 202.625 ;
        RECT 52.730 202.295 53.555 202.625 ;
        RECT 53.770 202.295 54.485 202.625 ;
        RECT 54.655 202.295 54.990 202.545 ;
        RECT 52.390 202.125 52.560 202.295 ;
        RECT 51.020 201.655 51.685 201.825 ;
        RECT 51.015 200.985 51.345 201.485 ;
        RECT 51.515 201.155 51.685 201.655 ;
        RECT 51.945 201.155 52.220 202.125 ;
        RECT 52.390 201.955 53.050 202.125 ;
        RECT 53.310 202.005 53.555 202.295 ;
        RECT 52.880 201.835 53.050 201.955 ;
        RECT 53.725 201.835 54.055 202.125 ;
        RECT 52.430 200.985 52.710 201.785 ;
        RECT 52.880 201.665 54.055 201.835 ;
        RECT 54.315 201.735 54.485 202.295 ;
        RECT 56.085 202.175 56.255 202.755 ;
        RECT 56.975 202.625 57.175 202.795 ;
        RECT 58.050 202.625 58.220 203.085 ;
        RECT 56.425 202.295 57.175 202.625 ;
        RECT 57.345 202.295 58.220 202.625 ;
        RECT 56.085 202.125 56.300 202.175 ;
        RECT 52.880 201.165 54.495 201.495 ;
        RECT 54.735 200.985 54.995 202.125 ;
        RECT 56.085 202.045 56.475 202.125 ;
        RECT 56.145 201.200 56.475 202.045 ;
        RECT 56.985 202.090 57.175 202.295 ;
        RECT 56.645 200.985 56.815 201.995 ;
        RECT 56.985 201.715 57.880 202.090 ;
        RECT 56.985 201.155 57.325 201.715 ;
        RECT 57.555 200.985 57.870 201.485 ;
        RECT 58.050 201.455 58.220 202.295 ;
        RECT 58.390 202.585 58.855 202.915 ;
        RECT 59.240 202.855 59.410 203.085 ;
        RECT 59.590 203.035 59.960 203.535 ;
        RECT 60.280 203.085 60.955 203.255 ;
        RECT 61.150 203.085 61.485 203.255 ;
        RECT 58.390 201.625 58.710 202.585 ;
        RECT 59.240 202.555 60.070 202.855 ;
        RECT 58.880 201.655 59.070 202.375 ;
        RECT 59.240 201.485 59.410 202.555 ;
        RECT 59.870 202.525 60.070 202.555 ;
        RECT 59.580 202.305 59.750 202.375 ;
        RECT 60.280 202.305 60.450 203.085 ;
        RECT 61.315 202.945 61.485 203.085 ;
        RECT 61.655 203.075 61.905 203.535 ;
        RECT 59.580 202.135 60.450 202.305 ;
        RECT 60.620 202.665 61.145 202.885 ;
        RECT 61.315 202.815 61.540 202.945 ;
        RECT 59.580 202.045 60.090 202.135 ;
        RECT 58.050 201.285 58.935 201.455 ;
        RECT 59.160 201.155 59.410 201.485 ;
        RECT 59.580 200.985 59.750 201.785 ;
        RECT 59.920 201.430 60.090 202.045 ;
        RECT 60.620 201.965 60.790 202.665 ;
        RECT 60.260 201.600 60.790 201.965 ;
        RECT 60.960 201.900 61.200 202.495 ;
        RECT 61.370 201.710 61.540 202.815 ;
        RECT 61.710 201.955 61.990 202.905 ;
        RECT 61.235 201.580 61.540 201.710 ;
        RECT 59.920 201.260 61.025 201.430 ;
        RECT 61.235 201.155 61.485 201.580 ;
        RECT 61.655 200.985 61.920 201.445 ;
        RECT 62.160 201.155 62.345 203.275 ;
        RECT 62.515 203.155 62.845 203.535 ;
        RECT 63.015 202.985 63.185 203.275 ;
        RECT 62.520 202.815 63.185 202.985 ;
        RECT 62.520 201.825 62.750 202.815 ;
        RECT 63.445 202.765 66.035 203.535 ;
        RECT 62.920 201.995 63.270 202.645 ;
        RECT 63.445 202.245 64.655 202.765 ;
        RECT 64.825 202.075 66.035 202.595 ;
        RECT 62.520 201.655 63.185 201.825 ;
        RECT 62.515 200.985 62.845 201.485 ;
        RECT 63.015 201.155 63.185 201.655 ;
        RECT 63.445 200.985 66.035 202.075 ;
        RECT 66.225 201.955 66.455 203.295 ;
        RECT 66.635 202.455 66.865 203.355 ;
        RECT 67.065 202.755 67.310 203.535 ;
        RECT 67.480 202.995 67.910 203.355 ;
        RECT 68.490 203.165 69.220 203.535 ;
        RECT 67.480 202.805 69.220 202.995 ;
        RECT 67.480 202.575 67.700 202.805 ;
        RECT 66.635 201.775 66.975 202.455 ;
        RECT 66.225 201.575 66.975 201.775 ;
        RECT 67.155 202.275 67.700 202.575 ;
        RECT 66.225 201.185 66.465 201.575 ;
        RECT 66.635 200.985 66.985 201.395 ;
        RECT 67.155 201.165 67.485 202.275 ;
        RECT 67.870 202.005 68.295 202.625 ;
        RECT 68.490 202.005 68.750 202.625 ;
        RECT 68.960 202.295 69.220 202.805 ;
        RECT 67.655 201.635 68.680 201.835 ;
        RECT 67.655 201.165 67.835 201.635 ;
        RECT 68.005 200.985 68.335 201.465 ;
        RECT 68.510 201.165 68.680 201.635 ;
        RECT 68.945 200.985 69.230 202.125 ;
        RECT 69.420 201.165 69.700 203.355 ;
        RECT 69.885 202.810 70.175 203.535 ;
        RECT 70.395 202.880 70.725 203.315 ;
        RECT 70.895 202.925 71.065 203.535 ;
        RECT 70.345 202.795 70.725 202.880 ;
        RECT 71.235 202.795 71.565 203.320 ;
        RECT 71.825 203.005 72.035 203.535 ;
        RECT 72.310 203.085 73.095 203.255 ;
        RECT 73.265 203.085 73.670 203.255 ;
        RECT 70.345 202.755 70.570 202.795 ;
        RECT 70.345 202.175 70.515 202.755 ;
        RECT 71.235 202.625 71.435 202.795 ;
        RECT 72.310 202.625 72.480 203.085 ;
        RECT 70.685 202.295 71.435 202.625 ;
        RECT 71.605 202.295 72.480 202.625 ;
        RECT 69.885 200.985 70.175 202.150 ;
        RECT 70.345 202.125 70.560 202.175 ;
        RECT 70.345 202.045 70.735 202.125 ;
        RECT 70.405 201.200 70.735 202.045 ;
        RECT 71.245 202.090 71.435 202.295 ;
        RECT 70.905 200.985 71.075 201.995 ;
        RECT 71.245 201.715 72.140 202.090 ;
        RECT 71.245 201.155 71.585 201.715 ;
        RECT 71.815 200.985 72.130 201.485 ;
        RECT 72.310 201.455 72.480 202.295 ;
        RECT 72.650 202.585 73.115 202.915 ;
        RECT 73.500 202.855 73.670 203.085 ;
        RECT 73.850 203.035 74.220 203.535 ;
        RECT 74.540 203.085 75.215 203.255 ;
        RECT 75.410 203.085 75.745 203.255 ;
        RECT 72.650 201.625 72.970 202.585 ;
        RECT 73.500 202.555 74.330 202.855 ;
        RECT 73.140 201.655 73.330 202.375 ;
        RECT 73.500 201.485 73.670 202.555 ;
        RECT 74.130 202.525 74.330 202.555 ;
        RECT 73.840 202.305 74.010 202.375 ;
        RECT 74.540 202.305 74.710 203.085 ;
        RECT 75.575 202.945 75.745 203.085 ;
        RECT 75.915 203.075 76.165 203.535 ;
        RECT 73.840 202.135 74.710 202.305 ;
        RECT 74.880 202.665 75.405 202.885 ;
        RECT 75.575 202.815 75.800 202.945 ;
        RECT 73.840 202.045 74.350 202.135 ;
        RECT 72.310 201.285 73.195 201.455 ;
        RECT 73.420 201.155 73.670 201.485 ;
        RECT 73.840 200.985 74.010 201.785 ;
        RECT 74.180 201.430 74.350 202.045 ;
        RECT 74.880 201.965 75.050 202.665 ;
        RECT 74.520 201.600 75.050 201.965 ;
        RECT 75.220 201.900 75.460 202.495 ;
        RECT 75.630 201.710 75.800 202.815 ;
        RECT 75.970 201.955 76.250 202.905 ;
        RECT 75.495 201.580 75.800 201.710 ;
        RECT 74.180 201.260 75.285 201.430 ;
        RECT 75.495 201.155 75.745 201.580 ;
        RECT 75.915 200.985 76.180 201.445 ;
        RECT 76.420 201.155 76.605 203.275 ;
        RECT 76.775 203.155 77.105 203.535 ;
        RECT 77.275 202.985 77.445 203.275 ;
        RECT 76.780 202.815 77.445 202.985 ;
        RECT 77.710 202.985 77.965 203.275 ;
        RECT 78.135 203.155 78.465 203.535 ;
        RECT 77.710 202.815 78.460 202.985 ;
        RECT 76.780 201.825 77.010 202.815 ;
        RECT 77.180 201.995 77.530 202.645 ;
        RECT 77.710 201.995 78.060 202.645 ;
        RECT 78.230 201.825 78.460 202.815 ;
        RECT 76.780 201.655 77.445 201.825 ;
        RECT 76.775 200.985 77.105 201.485 ;
        RECT 77.275 201.155 77.445 201.655 ;
        RECT 77.710 201.655 78.460 201.825 ;
        RECT 77.710 201.155 77.965 201.655 ;
        RECT 78.135 200.985 78.465 201.485 ;
        RECT 78.635 201.155 78.805 203.275 ;
        RECT 79.165 203.175 79.495 203.535 ;
        RECT 79.665 203.145 80.160 203.315 ;
        RECT 80.365 203.145 81.220 203.315 ;
        RECT 79.035 201.955 79.495 203.005 ;
        RECT 78.975 201.170 79.300 201.955 ;
        RECT 79.665 201.785 79.835 203.145 ;
        RECT 80.005 202.235 80.355 202.855 ;
        RECT 80.525 202.635 80.880 202.855 ;
        RECT 80.525 202.045 80.695 202.635 ;
        RECT 81.050 202.435 81.220 203.145 ;
        RECT 82.095 203.075 82.425 203.535 ;
        RECT 82.635 203.175 82.985 203.345 ;
        RECT 81.425 202.605 82.215 202.855 ;
        RECT 82.635 202.785 82.895 203.175 ;
        RECT 83.205 203.085 84.155 203.365 ;
        RECT 84.325 203.095 84.515 203.535 ;
        RECT 84.685 203.155 85.755 203.325 ;
        RECT 82.385 202.435 82.555 202.615 ;
        RECT 79.665 201.615 80.060 201.785 ;
        RECT 80.230 201.655 80.695 202.045 ;
        RECT 80.865 202.265 82.555 202.435 ;
        RECT 79.890 201.485 80.060 201.615 ;
        RECT 80.865 201.485 81.035 202.265 ;
        RECT 82.725 202.095 82.895 202.785 ;
        RECT 81.395 201.925 82.895 202.095 ;
        RECT 83.085 202.125 83.295 202.915 ;
        RECT 83.465 202.295 83.815 202.915 ;
        RECT 83.985 202.305 84.155 203.085 ;
        RECT 84.685 202.925 84.855 203.155 ;
        RECT 84.325 202.755 84.855 202.925 ;
        RECT 84.325 202.475 84.545 202.755 ;
        RECT 85.025 202.585 85.265 202.985 ;
        RECT 83.985 202.135 84.390 202.305 ;
        RECT 84.725 202.215 85.265 202.585 ;
        RECT 85.435 202.800 85.755 203.155 ;
        RECT 86.000 203.075 86.305 203.535 ;
        RECT 86.475 202.825 86.725 203.355 ;
        RECT 85.435 202.625 85.760 202.800 ;
        RECT 85.435 202.325 86.350 202.625 ;
        RECT 85.610 202.295 86.350 202.325 ;
        RECT 83.085 201.965 83.760 202.125 ;
        RECT 84.220 202.045 84.390 202.135 ;
        RECT 83.085 201.955 84.050 201.965 ;
        RECT 82.725 201.785 82.895 201.925 ;
        RECT 79.470 200.985 79.720 201.445 ;
        RECT 79.890 201.155 80.140 201.485 ;
        RECT 80.355 201.155 81.035 201.485 ;
        RECT 81.205 201.585 82.280 201.755 ;
        RECT 82.725 201.615 83.285 201.785 ;
        RECT 83.590 201.665 84.050 201.955 ;
        RECT 84.220 201.875 85.440 202.045 ;
        RECT 81.205 201.245 81.375 201.585 ;
        RECT 81.610 200.985 81.940 201.415 ;
        RECT 82.110 201.245 82.280 201.585 ;
        RECT 82.575 200.985 82.945 201.445 ;
        RECT 83.115 201.155 83.285 201.615 ;
        RECT 84.220 201.495 84.390 201.875 ;
        RECT 85.610 201.705 85.780 202.295 ;
        RECT 86.520 202.175 86.725 202.825 ;
        RECT 86.895 202.780 87.145 203.535 ;
        RECT 87.405 202.715 87.635 203.535 ;
        RECT 87.805 202.735 88.135 203.365 ;
        RECT 87.385 202.295 87.715 202.545 ;
        RECT 83.520 201.155 84.390 201.495 ;
        RECT 84.980 201.535 85.780 201.705 ;
        RECT 84.560 200.985 84.810 201.445 ;
        RECT 84.980 201.245 85.150 201.535 ;
        RECT 85.330 200.985 85.660 201.365 ;
        RECT 86.000 200.985 86.305 202.125 ;
        RECT 86.475 201.295 86.725 202.175 ;
        RECT 87.885 202.135 88.135 202.735 ;
        RECT 88.305 202.715 88.515 203.535 ;
        RECT 88.745 202.765 90.415 203.535 ;
        RECT 91.045 202.785 92.255 203.535 ;
        RECT 88.745 202.245 89.495 202.765 ;
        RECT 86.895 200.985 87.145 202.125 ;
        RECT 87.405 200.985 87.635 202.125 ;
        RECT 87.805 201.155 88.135 202.135 ;
        RECT 88.305 200.985 88.515 202.125 ;
        RECT 89.665 202.075 90.415 202.595 ;
        RECT 88.745 200.985 90.415 202.075 ;
        RECT 91.045 202.075 91.565 202.615 ;
        RECT 91.735 202.245 92.255 202.785 ;
        RECT 91.045 200.985 92.255 202.075 ;
        RECT 18.280 200.815 92.340 200.985 ;
        RECT 18.365 199.725 19.575 200.815 ;
        RECT 19.745 200.380 25.090 200.815 ;
        RECT 25.265 200.380 30.610 200.815 ;
        RECT 18.365 199.015 18.885 199.555 ;
        RECT 19.055 199.185 19.575 199.725 ;
        RECT 18.365 198.265 19.575 199.015 ;
        RECT 21.330 198.810 21.670 199.640 ;
        RECT 23.150 199.130 23.500 200.380 ;
        RECT 26.850 198.810 27.190 199.640 ;
        RECT 28.670 199.130 29.020 200.380 ;
        RECT 31.245 199.650 31.535 200.815 ;
        RECT 31.705 200.380 37.050 200.815 ;
        RECT 19.745 198.265 25.090 198.810 ;
        RECT 25.265 198.265 30.610 198.810 ;
        RECT 31.245 198.265 31.535 198.990 ;
        RECT 33.290 198.810 33.630 199.640 ;
        RECT 35.110 199.130 35.460 200.380 ;
        RECT 37.245 200.225 37.485 200.615 ;
        RECT 37.655 200.405 38.005 200.815 ;
        RECT 37.245 200.025 37.995 200.225 ;
        RECT 31.705 198.265 37.050 198.810 ;
        RECT 37.245 198.505 37.475 199.845 ;
        RECT 37.655 199.345 37.995 200.025 ;
        RECT 38.175 199.525 38.505 200.635 ;
        RECT 38.675 200.165 38.855 200.635 ;
        RECT 39.025 200.335 39.355 200.815 ;
        RECT 39.530 200.165 39.700 200.635 ;
        RECT 38.675 199.965 39.700 200.165 ;
        RECT 37.655 198.445 37.885 199.345 ;
        RECT 38.175 199.225 38.720 199.525 ;
        RECT 38.085 198.265 38.330 199.045 ;
        RECT 38.500 198.995 38.720 199.225 ;
        RECT 38.890 199.175 39.315 199.795 ;
        RECT 39.510 199.175 39.770 199.795 ;
        RECT 39.965 199.675 40.250 200.815 ;
        RECT 39.980 198.995 40.240 199.505 ;
        RECT 38.500 198.805 40.240 198.995 ;
        RECT 38.500 198.445 38.930 198.805 ;
        RECT 39.510 198.265 40.240 198.635 ;
        RECT 40.440 198.445 40.720 200.635 ;
        RECT 40.905 200.380 46.250 200.815 ;
        RECT 42.490 198.810 42.830 199.640 ;
        RECT 44.310 199.130 44.660 200.380 ;
        RECT 47.365 200.225 47.605 200.615 ;
        RECT 47.775 200.405 48.125 200.815 ;
        RECT 47.365 200.025 48.115 200.225 ;
        RECT 40.905 198.265 46.250 198.810 ;
        RECT 47.365 198.505 47.595 199.845 ;
        RECT 47.775 199.345 48.115 200.025 ;
        RECT 48.295 199.525 48.625 200.635 ;
        RECT 48.795 200.165 48.975 200.635 ;
        RECT 49.145 200.335 49.475 200.815 ;
        RECT 49.650 200.165 49.820 200.635 ;
        RECT 48.795 199.965 49.820 200.165 ;
        RECT 47.775 198.445 48.005 199.345 ;
        RECT 48.295 199.225 48.840 199.525 ;
        RECT 48.205 198.265 48.450 199.045 ;
        RECT 48.620 198.995 48.840 199.225 ;
        RECT 49.010 199.175 49.435 199.795 ;
        RECT 49.630 199.175 49.890 199.795 ;
        RECT 50.085 199.675 50.370 200.815 ;
        RECT 50.100 198.995 50.360 199.505 ;
        RECT 48.620 198.805 50.360 198.995 ;
        RECT 48.620 198.445 49.050 198.805 ;
        RECT 49.630 198.265 50.360 198.635 ;
        RECT 50.560 198.445 50.840 200.635 ;
        RECT 51.025 200.380 56.370 200.815 ;
        RECT 52.610 198.810 52.950 199.640 ;
        RECT 54.430 199.130 54.780 200.380 ;
        RECT 57.005 199.650 57.295 200.815 ;
        RECT 58.405 200.225 58.645 200.615 ;
        RECT 58.815 200.405 59.165 200.815 ;
        RECT 58.405 200.025 59.155 200.225 ;
        RECT 51.025 198.265 56.370 198.810 ;
        RECT 57.005 198.265 57.295 198.990 ;
        RECT 58.405 198.505 58.635 199.845 ;
        RECT 58.815 199.345 59.155 200.025 ;
        RECT 59.335 199.525 59.665 200.635 ;
        RECT 59.835 200.165 60.015 200.635 ;
        RECT 60.185 200.335 60.515 200.815 ;
        RECT 60.690 200.165 60.860 200.635 ;
        RECT 59.835 199.965 60.860 200.165 ;
        RECT 58.815 198.445 59.045 199.345 ;
        RECT 59.335 199.225 59.880 199.525 ;
        RECT 59.245 198.265 59.490 199.045 ;
        RECT 59.660 198.995 59.880 199.225 ;
        RECT 60.050 199.175 60.475 199.795 ;
        RECT 60.670 199.175 60.930 199.795 ;
        RECT 61.125 199.675 61.410 200.815 ;
        RECT 61.140 198.995 61.400 199.505 ;
        RECT 59.660 198.805 61.400 198.995 ;
        RECT 59.660 198.445 60.090 198.805 ;
        RECT 60.670 198.265 61.400 198.635 ;
        RECT 61.600 198.445 61.880 200.635 ;
        RECT 62.065 200.380 67.410 200.815 ;
        RECT 63.650 198.810 63.990 199.640 ;
        RECT 65.470 199.130 65.820 200.380 ;
        RECT 67.585 199.675 67.860 200.645 ;
        RECT 68.070 200.015 68.350 200.815 ;
        RECT 68.520 200.305 70.135 200.635 ;
        RECT 68.520 199.965 69.695 200.135 ;
        RECT 68.520 199.845 68.690 199.965 ;
        RECT 68.030 199.675 68.690 199.845 ;
        RECT 67.585 198.940 67.755 199.675 ;
        RECT 68.030 199.505 68.200 199.675 ;
        RECT 68.950 199.505 69.195 199.795 ;
        RECT 69.365 199.675 69.695 199.965 ;
        RECT 69.955 199.505 70.125 200.065 ;
        RECT 70.375 199.675 70.635 200.815 ;
        RECT 71.320 199.945 71.605 200.815 ;
        RECT 71.775 200.185 72.035 200.645 ;
        RECT 72.210 200.355 72.465 200.815 ;
        RECT 72.635 200.185 72.895 200.645 ;
        RECT 71.775 200.015 72.895 200.185 ;
        RECT 73.065 200.015 73.375 200.815 ;
        RECT 71.775 199.765 72.035 200.015 ;
        RECT 73.545 199.845 73.855 200.645 ;
        RECT 71.280 199.595 72.035 199.765 ;
        RECT 72.825 199.675 73.855 199.845 ;
        RECT 74.945 199.675 75.225 200.815 ;
        RECT 67.925 199.175 68.200 199.505 ;
        RECT 68.370 199.175 69.195 199.505 ;
        RECT 69.410 199.175 70.125 199.505 ;
        RECT 70.295 199.255 70.630 199.505 ;
        RECT 68.030 199.005 68.200 199.175 ;
        RECT 69.875 199.085 70.125 199.175 ;
        RECT 71.280 199.085 71.685 199.595 ;
        RECT 72.825 199.425 72.995 199.675 ;
        RECT 71.855 199.255 72.995 199.425 ;
        RECT 62.065 198.265 67.410 198.810 ;
        RECT 67.585 198.595 67.860 198.940 ;
        RECT 68.030 198.835 69.695 199.005 ;
        RECT 68.050 198.265 68.425 198.665 ;
        RECT 68.595 198.485 68.765 198.835 ;
        RECT 68.935 198.265 69.265 198.665 ;
        RECT 69.435 198.435 69.695 198.835 ;
        RECT 69.875 198.665 70.205 199.085 ;
        RECT 70.375 198.265 70.635 199.085 ;
        RECT 71.280 198.915 72.930 199.085 ;
        RECT 73.165 198.935 73.515 199.505 ;
        RECT 71.325 198.265 71.605 198.745 ;
        RECT 71.775 198.525 72.035 198.915 ;
        RECT 72.210 198.265 72.465 198.745 ;
        RECT 72.635 198.525 72.930 198.915 ;
        RECT 73.685 198.765 73.855 199.675 ;
        RECT 75.395 199.665 75.725 200.645 ;
        RECT 75.895 199.675 76.155 200.815 ;
        RECT 76.335 199.675 76.665 200.815 ;
        RECT 77.195 199.845 77.525 200.630 ;
        RECT 76.845 199.675 77.525 199.845 ;
        RECT 78.635 200.205 78.965 200.635 ;
        RECT 79.145 200.375 79.340 200.815 ;
        RECT 79.510 200.205 79.840 200.635 ;
        RECT 78.635 200.035 79.840 200.205 ;
        RECT 78.635 199.705 79.530 200.035 ;
        RECT 80.010 199.865 80.285 200.635 ;
        RECT 79.700 199.675 80.285 199.865 ;
        RECT 80.465 199.725 82.135 200.815 ;
        RECT 74.955 199.235 75.290 199.505 ;
        RECT 75.460 199.115 75.630 199.665 ;
        RECT 75.800 199.255 76.135 199.505 ;
        RECT 76.325 199.255 76.675 199.505 ;
        RECT 75.460 199.065 75.635 199.115 ;
        RECT 76.845 199.075 77.015 199.675 ;
        RECT 77.185 199.255 77.535 199.505 ;
        RECT 78.640 199.175 78.935 199.505 ;
        RECT 79.115 199.175 79.530 199.505 ;
        RECT 73.110 198.265 73.385 198.745 ;
        RECT 73.555 198.435 73.855 198.765 ;
        RECT 74.945 198.265 75.255 199.065 ;
        RECT 75.460 198.435 76.155 199.065 ;
        RECT 76.335 198.265 76.605 199.075 ;
        RECT 76.775 198.435 77.105 199.075 ;
        RECT 77.275 198.265 77.515 199.075 ;
        RECT 78.635 198.265 78.935 198.995 ;
        RECT 79.115 198.555 79.345 199.175 ;
        RECT 79.700 199.005 79.875 199.675 ;
        RECT 79.545 198.825 79.875 199.005 ;
        RECT 80.045 198.855 80.285 199.505 ;
        RECT 80.465 199.035 81.215 199.555 ;
        RECT 81.385 199.205 82.135 199.725 ;
        RECT 82.765 199.650 83.055 200.815 ;
        RECT 83.225 199.725 84.435 200.815 ;
        RECT 79.545 198.445 79.770 198.825 ;
        RECT 79.940 198.265 80.270 198.655 ;
        RECT 80.465 198.265 82.135 199.035 ;
        RECT 83.225 199.015 83.745 199.555 ;
        RECT 83.915 199.185 84.435 199.725 ;
        RECT 84.605 199.675 84.990 200.645 ;
        RECT 85.160 200.355 85.485 200.815 ;
        RECT 86.005 200.185 86.285 200.645 ;
        RECT 85.160 199.965 86.285 200.185 ;
        RECT 82.765 198.265 83.055 198.990 ;
        RECT 83.225 198.265 84.435 199.015 ;
        RECT 84.605 199.005 84.885 199.675 ;
        RECT 85.160 199.505 85.610 199.965 ;
        RECT 86.475 199.795 86.875 200.645 ;
        RECT 87.275 200.355 87.545 200.815 ;
        RECT 87.715 200.185 88.000 200.645 ;
        RECT 85.055 199.175 85.610 199.505 ;
        RECT 85.780 199.235 86.875 199.795 ;
        RECT 85.160 199.065 85.610 199.175 ;
        RECT 84.605 198.435 84.990 199.005 ;
        RECT 85.160 198.895 86.285 199.065 ;
        RECT 85.160 198.265 85.485 198.725 ;
        RECT 86.005 198.435 86.285 198.895 ;
        RECT 86.475 198.435 86.875 199.235 ;
        RECT 87.045 199.965 88.000 200.185 ;
        RECT 87.045 199.065 87.255 199.965 ;
        RECT 87.425 199.235 88.115 199.795 ;
        RECT 88.325 199.675 88.555 200.815 ;
        RECT 88.725 199.665 89.055 200.645 ;
        RECT 89.225 199.675 89.435 200.815 ;
        RECT 89.665 199.725 90.875 200.815 ;
        RECT 88.305 199.255 88.635 199.505 ;
        RECT 87.045 198.895 88.000 199.065 ;
        RECT 87.275 198.265 87.545 198.725 ;
        RECT 87.715 198.435 88.000 198.895 ;
        RECT 88.325 198.265 88.555 199.085 ;
        RECT 88.805 199.065 89.055 199.665 ;
        RECT 88.725 198.435 89.055 199.065 ;
        RECT 89.225 198.265 89.435 199.085 ;
        RECT 89.665 199.015 90.185 199.555 ;
        RECT 90.355 199.185 90.875 199.725 ;
        RECT 91.045 199.725 92.255 200.815 ;
        RECT 91.045 199.185 91.565 199.725 ;
        RECT 91.735 199.015 92.255 199.555 ;
        RECT 89.665 198.265 90.875 199.015 ;
        RECT 91.045 198.265 92.255 199.015 ;
        RECT 18.280 198.095 92.340 198.265 ;
        RECT 18.365 197.345 19.575 198.095 ;
        RECT 19.745 197.550 25.090 198.095 ;
        RECT 25.265 197.550 30.610 198.095 ;
        RECT 18.365 196.805 18.885 197.345 ;
        RECT 19.055 196.635 19.575 197.175 ;
        RECT 21.330 196.720 21.670 197.550 ;
        RECT 18.365 195.545 19.575 196.635 ;
        RECT 23.150 195.980 23.500 197.230 ;
        RECT 26.850 196.720 27.190 197.550 ;
        RECT 30.785 197.325 34.295 198.095 ;
        RECT 28.670 195.980 29.020 197.230 ;
        RECT 30.785 196.805 32.435 197.325 ;
        RECT 32.605 196.635 34.295 197.155 ;
        RECT 19.745 195.545 25.090 195.980 ;
        RECT 25.265 195.545 30.610 195.980 ;
        RECT 30.785 195.545 34.295 196.635 ;
        RECT 34.945 196.515 35.175 197.855 ;
        RECT 35.355 197.015 35.585 197.915 ;
        RECT 35.785 197.315 36.030 198.095 ;
        RECT 36.200 197.555 36.630 197.915 ;
        RECT 37.210 197.725 37.940 198.095 ;
        RECT 36.200 197.365 37.940 197.555 ;
        RECT 36.200 197.135 36.420 197.365 ;
        RECT 35.355 196.335 35.695 197.015 ;
        RECT 34.945 196.135 35.695 196.335 ;
        RECT 35.875 196.835 36.420 197.135 ;
        RECT 34.945 195.745 35.185 196.135 ;
        RECT 35.355 195.545 35.705 195.955 ;
        RECT 35.875 195.725 36.205 196.835 ;
        RECT 36.590 196.565 37.015 197.185 ;
        RECT 37.210 196.565 37.470 197.185 ;
        RECT 37.680 196.855 37.940 197.365 ;
        RECT 36.375 196.195 37.400 196.395 ;
        RECT 36.375 195.725 36.555 196.195 ;
        RECT 36.725 195.545 37.055 196.025 ;
        RECT 37.230 195.725 37.400 196.195 ;
        RECT 37.665 195.545 37.950 196.685 ;
        RECT 38.140 195.725 38.420 197.915 ;
        RECT 38.605 197.550 43.950 198.095 ;
        RECT 40.190 196.720 40.530 197.550 ;
        RECT 44.125 197.370 44.415 198.095 ;
        RECT 42.010 195.980 42.360 197.230 ;
        RECT 38.605 195.545 43.950 195.980 ;
        RECT 44.125 195.545 44.415 196.710 ;
        RECT 44.600 195.725 44.880 197.915 ;
        RECT 45.080 197.725 45.810 198.095 ;
        RECT 46.390 197.555 46.820 197.915 ;
        RECT 45.080 197.365 46.820 197.555 ;
        RECT 45.080 196.855 45.340 197.365 ;
        RECT 45.070 195.545 45.355 196.685 ;
        RECT 45.550 196.565 45.810 197.185 ;
        RECT 46.005 196.565 46.430 197.185 ;
        RECT 46.600 197.135 46.820 197.365 ;
        RECT 46.990 197.315 47.235 198.095 ;
        RECT 46.600 196.835 47.145 197.135 ;
        RECT 47.435 197.015 47.665 197.915 ;
        RECT 45.620 196.195 46.645 196.395 ;
        RECT 45.620 195.725 45.790 196.195 ;
        RECT 45.965 195.545 46.295 196.025 ;
        RECT 46.465 195.725 46.645 196.195 ;
        RECT 46.815 195.725 47.145 196.835 ;
        RECT 47.325 196.335 47.665 197.015 ;
        RECT 47.845 196.515 48.075 197.855 ;
        RECT 48.265 197.325 50.855 198.095 ;
        RECT 51.535 197.440 51.865 197.875 ;
        RECT 52.035 197.485 52.205 198.095 ;
        RECT 51.485 197.355 51.865 197.440 ;
        RECT 52.375 197.355 52.705 197.880 ;
        RECT 52.965 197.565 53.175 198.095 ;
        RECT 53.450 197.645 54.235 197.815 ;
        RECT 54.405 197.645 54.810 197.815 ;
        RECT 48.265 196.805 49.475 197.325 ;
        RECT 51.485 197.315 51.710 197.355 ;
        RECT 49.645 196.635 50.855 197.155 ;
        RECT 47.325 196.135 48.075 196.335 ;
        RECT 47.315 195.545 47.665 195.955 ;
        RECT 47.835 195.745 48.075 196.135 ;
        RECT 48.265 195.545 50.855 196.635 ;
        RECT 51.485 196.735 51.655 197.315 ;
        RECT 52.375 197.185 52.575 197.355 ;
        RECT 53.450 197.185 53.620 197.645 ;
        RECT 51.825 196.855 52.575 197.185 ;
        RECT 52.745 196.855 53.620 197.185 ;
        RECT 51.485 196.685 51.700 196.735 ;
        RECT 51.485 196.605 51.875 196.685 ;
        RECT 51.545 195.760 51.875 196.605 ;
        RECT 52.385 196.650 52.575 196.855 ;
        RECT 52.045 195.545 52.215 196.555 ;
        RECT 52.385 196.275 53.280 196.650 ;
        RECT 52.385 195.715 52.725 196.275 ;
        RECT 52.955 195.545 53.270 196.045 ;
        RECT 53.450 196.015 53.620 196.855 ;
        RECT 53.790 197.145 54.255 197.475 ;
        RECT 54.640 197.415 54.810 197.645 ;
        RECT 54.990 197.595 55.360 198.095 ;
        RECT 55.680 197.645 56.355 197.815 ;
        RECT 56.550 197.645 56.885 197.815 ;
        RECT 53.790 196.185 54.110 197.145 ;
        RECT 54.640 197.115 55.470 197.415 ;
        RECT 54.280 196.215 54.470 196.935 ;
        RECT 54.640 196.045 54.810 197.115 ;
        RECT 55.270 197.085 55.470 197.115 ;
        RECT 54.980 196.865 55.150 196.935 ;
        RECT 55.680 196.865 55.850 197.645 ;
        RECT 56.715 197.505 56.885 197.645 ;
        RECT 57.055 197.635 57.305 198.095 ;
        RECT 54.980 196.695 55.850 196.865 ;
        RECT 56.020 197.225 56.545 197.445 ;
        RECT 56.715 197.375 56.940 197.505 ;
        RECT 54.980 196.605 55.490 196.695 ;
        RECT 53.450 195.845 54.335 196.015 ;
        RECT 54.560 195.715 54.810 196.045 ;
        RECT 54.980 195.545 55.150 196.345 ;
        RECT 55.320 195.990 55.490 196.605 ;
        RECT 56.020 196.525 56.190 197.225 ;
        RECT 55.660 196.160 56.190 196.525 ;
        RECT 56.360 196.460 56.600 197.055 ;
        RECT 56.770 196.270 56.940 197.375 ;
        RECT 57.110 196.515 57.390 197.465 ;
        RECT 56.635 196.140 56.940 196.270 ;
        RECT 55.320 195.820 56.425 195.990 ;
        RECT 56.635 195.715 56.885 196.140 ;
        RECT 57.055 195.545 57.320 196.005 ;
        RECT 57.560 195.715 57.745 197.835 ;
        RECT 57.915 197.715 58.245 198.095 ;
        RECT 58.415 197.545 58.585 197.835 ;
        RECT 57.920 197.375 58.585 197.545 ;
        RECT 57.920 196.385 58.150 197.375 ;
        RECT 58.845 197.325 60.515 198.095 ;
        RECT 60.775 197.545 60.945 197.835 ;
        RECT 61.115 197.715 61.445 198.095 ;
        RECT 60.775 197.375 61.440 197.545 ;
        RECT 58.320 196.555 58.670 197.205 ;
        RECT 58.845 196.805 59.595 197.325 ;
        RECT 59.765 196.635 60.515 197.155 ;
        RECT 57.920 196.215 58.585 196.385 ;
        RECT 57.915 195.545 58.245 196.045 ;
        RECT 58.415 195.715 58.585 196.215 ;
        RECT 58.845 195.545 60.515 196.635 ;
        RECT 60.690 196.555 61.040 197.205 ;
        RECT 61.210 196.385 61.440 197.375 ;
        RECT 60.775 196.215 61.440 196.385 ;
        RECT 60.775 195.715 60.945 196.215 ;
        RECT 61.115 195.545 61.445 196.045 ;
        RECT 61.615 195.715 61.800 197.835 ;
        RECT 62.055 197.635 62.305 198.095 ;
        RECT 62.475 197.645 62.810 197.815 ;
        RECT 63.005 197.645 63.680 197.815 ;
        RECT 62.475 197.505 62.645 197.645 ;
        RECT 61.970 196.515 62.250 197.465 ;
        RECT 62.420 197.375 62.645 197.505 ;
        RECT 62.420 196.270 62.590 197.375 ;
        RECT 62.815 197.225 63.340 197.445 ;
        RECT 62.760 196.460 63.000 197.055 ;
        RECT 63.170 196.525 63.340 197.225 ;
        RECT 63.510 196.865 63.680 197.645 ;
        RECT 64.000 197.595 64.370 198.095 ;
        RECT 64.550 197.645 64.955 197.815 ;
        RECT 65.125 197.645 65.910 197.815 ;
        RECT 64.550 197.415 64.720 197.645 ;
        RECT 63.890 197.115 64.720 197.415 ;
        RECT 65.105 197.145 65.570 197.475 ;
        RECT 63.890 197.085 64.090 197.115 ;
        RECT 64.210 196.865 64.380 196.935 ;
        RECT 63.510 196.695 64.380 196.865 ;
        RECT 63.870 196.605 64.380 196.695 ;
        RECT 62.420 196.140 62.725 196.270 ;
        RECT 63.170 196.160 63.700 196.525 ;
        RECT 62.040 195.545 62.305 196.005 ;
        RECT 62.475 195.715 62.725 196.140 ;
        RECT 63.870 195.990 64.040 196.605 ;
        RECT 62.935 195.820 64.040 195.990 ;
        RECT 64.210 195.545 64.380 196.345 ;
        RECT 64.550 196.045 64.720 197.115 ;
        RECT 64.890 196.215 65.080 196.935 ;
        RECT 65.250 196.185 65.570 197.145 ;
        RECT 65.740 197.185 65.910 197.645 ;
        RECT 66.185 197.565 66.395 198.095 ;
        RECT 66.655 197.355 66.985 197.880 ;
        RECT 67.155 197.485 67.325 198.095 ;
        RECT 67.495 197.440 67.825 197.875 ;
        RECT 67.495 197.355 67.875 197.440 ;
        RECT 66.785 197.185 66.985 197.355 ;
        RECT 67.650 197.315 67.875 197.355 ;
        RECT 65.740 196.855 66.615 197.185 ;
        RECT 66.785 196.855 67.535 197.185 ;
        RECT 64.550 195.715 64.800 196.045 ;
        RECT 65.740 196.015 65.910 196.855 ;
        RECT 66.785 196.650 66.975 196.855 ;
        RECT 67.705 196.735 67.875 197.315 ;
        RECT 68.045 197.325 69.715 198.095 ;
        RECT 69.885 197.370 70.175 198.095 ;
        RECT 70.345 197.325 72.935 198.095 ;
        RECT 73.115 197.375 73.445 198.095 ;
        RECT 73.990 197.695 75.605 197.865 ;
        RECT 75.775 197.695 76.105 198.095 ;
        RECT 75.435 197.525 75.605 197.695 ;
        RECT 76.275 197.620 76.610 197.880 ;
        RECT 68.045 196.805 68.795 197.325 ;
        RECT 67.660 196.685 67.875 196.735 ;
        RECT 66.080 196.275 66.975 196.650 ;
        RECT 67.485 196.605 67.875 196.685 ;
        RECT 68.965 196.635 69.715 197.155 ;
        RECT 70.345 196.805 71.555 197.325 ;
        RECT 65.025 195.845 65.910 196.015 ;
        RECT 66.090 195.545 66.405 196.045 ;
        RECT 66.635 195.715 66.975 196.275 ;
        RECT 67.145 195.545 67.315 196.555 ;
        RECT 67.485 195.760 67.815 196.605 ;
        RECT 68.045 195.545 69.715 196.635 ;
        RECT 69.885 195.545 70.175 196.710 ;
        RECT 71.725 196.635 72.935 197.155 ;
        RECT 73.170 196.855 73.520 197.185 ;
        RECT 73.830 196.855 74.250 197.520 ;
        RECT 74.420 197.075 74.710 197.515 ;
        RECT 74.900 197.075 75.170 197.515 ;
        RECT 75.435 197.355 75.995 197.525 ;
        RECT 75.825 197.185 75.995 197.355 ;
        RECT 75.380 197.075 75.630 197.185 ;
        RECT 74.420 196.905 74.715 197.075 ;
        RECT 74.900 196.905 75.175 197.075 ;
        RECT 75.380 196.905 75.635 197.075 ;
        RECT 74.420 196.855 74.710 196.905 ;
        RECT 74.900 196.855 75.170 196.905 ;
        RECT 75.380 196.855 75.630 196.905 ;
        RECT 75.825 196.855 76.130 197.185 ;
        RECT 73.170 196.735 73.375 196.855 ;
        RECT 70.345 195.545 72.935 196.635 ;
        RECT 73.165 196.565 73.375 196.735 ;
        RECT 75.825 196.685 75.995 196.855 ;
        RECT 73.625 196.515 75.995 196.685 ;
        RECT 73.195 195.885 73.365 196.385 ;
        RECT 73.625 196.055 73.795 196.515 ;
        RECT 74.025 196.135 75.450 196.305 ;
        RECT 74.025 195.885 74.355 196.135 ;
        RECT 73.195 195.715 74.355 195.885 ;
        RECT 74.580 195.545 74.910 195.965 ;
        RECT 75.165 195.715 75.450 196.135 ;
        RECT 75.695 195.545 76.025 196.345 ;
        RECT 76.355 196.265 76.610 197.620 ;
        RECT 77.710 197.565 78.000 197.915 ;
        RECT 78.195 197.735 78.525 198.095 ;
        RECT 78.695 197.565 78.925 197.870 ;
        RECT 77.710 197.395 78.925 197.565 ;
        RECT 79.115 197.755 79.285 197.790 ;
        RECT 79.115 197.585 79.315 197.755 ;
        RECT 79.115 197.225 79.285 197.585 ;
        RECT 77.770 197.075 78.030 197.185 ;
        RECT 77.765 196.905 78.030 197.075 ;
        RECT 77.770 196.855 78.030 196.905 ;
        RECT 78.210 196.855 78.595 197.185 ;
        RECT 78.765 197.055 79.285 197.225 ;
        RECT 79.545 197.325 82.135 198.095 ;
        RECT 82.395 197.545 82.565 197.835 ;
        RECT 82.735 197.715 83.065 198.095 ;
        RECT 82.395 197.375 83.060 197.545 ;
        RECT 76.275 195.755 76.610 196.265 ;
        RECT 77.710 195.545 78.030 196.685 ;
        RECT 78.210 195.805 78.405 196.855 ;
        RECT 78.765 196.675 78.935 197.055 ;
        RECT 78.585 196.395 78.935 196.675 ;
        RECT 79.125 196.525 79.370 196.885 ;
        RECT 79.545 196.805 80.755 197.325 ;
        RECT 80.925 196.635 82.135 197.155 ;
        RECT 78.585 195.715 78.915 196.395 ;
        RECT 79.115 195.545 79.370 196.345 ;
        RECT 79.545 195.545 82.135 196.635 ;
        RECT 82.310 196.555 82.660 197.205 ;
        RECT 82.830 196.385 83.060 197.375 ;
        RECT 82.395 196.215 83.060 196.385 ;
        RECT 82.395 195.715 82.565 196.215 ;
        RECT 82.735 195.545 83.065 196.045 ;
        RECT 83.235 195.715 83.460 197.835 ;
        RECT 83.675 197.635 83.925 198.095 ;
        RECT 84.110 197.645 84.440 197.815 ;
        RECT 84.620 197.645 85.370 197.815 ;
        RECT 83.660 196.515 83.940 197.115 ;
        RECT 84.110 196.115 84.280 197.645 ;
        RECT 84.450 197.145 85.030 197.475 ;
        RECT 84.450 196.275 84.690 197.145 ;
        RECT 85.200 196.865 85.370 197.645 ;
        RECT 85.620 197.595 85.990 198.095 ;
        RECT 86.170 197.645 86.630 197.815 ;
        RECT 86.860 197.645 87.530 197.815 ;
        RECT 86.170 197.415 86.340 197.645 ;
        RECT 85.540 197.115 86.340 197.415 ;
        RECT 86.510 197.145 87.060 197.475 ;
        RECT 85.540 197.085 85.710 197.115 ;
        RECT 85.830 196.865 86.000 196.935 ;
        RECT 85.200 196.695 86.000 196.865 ;
        RECT 85.490 196.605 86.000 196.695 ;
        RECT 84.880 196.170 85.320 196.525 ;
        RECT 83.660 195.545 83.925 196.005 ;
        RECT 84.110 195.740 84.345 196.115 ;
        RECT 85.490 195.990 85.660 196.605 ;
        RECT 84.590 195.820 85.660 195.990 ;
        RECT 85.830 195.545 86.000 196.345 ;
        RECT 86.170 196.045 86.340 197.115 ;
        RECT 86.510 196.215 86.700 196.935 ;
        RECT 86.870 196.605 87.060 197.145 ;
        RECT 87.360 197.105 87.530 197.645 ;
        RECT 87.845 197.565 88.015 198.095 ;
        RECT 88.310 197.445 88.670 197.885 ;
        RECT 88.845 197.615 89.015 198.095 ;
        RECT 89.205 197.450 89.540 197.875 ;
        RECT 89.715 197.620 89.885 198.095 ;
        RECT 90.060 197.450 90.395 197.875 ;
        RECT 90.565 197.620 90.735 198.095 ;
        RECT 88.310 197.275 88.810 197.445 ;
        RECT 89.205 197.280 90.875 197.450 ;
        RECT 91.045 197.345 92.255 198.095 ;
        RECT 88.640 197.105 88.810 197.275 ;
        RECT 87.360 196.935 88.450 197.105 ;
        RECT 88.640 196.935 90.460 197.105 ;
        RECT 86.870 196.275 87.190 196.605 ;
        RECT 86.170 195.715 86.420 196.045 ;
        RECT 87.360 196.015 87.530 196.935 ;
        RECT 88.640 196.680 88.810 196.935 ;
        RECT 90.630 196.715 90.875 197.280 ;
        RECT 87.700 196.510 88.810 196.680 ;
        RECT 89.205 196.545 90.875 196.715 ;
        RECT 91.045 196.635 91.565 197.175 ;
        RECT 91.735 196.805 92.255 197.345 ;
        RECT 87.700 196.350 88.560 196.510 ;
        RECT 86.645 195.845 87.530 196.015 ;
        RECT 87.710 195.545 87.925 196.045 ;
        RECT 88.390 195.725 88.560 196.350 ;
        RECT 88.845 195.545 89.025 196.325 ;
        RECT 89.205 195.785 89.540 196.545 ;
        RECT 89.720 195.545 89.890 196.375 ;
        RECT 90.060 195.785 90.390 196.545 ;
        RECT 90.560 195.545 90.730 196.375 ;
        RECT 91.045 195.545 92.255 196.635 ;
        RECT 18.280 195.375 92.340 195.545 ;
        RECT 18.365 194.285 19.575 195.375 ;
        RECT 19.745 194.940 25.090 195.375 ;
        RECT 25.265 194.940 30.610 195.375 ;
        RECT 18.365 193.575 18.885 194.115 ;
        RECT 19.055 193.745 19.575 194.285 ;
        RECT 18.365 192.825 19.575 193.575 ;
        RECT 21.330 193.370 21.670 194.200 ;
        RECT 23.150 193.690 23.500 194.940 ;
        RECT 26.850 193.370 27.190 194.200 ;
        RECT 28.670 193.690 29.020 194.940 ;
        RECT 31.245 194.210 31.535 195.375 ;
        RECT 31.765 194.315 32.095 195.160 ;
        RECT 32.265 194.365 32.435 195.375 ;
        RECT 32.605 194.645 32.945 195.205 ;
        RECT 33.175 194.875 33.490 195.375 ;
        RECT 33.670 194.905 34.555 195.075 ;
        RECT 31.705 194.235 32.095 194.315 ;
        RECT 32.605 194.270 33.500 194.645 ;
        RECT 31.705 194.185 31.920 194.235 ;
        RECT 31.705 193.605 31.875 194.185 ;
        RECT 32.605 194.065 32.795 194.270 ;
        RECT 33.670 194.065 33.840 194.905 ;
        RECT 34.780 194.875 35.030 195.205 ;
        RECT 32.045 193.735 32.795 194.065 ;
        RECT 32.965 193.735 33.840 194.065 ;
        RECT 31.705 193.565 31.930 193.605 ;
        RECT 32.595 193.565 32.795 193.735 ;
        RECT 19.745 192.825 25.090 193.370 ;
        RECT 25.265 192.825 30.610 193.370 ;
        RECT 31.245 192.825 31.535 193.550 ;
        RECT 31.705 193.480 32.085 193.565 ;
        RECT 31.755 193.045 32.085 193.480 ;
        RECT 32.255 192.825 32.425 193.435 ;
        RECT 32.595 193.040 32.925 193.565 ;
        RECT 33.185 192.825 33.395 193.355 ;
        RECT 33.670 193.275 33.840 193.735 ;
        RECT 34.010 193.775 34.330 194.735 ;
        RECT 34.500 193.985 34.690 194.705 ;
        RECT 34.860 193.805 35.030 194.875 ;
        RECT 35.200 194.575 35.370 195.375 ;
        RECT 35.540 194.930 36.645 195.100 ;
        RECT 35.540 194.315 35.710 194.930 ;
        RECT 36.855 194.780 37.105 195.205 ;
        RECT 37.275 194.915 37.540 195.375 ;
        RECT 35.880 194.395 36.410 194.760 ;
        RECT 36.855 194.650 37.160 194.780 ;
        RECT 35.200 194.225 35.710 194.315 ;
        RECT 35.200 194.055 36.070 194.225 ;
        RECT 35.200 193.985 35.370 194.055 ;
        RECT 35.490 193.805 35.690 193.835 ;
        RECT 34.010 193.445 34.475 193.775 ;
        RECT 34.860 193.505 35.690 193.805 ;
        RECT 34.860 193.275 35.030 193.505 ;
        RECT 33.670 193.105 34.455 193.275 ;
        RECT 34.625 193.105 35.030 193.275 ;
        RECT 35.210 192.825 35.580 193.325 ;
        RECT 35.900 193.275 36.070 194.055 ;
        RECT 36.240 193.695 36.410 194.395 ;
        RECT 36.580 193.865 36.820 194.460 ;
        RECT 36.240 193.475 36.765 193.695 ;
        RECT 36.990 193.545 37.160 194.650 ;
        RECT 36.935 193.415 37.160 193.545 ;
        RECT 37.330 193.455 37.610 194.405 ;
        RECT 36.935 193.275 37.105 193.415 ;
        RECT 35.900 193.105 36.575 193.275 ;
        RECT 36.770 193.105 37.105 193.275 ;
        RECT 37.275 192.825 37.525 193.285 ;
        RECT 37.780 193.085 37.965 195.205 ;
        RECT 38.135 194.875 38.465 195.375 ;
        RECT 38.635 194.705 38.805 195.205 ;
        RECT 38.140 194.535 38.805 194.705 ;
        RECT 38.140 193.545 38.370 194.535 ;
        RECT 38.540 193.715 38.890 194.365 ;
        RECT 39.065 194.285 41.655 195.375 ;
        RECT 41.915 194.705 42.085 195.205 ;
        RECT 42.255 194.875 42.585 195.375 ;
        RECT 41.915 194.535 42.580 194.705 ;
        RECT 39.065 193.595 40.275 194.115 ;
        RECT 40.445 193.765 41.655 194.285 ;
        RECT 41.830 193.715 42.180 194.365 ;
        RECT 38.140 193.375 38.805 193.545 ;
        RECT 38.135 192.825 38.465 193.205 ;
        RECT 38.635 193.085 38.805 193.375 ;
        RECT 39.065 192.825 41.655 193.595 ;
        RECT 42.350 193.545 42.580 194.535 ;
        RECT 41.915 193.375 42.580 193.545 ;
        RECT 41.915 193.085 42.085 193.375 ;
        RECT 42.255 192.825 42.585 193.205 ;
        RECT 42.755 193.085 42.940 195.205 ;
        RECT 43.180 194.915 43.445 195.375 ;
        RECT 43.615 194.780 43.865 195.205 ;
        RECT 44.075 194.930 45.180 195.100 ;
        RECT 43.560 194.650 43.865 194.780 ;
        RECT 43.110 193.455 43.390 194.405 ;
        RECT 43.560 193.545 43.730 194.650 ;
        RECT 43.900 193.865 44.140 194.460 ;
        RECT 44.310 194.395 44.840 194.760 ;
        RECT 44.310 193.695 44.480 194.395 ;
        RECT 45.010 194.315 45.180 194.930 ;
        RECT 45.350 194.575 45.520 195.375 ;
        RECT 45.690 194.875 45.940 195.205 ;
        RECT 46.165 194.905 47.050 195.075 ;
        RECT 45.010 194.225 45.520 194.315 ;
        RECT 43.560 193.415 43.785 193.545 ;
        RECT 43.955 193.475 44.480 193.695 ;
        RECT 44.650 194.055 45.520 194.225 ;
        RECT 43.195 192.825 43.445 193.285 ;
        RECT 43.615 193.275 43.785 193.415 ;
        RECT 44.650 193.275 44.820 194.055 ;
        RECT 45.350 193.985 45.520 194.055 ;
        RECT 45.030 193.805 45.230 193.835 ;
        RECT 45.690 193.805 45.860 194.875 ;
        RECT 46.030 193.985 46.220 194.705 ;
        RECT 45.030 193.505 45.860 193.805 ;
        RECT 46.390 193.775 46.710 194.735 ;
        RECT 43.615 193.105 43.950 193.275 ;
        RECT 44.145 193.105 44.820 193.275 ;
        RECT 45.140 192.825 45.510 193.325 ;
        RECT 45.690 193.275 45.860 193.505 ;
        RECT 46.245 193.445 46.710 193.775 ;
        RECT 46.880 194.065 47.050 194.905 ;
        RECT 47.230 194.875 47.545 195.375 ;
        RECT 47.775 194.645 48.115 195.205 ;
        RECT 47.220 194.270 48.115 194.645 ;
        RECT 48.285 194.365 48.455 195.375 ;
        RECT 47.925 194.065 48.115 194.270 ;
        RECT 48.625 194.315 48.955 195.160 ;
        RECT 48.625 194.235 49.015 194.315 ;
        RECT 48.800 194.185 49.015 194.235 ;
        RECT 46.880 193.735 47.755 194.065 ;
        RECT 47.925 193.735 48.675 194.065 ;
        RECT 46.880 193.275 47.050 193.735 ;
        RECT 47.925 193.565 48.125 193.735 ;
        RECT 48.845 193.605 49.015 194.185 ;
        RECT 48.790 193.565 49.015 193.605 ;
        RECT 45.690 193.105 46.095 193.275 ;
        RECT 46.265 193.105 47.050 193.275 ;
        RECT 47.325 192.825 47.535 193.355 ;
        RECT 47.795 193.040 48.125 193.565 ;
        RECT 48.635 193.480 49.015 193.565 ;
        RECT 49.190 194.235 49.465 195.205 ;
        RECT 49.675 194.575 49.955 195.375 ;
        RECT 50.125 194.865 51.315 195.155 ;
        RECT 50.125 194.525 51.295 194.695 ;
        RECT 50.125 194.405 50.295 194.525 ;
        RECT 49.635 194.235 50.295 194.405 ;
        RECT 49.190 193.500 49.360 194.235 ;
        RECT 49.635 194.065 49.805 194.235 ;
        RECT 50.605 194.065 50.800 194.355 ;
        RECT 50.970 194.235 51.295 194.525 ;
        RECT 51.525 194.235 51.755 195.375 ;
        RECT 51.925 194.225 52.255 195.205 ;
        RECT 52.425 194.235 52.635 195.375 ;
        RECT 53.785 194.235 54.045 195.375 ;
        RECT 54.285 194.865 55.900 195.195 ;
        RECT 49.530 193.735 49.805 194.065 ;
        RECT 49.975 193.735 50.800 194.065 ;
        RECT 50.970 193.735 51.315 194.065 ;
        RECT 51.505 193.815 51.835 194.065 ;
        RECT 49.635 193.565 49.805 193.735 ;
        RECT 48.295 192.825 48.465 193.435 ;
        RECT 48.635 193.045 48.965 193.480 ;
        RECT 49.190 193.155 49.465 193.500 ;
        RECT 49.635 193.395 51.300 193.565 ;
        RECT 49.655 192.825 50.035 193.225 ;
        RECT 50.205 193.045 50.375 193.395 ;
        RECT 50.545 192.825 50.875 193.225 ;
        RECT 51.045 193.045 51.300 193.395 ;
        RECT 51.525 192.825 51.755 193.645 ;
        RECT 52.005 193.625 52.255 194.225 ;
        RECT 54.295 194.065 54.465 194.625 ;
        RECT 54.725 194.525 55.900 194.695 ;
        RECT 56.070 194.575 56.350 195.375 ;
        RECT 54.725 194.235 55.055 194.525 ;
        RECT 55.730 194.405 55.900 194.525 ;
        RECT 55.225 194.065 55.470 194.355 ;
        RECT 55.730 194.235 56.390 194.405 ;
        RECT 56.560 194.235 56.835 195.205 ;
        RECT 56.220 194.065 56.390 194.235 ;
        RECT 53.790 193.815 54.125 194.065 ;
        RECT 54.295 193.735 55.010 194.065 ;
        RECT 55.225 193.735 56.050 194.065 ;
        RECT 56.220 193.735 56.495 194.065 ;
        RECT 54.295 193.645 54.545 193.735 ;
        RECT 51.925 192.995 52.255 193.625 ;
        RECT 52.425 192.825 52.635 193.645 ;
        RECT 53.785 192.825 54.045 193.645 ;
        RECT 54.215 193.225 54.545 193.645 ;
        RECT 56.220 193.565 56.390 193.735 ;
        RECT 54.725 193.395 56.390 193.565 ;
        RECT 56.665 193.500 56.835 194.235 ;
        RECT 57.005 194.210 57.295 195.375 ;
        RECT 57.485 194.785 57.725 195.175 ;
        RECT 57.895 194.965 58.245 195.375 ;
        RECT 57.485 194.585 58.235 194.785 ;
        RECT 54.725 192.995 54.985 193.395 ;
        RECT 55.155 192.825 55.485 193.225 ;
        RECT 55.655 193.045 55.825 193.395 ;
        RECT 55.995 192.825 56.370 193.225 ;
        RECT 56.560 193.155 56.835 193.500 ;
        RECT 57.005 192.825 57.295 193.550 ;
        RECT 57.485 193.065 57.715 194.405 ;
        RECT 57.895 193.905 58.235 194.585 ;
        RECT 58.415 194.085 58.745 195.195 ;
        RECT 58.915 194.725 59.095 195.195 ;
        RECT 59.265 194.895 59.595 195.375 ;
        RECT 59.770 194.725 59.940 195.195 ;
        RECT 58.915 194.525 59.940 194.725 ;
        RECT 57.895 193.005 58.125 193.905 ;
        RECT 58.415 193.785 58.960 194.085 ;
        RECT 58.325 192.825 58.570 193.605 ;
        RECT 58.740 193.555 58.960 193.785 ;
        RECT 59.130 193.735 59.555 194.355 ;
        RECT 59.750 193.735 60.010 194.355 ;
        RECT 60.205 194.235 60.490 195.375 ;
        RECT 60.220 193.555 60.480 194.065 ;
        RECT 58.740 193.365 60.480 193.555 ;
        RECT 58.740 193.005 59.170 193.365 ;
        RECT 59.750 192.825 60.480 193.195 ;
        RECT 60.680 193.005 60.960 195.195 ;
        RECT 61.145 194.285 64.655 195.375 ;
        RECT 61.145 193.595 62.795 194.115 ;
        RECT 62.965 193.765 64.655 194.285 ;
        RECT 61.145 192.825 64.655 193.595 ;
        RECT 65.300 193.005 65.580 195.195 ;
        RECT 65.770 194.235 66.055 195.375 ;
        RECT 66.320 194.725 66.490 195.195 ;
        RECT 66.665 194.895 66.995 195.375 ;
        RECT 67.165 194.725 67.345 195.195 ;
        RECT 66.320 194.525 67.345 194.725 ;
        RECT 65.780 193.555 66.040 194.065 ;
        RECT 66.250 193.735 66.510 194.355 ;
        RECT 66.705 193.735 67.130 194.355 ;
        RECT 67.515 194.085 67.845 195.195 ;
        RECT 68.015 194.965 68.365 195.375 ;
        RECT 68.535 194.785 68.775 195.175 ;
        RECT 67.300 193.785 67.845 194.085 ;
        RECT 68.025 194.585 68.775 194.785 ;
        RECT 68.025 193.905 68.365 194.585 ;
        RECT 67.300 193.555 67.520 193.785 ;
        RECT 65.780 193.365 67.520 193.555 ;
        RECT 65.780 192.825 66.510 193.195 ;
        RECT 67.090 193.005 67.520 193.365 ;
        RECT 67.690 192.825 67.935 193.605 ;
        RECT 68.135 193.005 68.365 193.905 ;
        RECT 68.545 193.065 68.775 194.405 ;
        RECT 68.965 194.235 69.240 195.205 ;
        RECT 69.450 194.575 69.730 195.375 ;
        RECT 69.900 194.865 71.515 195.195 ;
        RECT 69.900 194.525 71.075 194.695 ;
        RECT 69.900 194.405 70.070 194.525 ;
        RECT 69.410 194.235 70.070 194.405 ;
        RECT 68.965 193.500 69.135 194.235 ;
        RECT 69.410 194.065 69.580 194.235 ;
        RECT 70.330 194.065 70.575 194.355 ;
        RECT 70.745 194.235 71.075 194.525 ;
        RECT 71.335 194.065 71.505 194.625 ;
        RECT 71.755 194.235 72.015 195.375 ;
        RECT 72.385 194.705 72.665 195.375 ;
        RECT 72.835 194.485 73.135 195.035 ;
        RECT 73.335 194.655 73.665 195.375 ;
        RECT 73.855 194.655 74.315 195.205 ;
        RECT 72.200 194.065 72.465 194.425 ;
        RECT 72.835 194.315 73.775 194.485 ;
        RECT 73.605 194.065 73.775 194.315 ;
        RECT 69.305 193.735 69.580 194.065 ;
        RECT 69.750 193.735 70.575 194.065 ;
        RECT 70.790 193.735 71.505 194.065 ;
        RECT 71.675 193.815 72.010 194.065 ;
        RECT 72.200 193.815 72.875 194.065 ;
        RECT 73.095 193.815 73.435 194.065 ;
        RECT 69.410 193.565 69.580 193.735 ;
        RECT 71.255 193.645 71.505 193.735 ;
        RECT 73.605 193.735 73.895 194.065 ;
        RECT 73.605 193.645 73.775 193.735 ;
        RECT 68.965 193.155 69.240 193.500 ;
        RECT 69.410 193.395 71.075 193.565 ;
        RECT 69.430 192.825 69.805 193.225 ;
        RECT 69.975 193.045 70.145 193.395 ;
        RECT 70.315 192.825 70.645 193.225 ;
        RECT 70.815 192.995 71.075 193.395 ;
        RECT 71.255 193.225 71.585 193.645 ;
        RECT 71.755 192.825 72.015 193.645 ;
        RECT 72.385 193.455 73.775 193.645 ;
        RECT 72.385 193.095 72.715 193.455 ;
        RECT 74.065 193.285 74.315 194.655 ;
        RECT 74.485 194.235 74.745 195.375 ;
        RECT 74.915 194.225 75.245 195.205 ;
        RECT 75.415 194.235 75.695 195.375 ;
        RECT 75.955 194.405 76.125 195.205 ;
        RECT 76.885 194.745 77.135 195.205 ;
        RECT 77.335 194.995 78.005 195.375 ;
        RECT 78.195 194.745 78.445 195.205 ;
        RECT 78.620 194.915 78.865 195.375 ;
        RECT 76.885 194.575 78.445 194.745 ;
        RECT 79.035 194.525 79.375 195.165 ;
        RECT 75.955 194.235 78.895 194.405 ;
        RECT 74.505 193.815 74.840 194.065 ;
        RECT 75.010 193.625 75.180 194.225 ;
        RECT 78.725 194.065 78.895 194.235 ;
        RECT 75.350 193.795 75.685 194.065 ;
        RECT 75.925 193.735 76.110 194.065 ;
        RECT 76.365 193.735 76.840 194.065 ;
        RECT 77.150 193.735 77.495 194.065 ;
        RECT 73.335 192.825 73.585 193.285 ;
        RECT 73.755 192.995 74.315 193.285 ;
        RECT 74.485 192.995 75.180 193.625 ;
        RECT 75.385 192.825 75.695 193.625 ;
        RECT 75.955 193.395 77.135 193.565 ;
        RECT 77.305 193.505 77.495 193.735 ;
        RECT 77.755 193.490 77.950 194.065 ;
        RECT 78.220 193.735 78.555 194.065 ;
        RECT 78.725 193.735 79.035 194.065 ;
        RECT 78.725 193.565 78.895 193.735 ;
        RECT 75.955 192.995 76.125 193.395 ;
        RECT 76.365 192.825 76.695 193.225 ;
        RECT 76.965 193.165 77.135 193.395 ;
        RECT 78.200 193.395 78.895 193.565 ;
        RECT 79.205 193.410 79.375 194.525 ;
        RECT 79.730 194.405 80.120 194.580 ;
        RECT 80.605 194.575 80.935 195.375 ;
        RECT 81.105 194.585 81.640 195.205 ;
        RECT 79.730 194.235 81.155 194.405 ;
        RECT 79.605 193.505 79.960 194.065 ;
        RECT 78.200 193.165 78.370 193.395 ;
        RECT 76.965 192.995 78.370 193.165 ;
        RECT 78.540 192.825 78.870 193.205 ;
        RECT 79.065 192.995 79.375 193.410 ;
        RECT 80.130 193.335 80.300 194.235 ;
        RECT 80.470 193.505 80.735 194.065 ;
        RECT 80.985 193.735 81.155 194.235 ;
        RECT 81.325 193.565 81.640 194.585 ;
        RECT 82.765 194.210 83.055 195.375 ;
        RECT 83.225 194.235 83.565 195.205 ;
        RECT 83.735 194.235 83.905 195.375 ;
        RECT 84.175 194.575 84.425 195.375 ;
        RECT 85.070 194.405 85.400 195.205 ;
        RECT 85.700 194.575 86.030 195.375 ;
        RECT 86.200 194.405 86.530 195.205 ;
        RECT 84.095 194.235 86.530 194.405 ;
        RECT 86.905 194.285 90.415 195.375 ;
        RECT 79.710 192.825 79.950 193.335 ;
        RECT 80.130 193.005 80.410 193.335 ;
        RECT 80.640 192.825 80.855 193.335 ;
        RECT 81.025 192.995 81.640 193.565 ;
        RECT 83.225 193.625 83.400 194.235 ;
        RECT 84.095 193.985 84.265 194.235 ;
        RECT 83.570 193.815 84.265 193.985 ;
        RECT 84.440 193.815 84.860 194.015 ;
        RECT 85.030 193.815 85.360 194.015 ;
        RECT 85.530 193.815 85.860 194.015 ;
        RECT 82.765 192.825 83.055 193.550 ;
        RECT 83.225 192.995 83.565 193.625 ;
        RECT 83.735 192.825 83.985 193.625 ;
        RECT 84.175 193.475 85.400 193.645 ;
        RECT 84.175 192.995 84.505 193.475 ;
        RECT 84.675 192.825 84.900 193.285 ;
        RECT 85.070 192.995 85.400 193.475 ;
        RECT 86.030 193.605 86.200 194.235 ;
        RECT 86.385 193.815 86.735 194.065 ;
        RECT 86.030 192.995 86.530 193.605 ;
        RECT 86.905 193.595 88.555 194.115 ;
        RECT 88.725 193.765 90.415 194.285 ;
        RECT 91.045 194.285 92.255 195.375 ;
        RECT 91.045 193.745 91.565 194.285 ;
        RECT 86.905 192.825 90.415 193.595 ;
        RECT 91.735 193.575 92.255 194.115 ;
        RECT 91.045 192.825 92.255 193.575 ;
        RECT 18.280 192.655 92.340 192.825 ;
        RECT 18.365 191.905 19.575 192.655 ;
        RECT 19.745 192.110 25.090 192.655 ;
        RECT 25.265 192.110 30.610 192.655 ;
        RECT 30.785 192.110 36.130 192.655 ;
        RECT 18.365 191.365 18.885 191.905 ;
        RECT 19.055 191.195 19.575 191.735 ;
        RECT 21.330 191.280 21.670 192.110 ;
        RECT 18.365 190.105 19.575 191.195 ;
        RECT 23.150 190.540 23.500 191.790 ;
        RECT 26.850 191.280 27.190 192.110 ;
        RECT 28.670 190.540 29.020 191.790 ;
        RECT 32.370 191.280 32.710 192.110 ;
        RECT 36.765 191.980 37.040 192.325 ;
        RECT 37.230 192.255 37.605 192.655 ;
        RECT 37.775 192.085 37.945 192.435 ;
        RECT 38.115 192.255 38.445 192.655 ;
        RECT 38.615 192.085 38.875 192.485 ;
        RECT 34.190 190.540 34.540 191.790 ;
        RECT 36.765 191.245 36.935 191.980 ;
        RECT 37.210 191.915 38.875 192.085 ;
        RECT 37.210 191.745 37.380 191.915 ;
        RECT 39.055 191.835 39.385 192.255 ;
        RECT 39.555 191.835 39.815 192.655 ;
        RECT 39.985 191.885 43.495 192.655 ;
        RECT 44.125 191.930 44.415 192.655 ;
        RECT 44.585 192.110 49.930 192.655 ;
        RECT 39.055 191.745 39.305 191.835 ;
        RECT 37.105 191.415 37.380 191.745 ;
        RECT 37.550 191.415 38.375 191.745 ;
        RECT 38.590 191.415 39.305 191.745 ;
        RECT 39.475 191.415 39.810 191.665 ;
        RECT 37.210 191.245 37.380 191.415 ;
        RECT 19.745 190.105 25.090 190.540 ;
        RECT 25.265 190.105 30.610 190.540 ;
        RECT 30.785 190.105 36.130 190.540 ;
        RECT 36.765 190.275 37.040 191.245 ;
        RECT 37.210 191.075 37.870 191.245 ;
        RECT 38.130 191.125 38.375 191.415 ;
        RECT 37.700 190.955 37.870 191.075 ;
        RECT 38.545 190.955 38.875 191.245 ;
        RECT 37.250 190.105 37.530 190.905 ;
        RECT 37.700 190.785 38.875 190.955 ;
        RECT 39.135 190.855 39.305 191.415 ;
        RECT 39.985 191.365 41.635 191.885 ;
        RECT 37.700 190.285 39.315 190.615 ;
        RECT 39.555 190.105 39.815 191.245 ;
        RECT 41.805 191.195 43.495 191.715 ;
        RECT 46.170 191.280 46.510 192.110 ;
        RECT 50.105 191.885 53.615 192.655 ;
        RECT 54.705 192.045 55.045 192.460 ;
        RECT 55.215 192.215 55.385 192.655 ;
        RECT 55.555 192.265 56.805 192.445 ;
        RECT 55.555 192.045 55.885 192.265 ;
        RECT 57.075 192.195 57.245 192.655 ;
        RECT 39.985 190.105 43.495 191.195 ;
        RECT 44.125 190.105 44.415 191.270 ;
        RECT 47.990 190.540 48.340 191.790 ;
        RECT 50.105 191.365 51.755 191.885 ;
        RECT 54.705 191.875 55.885 192.045 ;
        RECT 56.055 192.025 56.420 192.095 ;
        RECT 56.055 191.845 57.305 192.025 ;
        RECT 51.925 191.195 53.615 191.715 ;
        RECT 54.705 191.465 55.170 191.665 ;
        RECT 55.345 191.415 55.675 191.665 ;
        RECT 55.845 191.635 56.310 191.665 ;
        RECT 55.845 191.465 56.315 191.635 ;
        RECT 55.845 191.415 56.310 191.465 ;
        RECT 56.505 191.415 56.860 191.665 ;
        RECT 55.345 191.295 55.525 191.415 ;
        RECT 44.585 190.105 49.930 190.540 ;
        RECT 50.105 190.105 53.615 191.195 ;
        RECT 54.705 190.105 55.025 191.285 ;
        RECT 55.195 191.125 55.525 191.295 ;
        RECT 57.030 191.245 57.305 191.845 ;
        RECT 55.195 190.335 55.395 191.125 ;
        RECT 55.695 191.035 57.305 191.245 ;
        RECT 55.695 190.935 56.105 191.035 ;
        RECT 55.720 190.275 56.105 190.935 ;
        RECT 56.500 190.105 57.285 190.865 ;
        RECT 57.475 190.275 57.755 192.375 ;
        RECT 57.930 192.150 58.265 192.655 ;
        RECT 58.435 192.085 58.675 192.460 ;
        RECT 58.955 192.325 59.125 192.470 ;
        RECT 58.955 192.130 59.330 192.325 ;
        RECT 59.690 192.160 60.085 192.655 ;
        RECT 57.985 191.125 58.285 191.975 ;
        RECT 58.455 191.935 58.675 192.085 ;
        RECT 58.455 191.605 58.990 191.935 ;
        RECT 59.160 191.795 59.330 192.130 ;
        RECT 60.255 191.965 60.495 192.485 ;
        RECT 58.455 190.955 58.690 191.605 ;
        RECT 59.160 191.435 60.145 191.795 ;
        RECT 58.015 190.725 58.690 190.955 ;
        RECT 58.860 191.415 60.145 191.435 ;
        RECT 58.860 191.265 59.720 191.415 ;
        RECT 58.015 190.295 58.185 190.725 ;
        RECT 58.355 190.105 58.685 190.555 ;
        RECT 58.860 190.320 59.145 191.265 ;
        RECT 60.320 191.160 60.495 191.965 ;
        RECT 60.685 191.885 62.355 192.655 ;
        RECT 62.990 192.150 63.325 192.655 ;
        RECT 63.495 192.085 63.735 192.460 ;
        RECT 64.015 192.325 64.185 192.470 ;
        RECT 64.015 192.130 64.390 192.325 ;
        RECT 64.750 192.160 65.145 192.655 ;
        RECT 60.685 191.365 61.435 191.885 ;
        RECT 61.605 191.195 62.355 191.715 ;
        RECT 59.320 190.785 60.015 191.095 ;
        RECT 59.325 190.105 60.010 190.575 ;
        RECT 60.190 190.375 60.495 191.160 ;
        RECT 60.685 190.105 62.355 191.195 ;
        RECT 63.045 191.125 63.345 191.975 ;
        RECT 63.515 191.935 63.735 192.085 ;
        RECT 63.515 191.605 64.050 191.935 ;
        RECT 64.220 191.795 64.390 192.130 ;
        RECT 65.315 191.965 65.555 192.485 ;
        RECT 63.515 190.955 63.750 191.605 ;
        RECT 64.220 191.435 65.205 191.795 ;
        RECT 63.075 190.725 63.750 190.955 ;
        RECT 63.920 191.415 65.205 191.435 ;
        RECT 63.920 191.265 64.780 191.415 ;
        RECT 63.075 190.295 63.245 190.725 ;
        RECT 63.415 190.105 63.745 190.555 ;
        RECT 63.920 190.320 64.205 191.265 ;
        RECT 65.380 191.160 65.555 191.965 ;
        RECT 65.745 191.885 69.255 192.655 ;
        RECT 69.885 191.930 70.175 192.655 ;
        RECT 70.345 192.110 75.690 192.655 ;
        RECT 65.745 191.365 67.395 191.885 ;
        RECT 67.565 191.195 69.255 191.715 ;
        RECT 71.930 191.280 72.270 192.110 ;
        RECT 76.985 192.025 77.315 192.385 ;
        RECT 77.935 192.195 78.185 192.655 ;
        RECT 78.355 192.195 78.915 192.485 ;
        RECT 76.985 191.835 78.375 192.025 ;
        RECT 64.380 190.785 65.075 191.095 ;
        RECT 64.385 190.105 65.070 190.575 ;
        RECT 65.250 190.375 65.555 191.160 ;
        RECT 65.745 190.105 69.255 191.195 ;
        RECT 69.885 190.105 70.175 191.270 ;
        RECT 73.750 190.540 74.100 191.790 ;
        RECT 78.205 191.745 78.375 191.835 ;
        RECT 76.800 191.415 77.475 191.665 ;
        RECT 77.695 191.415 78.035 191.665 ;
        RECT 78.205 191.415 78.495 191.745 ;
        RECT 76.800 191.055 77.065 191.415 ;
        RECT 78.205 191.165 78.375 191.415 ;
        RECT 77.435 190.995 78.375 191.165 ;
        RECT 70.345 190.105 75.690 190.540 ;
        RECT 76.985 190.105 77.265 190.775 ;
        RECT 77.435 190.445 77.735 190.995 ;
        RECT 78.665 190.825 78.915 192.195 ;
        RECT 79.085 191.885 81.675 192.655 ;
        RECT 82.395 192.105 82.565 192.395 ;
        RECT 82.735 192.275 83.065 192.655 ;
        RECT 82.395 191.935 83.060 192.105 ;
        RECT 79.085 191.365 80.295 191.885 ;
        RECT 80.465 191.195 81.675 191.715 ;
        RECT 77.935 190.105 78.265 190.825 ;
        RECT 78.455 190.275 78.915 190.825 ;
        RECT 79.085 190.105 81.675 191.195 ;
        RECT 82.310 191.115 82.660 191.765 ;
        RECT 82.830 190.945 83.060 191.935 ;
        RECT 82.395 190.775 83.060 190.945 ;
        RECT 82.395 190.275 82.565 190.775 ;
        RECT 82.735 190.105 83.065 190.605 ;
        RECT 83.235 190.275 83.460 192.395 ;
        RECT 83.675 192.195 83.925 192.655 ;
        RECT 84.110 192.205 84.440 192.375 ;
        RECT 84.620 192.205 85.370 192.375 ;
        RECT 83.660 191.075 83.940 191.675 ;
        RECT 84.110 190.675 84.280 192.205 ;
        RECT 84.450 191.705 85.030 192.035 ;
        RECT 84.450 190.835 84.690 191.705 ;
        RECT 85.200 191.425 85.370 192.205 ;
        RECT 85.620 192.155 85.990 192.655 ;
        RECT 86.170 192.205 86.630 192.375 ;
        RECT 86.860 192.205 87.530 192.375 ;
        RECT 86.170 191.975 86.340 192.205 ;
        RECT 85.540 191.675 86.340 191.975 ;
        RECT 86.510 191.705 87.060 192.035 ;
        RECT 85.540 191.645 85.710 191.675 ;
        RECT 85.830 191.425 86.000 191.495 ;
        RECT 85.200 191.255 86.000 191.425 ;
        RECT 85.490 191.165 86.000 191.255 ;
        RECT 84.880 190.730 85.320 191.085 ;
        RECT 83.660 190.105 83.925 190.565 ;
        RECT 84.110 190.300 84.345 190.675 ;
        RECT 85.490 190.550 85.660 191.165 ;
        RECT 84.590 190.380 85.660 190.550 ;
        RECT 85.830 190.105 86.000 190.905 ;
        RECT 86.170 190.605 86.340 191.675 ;
        RECT 86.510 190.775 86.700 191.495 ;
        RECT 86.870 191.165 87.060 191.705 ;
        RECT 87.360 191.665 87.530 192.205 ;
        RECT 87.845 192.125 88.015 192.655 ;
        RECT 88.310 192.005 88.670 192.445 ;
        RECT 88.845 192.175 89.015 192.655 ;
        RECT 89.205 192.010 89.540 192.435 ;
        RECT 89.715 192.180 89.885 192.655 ;
        RECT 90.060 192.010 90.395 192.435 ;
        RECT 90.565 192.180 90.735 192.655 ;
        RECT 88.310 191.835 88.810 192.005 ;
        RECT 89.205 191.840 90.875 192.010 ;
        RECT 91.045 191.905 92.255 192.655 ;
        RECT 88.640 191.665 88.810 191.835 ;
        RECT 87.360 191.495 88.450 191.665 ;
        RECT 88.640 191.495 90.460 191.665 ;
        RECT 86.870 190.835 87.190 191.165 ;
        RECT 86.170 190.275 86.420 190.605 ;
        RECT 87.360 190.575 87.530 191.495 ;
        RECT 88.640 191.240 88.810 191.495 ;
        RECT 90.630 191.275 90.875 191.840 ;
        RECT 87.700 191.070 88.810 191.240 ;
        RECT 89.205 191.105 90.875 191.275 ;
        RECT 91.045 191.195 91.565 191.735 ;
        RECT 91.735 191.365 92.255 191.905 ;
        RECT 87.700 190.910 88.560 191.070 ;
        RECT 86.645 190.405 87.530 190.575 ;
        RECT 87.710 190.105 87.925 190.605 ;
        RECT 88.390 190.285 88.560 190.910 ;
        RECT 88.845 190.105 89.025 190.885 ;
        RECT 89.205 190.345 89.540 191.105 ;
        RECT 89.720 190.105 89.890 190.935 ;
        RECT 90.060 190.345 90.390 191.105 ;
        RECT 90.560 190.105 90.730 190.935 ;
        RECT 91.045 190.105 92.255 191.195 ;
        RECT 18.280 189.935 92.340 190.105 ;
        RECT 18.365 188.845 19.575 189.935 ;
        RECT 19.745 189.500 25.090 189.935 ;
        RECT 25.265 189.500 30.610 189.935 ;
        RECT 18.365 188.135 18.885 188.675 ;
        RECT 19.055 188.305 19.575 188.845 ;
        RECT 18.365 187.385 19.575 188.135 ;
        RECT 21.330 187.930 21.670 188.760 ;
        RECT 23.150 188.250 23.500 189.500 ;
        RECT 26.850 187.930 27.190 188.760 ;
        RECT 28.670 188.250 29.020 189.500 ;
        RECT 31.245 188.770 31.535 189.935 ;
        RECT 31.705 188.845 34.295 189.935 ;
        RECT 31.705 188.155 32.915 188.675 ;
        RECT 33.085 188.325 34.295 188.845 ;
        RECT 34.465 189.085 34.845 189.765 ;
        RECT 35.435 189.085 35.605 189.935 ;
        RECT 35.775 189.255 36.105 189.765 ;
        RECT 36.275 189.425 36.445 189.935 ;
        RECT 36.615 189.255 37.015 189.765 ;
        RECT 35.775 189.085 37.015 189.255 ;
        RECT 19.745 187.385 25.090 187.930 ;
        RECT 25.265 187.385 30.610 187.930 ;
        RECT 31.245 187.385 31.535 188.110 ;
        RECT 31.705 187.385 34.295 188.155 ;
        RECT 34.465 188.125 34.635 189.085 ;
        RECT 34.805 188.745 36.110 188.915 ;
        RECT 37.195 188.835 37.515 189.765 ;
        RECT 37.685 188.845 40.275 189.935 ;
        RECT 34.805 188.295 35.050 188.745 ;
        RECT 35.220 188.375 35.770 188.575 ;
        RECT 35.940 188.545 36.110 188.745 ;
        RECT 36.885 188.665 37.515 188.835 ;
        RECT 35.940 188.375 36.315 188.545 ;
        RECT 36.485 188.125 36.715 188.625 ;
        RECT 34.465 187.955 36.715 188.125 ;
        RECT 34.515 187.385 34.845 187.775 ;
        RECT 35.015 187.635 35.185 187.955 ;
        RECT 36.885 187.785 37.055 188.665 ;
        RECT 35.355 187.385 35.685 187.775 ;
        RECT 36.100 187.615 37.055 187.785 ;
        RECT 37.225 187.385 37.515 188.220 ;
        RECT 37.685 188.155 38.895 188.675 ;
        RECT 39.065 188.325 40.275 188.845 ;
        RECT 41.110 188.965 41.440 189.765 ;
        RECT 41.610 189.135 41.940 189.935 ;
        RECT 42.240 188.965 42.570 189.765 ;
        RECT 43.215 189.135 43.465 189.935 ;
        RECT 41.110 188.795 43.545 188.965 ;
        RECT 43.735 188.795 43.905 189.935 ;
        RECT 44.075 188.795 44.415 189.765 ;
        RECT 44.585 188.845 46.255 189.935 ;
        RECT 46.975 189.315 47.145 189.745 ;
        RECT 47.315 189.485 47.645 189.935 ;
        RECT 46.975 189.085 47.650 189.315 ;
        RECT 40.905 188.375 41.255 188.625 ;
        RECT 41.440 188.165 41.610 188.795 ;
        RECT 41.780 188.375 42.110 188.575 ;
        RECT 42.280 188.375 42.610 188.575 ;
        RECT 42.780 188.375 43.200 188.575 ;
        RECT 43.375 188.545 43.545 188.795 ;
        RECT 43.375 188.375 44.070 188.545 ;
        RECT 37.685 187.385 40.275 188.155 ;
        RECT 41.110 187.555 41.610 188.165 ;
        RECT 42.240 188.035 43.465 188.205 ;
        RECT 44.240 188.185 44.415 188.795 ;
        RECT 42.240 187.555 42.570 188.035 ;
        RECT 42.740 187.385 42.965 187.845 ;
        RECT 43.135 187.555 43.465 188.035 ;
        RECT 43.655 187.385 43.905 188.185 ;
        RECT 44.075 187.555 44.415 188.185 ;
        RECT 44.585 188.155 45.335 188.675 ;
        RECT 45.505 188.325 46.255 188.845 ;
        RECT 44.585 187.385 46.255 188.155 ;
        RECT 46.945 188.065 47.245 188.915 ;
        RECT 47.415 188.435 47.650 189.085 ;
        RECT 47.820 188.775 48.105 189.720 ;
        RECT 48.285 189.465 48.970 189.935 ;
        RECT 48.280 188.945 48.975 189.255 ;
        RECT 49.150 188.880 49.455 189.665 ;
        RECT 47.820 188.625 48.680 188.775 ;
        RECT 47.820 188.605 49.105 188.625 ;
        RECT 47.415 188.105 47.950 188.435 ;
        RECT 48.120 188.245 49.105 188.605 ;
        RECT 47.415 187.955 47.635 188.105 ;
        RECT 46.890 187.385 47.225 187.890 ;
        RECT 47.395 187.580 47.635 187.955 ;
        RECT 48.120 187.910 48.290 188.245 ;
        RECT 49.280 188.075 49.455 188.880 ;
        RECT 49.735 188.925 49.905 189.765 ;
        RECT 50.075 189.595 51.245 189.765 ;
        RECT 50.075 189.095 50.405 189.595 ;
        RECT 50.915 189.555 51.245 189.595 ;
        RECT 51.435 189.515 51.790 189.935 ;
        RECT 50.575 189.335 50.805 189.425 ;
        RECT 51.960 189.335 52.210 189.765 ;
        RECT 50.575 189.095 52.210 189.335 ;
        RECT 52.380 189.175 52.710 189.935 ;
        RECT 52.880 189.095 53.135 189.765 ;
        RECT 49.735 188.755 52.795 188.925 ;
        RECT 49.650 188.375 50.000 188.585 ;
        RECT 50.170 188.375 50.615 188.575 ;
        RECT 50.785 188.375 51.260 188.575 ;
        RECT 47.915 187.715 48.290 187.910 ;
        RECT 47.915 187.570 48.085 187.715 ;
        RECT 48.650 187.385 49.045 187.880 ;
        RECT 49.215 187.555 49.455 188.075 ;
        RECT 49.735 188.035 50.800 188.205 ;
        RECT 49.735 187.555 49.905 188.035 ;
        RECT 50.075 187.385 50.405 187.865 ;
        RECT 50.630 187.805 50.800 188.035 ;
        RECT 50.980 187.975 51.260 188.375 ;
        RECT 51.530 188.375 51.860 188.575 ;
        RECT 52.030 188.405 52.405 188.575 ;
        RECT 52.030 188.375 52.395 188.405 ;
        RECT 51.530 187.975 51.815 188.375 ;
        RECT 52.625 188.205 52.795 188.755 ;
        RECT 51.995 188.035 52.795 188.205 ;
        RECT 51.995 187.805 52.165 188.035 ;
        RECT 52.965 187.965 53.135 189.095 ;
        RECT 52.950 187.895 53.135 187.965 ;
        RECT 52.925 187.885 53.135 187.895 ;
        RECT 50.630 187.555 52.165 187.805 ;
        RECT 52.335 187.385 52.665 187.865 ;
        RECT 52.880 187.555 53.135 187.885 ;
        RECT 53.325 188.825 53.585 189.765 ;
        RECT 53.755 189.535 54.085 189.935 ;
        RECT 55.230 189.670 55.485 189.765 ;
        RECT 54.345 189.500 55.485 189.670 ;
        RECT 55.655 189.555 55.985 189.725 ;
        RECT 54.345 189.275 54.515 189.500 ;
        RECT 53.755 189.105 54.515 189.275 ;
        RECT 55.230 189.365 55.485 189.500 ;
        RECT 53.325 188.110 53.500 188.825 ;
        RECT 53.755 188.625 53.925 189.105 ;
        RECT 54.780 189.015 54.950 189.205 ;
        RECT 55.230 189.195 55.640 189.365 ;
        RECT 53.670 188.295 53.925 188.625 ;
        RECT 54.150 188.295 54.480 188.915 ;
        RECT 54.780 188.845 55.300 189.015 ;
        RECT 54.650 188.295 54.940 188.675 ;
        RECT 55.130 188.125 55.300 188.845 ;
        RECT 53.325 187.555 53.585 188.110 ;
        RECT 54.420 187.955 55.300 188.125 ;
        RECT 55.470 188.170 55.640 189.195 ;
        RECT 55.815 189.305 55.985 189.555 ;
        RECT 56.155 189.475 56.405 189.935 ;
        RECT 56.575 189.305 56.755 189.765 ;
        RECT 55.815 189.135 56.755 189.305 ;
        RECT 55.840 188.655 56.320 188.955 ;
        RECT 55.470 188.000 55.820 188.170 ;
        RECT 56.060 188.065 56.320 188.655 ;
        RECT 56.520 188.065 56.780 188.955 ;
        RECT 57.005 188.770 57.295 189.935 ;
        RECT 58.405 189.095 58.660 189.765 ;
        RECT 58.830 189.175 59.160 189.935 ;
        RECT 59.330 189.335 59.580 189.765 ;
        RECT 59.750 189.515 60.105 189.935 ;
        RECT 60.295 189.595 61.465 189.765 ;
        RECT 60.295 189.555 60.625 189.595 ;
        RECT 60.735 189.335 60.965 189.425 ;
        RECT 59.330 189.095 60.965 189.335 ;
        RECT 61.135 189.095 61.465 189.595 ;
        RECT 53.755 187.385 54.185 187.830 ;
        RECT 54.420 187.555 54.590 187.955 ;
        RECT 54.760 187.385 55.480 187.785 ;
        RECT 55.650 187.555 55.820 188.000 ;
        RECT 56.395 187.385 56.795 187.895 ;
        RECT 57.005 187.385 57.295 188.110 ;
        RECT 58.405 187.965 58.575 189.095 ;
        RECT 61.635 188.925 61.805 189.765 ;
        RECT 58.745 188.755 61.805 188.925 ;
        RECT 62.065 188.845 63.735 189.935 ;
        RECT 63.995 189.265 64.165 189.765 ;
        RECT 64.335 189.435 64.665 189.935 ;
        RECT 63.995 189.095 64.660 189.265 ;
        RECT 58.745 188.205 58.915 188.755 ;
        RECT 59.135 188.405 59.510 188.575 ;
        RECT 59.145 188.375 59.510 188.405 ;
        RECT 59.680 188.375 60.010 188.575 ;
        RECT 58.745 188.035 59.545 188.205 ;
        RECT 58.405 187.895 58.590 187.965 ;
        RECT 58.405 187.885 58.615 187.895 ;
        RECT 58.405 187.555 58.660 187.885 ;
        RECT 58.875 187.385 59.205 187.865 ;
        RECT 59.375 187.805 59.545 188.035 ;
        RECT 59.725 187.975 60.010 188.375 ;
        RECT 60.280 188.375 60.755 188.575 ;
        RECT 60.925 188.375 61.370 188.575 ;
        RECT 61.540 188.375 61.890 188.585 ;
        RECT 60.280 187.975 60.560 188.375 ;
        RECT 60.740 188.035 61.805 188.205 ;
        RECT 60.740 187.805 60.910 188.035 ;
        RECT 59.375 187.555 60.910 187.805 ;
        RECT 61.135 187.385 61.465 187.865 ;
        RECT 61.635 187.555 61.805 188.035 ;
        RECT 62.065 188.155 62.815 188.675 ;
        RECT 62.985 188.325 63.735 188.845 ;
        RECT 63.910 188.275 64.260 188.925 ;
        RECT 62.065 187.385 63.735 188.155 ;
        RECT 64.430 188.105 64.660 189.095 ;
        RECT 63.995 187.935 64.660 188.105 ;
        RECT 63.995 187.645 64.165 187.935 ;
        RECT 64.335 187.385 64.665 187.765 ;
        RECT 64.835 187.645 65.020 189.765 ;
        RECT 65.260 189.475 65.525 189.935 ;
        RECT 65.695 189.340 65.945 189.765 ;
        RECT 66.155 189.490 67.260 189.660 ;
        RECT 65.640 189.210 65.945 189.340 ;
        RECT 65.190 188.015 65.470 188.965 ;
        RECT 65.640 188.105 65.810 189.210 ;
        RECT 65.980 188.425 66.220 189.020 ;
        RECT 66.390 188.955 66.920 189.320 ;
        RECT 66.390 188.255 66.560 188.955 ;
        RECT 67.090 188.875 67.260 189.490 ;
        RECT 67.430 189.135 67.600 189.935 ;
        RECT 67.770 189.435 68.020 189.765 ;
        RECT 68.245 189.465 69.130 189.635 ;
        RECT 67.090 188.785 67.600 188.875 ;
        RECT 65.640 187.975 65.865 188.105 ;
        RECT 66.035 188.035 66.560 188.255 ;
        RECT 66.730 188.615 67.600 188.785 ;
        RECT 65.275 187.385 65.525 187.845 ;
        RECT 65.695 187.835 65.865 187.975 ;
        RECT 66.730 187.835 66.900 188.615 ;
        RECT 67.430 188.545 67.600 188.615 ;
        RECT 67.110 188.365 67.310 188.395 ;
        RECT 67.770 188.365 67.940 189.435 ;
        RECT 68.110 188.545 68.300 189.265 ;
        RECT 67.110 188.065 67.940 188.365 ;
        RECT 68.470 188.335 68.790 189.295 ;
        RECT 65.695 187.665 66.030 187.835 ;
        RECT 66.225 187.665 66.900 187.835 ;
        RECT 67.220 187.385 67.590 187.885 ;
        RECT 67.770 187.835 67.940 188.065 ;
        RECT 68.325 188.005 68.790 188.335 ;
        RECT 68.960 188.625 69.130 189.465 ;
        RECT 69.310 189.435 69.625 189.935 ;
        RECT 69.855 189.205 70.195 189.765 ;
        RECT 69.300 188.830 70.195 189.205 ;
        RECT 70.365 188.925 70.535 189.935 ;
        RECT 70.005 188.625 70.195 188.830 ;
        RECT 70.705 188.875 71.035 189.720 ;
        RECT 70.705 188.795 71.095 188.875 ;
        RECT 70.880 188.745 71.095 188.795 ;
        RECT 68.960 188.295 69.835 188.625 ;
        RECT 70.005 188.295 70.755 188.625 ;
        RECT 68.960 187.835 69.130 188.295 ;
        RECT 70.005 188.125 70.205 188.295 ;
        RECT 70.925 188.165 71.095 188.745 ;
        RECT 70.870 188.125 71.095 188.165 ;
        RECT 67.770 187.665 68.175 187.835 ;
        RECT 68.345 187.665 69.130 187.835 ;
        RECT 69.405 187.385 69.615 187.915 ;
        RECT 69.875 187.600 70.205 188.125 ;
        RECT 70.715 188.040 71.095 188.125 ;
        RECT 71.265 188.795 71.650 189.765 ;
        RECT 71.820 189.475 72.145 189.935 ;
        RECT 72.665 189.305 72.945 189.765 ;
        RECT 71.820 189.085 72.945 189.305 ;
        RECT 71.265 188.125 71.545 188.795 ;
        RECT 71.820 188.625 72.270 189.085 ;
        RECT 73.135 188.915 73.535 189.765 ;
        RECT 73.935 189.475 74.205 189.935 ;
        RECT 74.375 189.305 74.660 189.765 ;
        RECT 71.715 188.295 72.270 188.625 ;
        RECT 72.440 188.355 73.535 188.915 ;
        RECT 71.820 188.185 72.270 188.295 ;
        RECT 70.375 187.385 70.545 187.995 ;
        RECT 70.715 187.605 71.045 188.040 ;
        RECT 71.265 187.555 71.650 188.125 ;
        RECT 71.820 188.015 72.945 188.185 ;
        RECT 71.820 187.385 72.145 187.845 ;
        RECT 72.665 187.555 72.945 188.015 ;
        RECT 73.135 187.555 73.535 188.355 ;
        RECT 73.705 189.085 74.660 189.305 ;
        RECT 73.705 188.185 73.915 189.085 ;
        RECT 74.085 188.355 74.775 188.915 ;
        RECT 75.875 188.795 76.205 189.935 ;
        RECT 76.735 188.965 77.065 189.750 ;
        RECT 76.385 188.795 77.065 188.965 ;
        RECT 77.245 188.845 78.915 189.935 ;
        RECT 75.865 188.375 76.215 188.625 ;
        RECT 76.385 188.195 76.555 188.795 ;
        RECT 76.725 188.375 77.075 188.625 ;
        RECT 73.705 188.015 74.660 188.185 ;
        RECT 73.935 187.385 74.205 187.845 ;
        RECT 74.375 187.555 74.660 188.015 ;
        RECT 75.875 187.385 76.145 188.195 ;
        RECT 76.315 187.555 76.645 188.195 ;
        RECT 76.815 187.385 77.055 188.195 ;
        RECT 77.245 188.155 77.995 188.675 ;
        RECT 78.165 188.325 78.915 188.845 ;
        RECT 79.085 189.065 79.360 189.765 ;
        RECT 79.530 189.390 79.785 189.935 ;
        RECT 79.955 189.425 80.435 189.765 ;
        RECT 80.610 189.380 81.215 189.935 ;
        RECT 80.600 189.280 81.215 189.380 ;
        RECT 80.600 189.255 80.785 189.280 ;
        RECT 77.245 187.385 78.915 188.155 ;
        RECT 79.085 188.035 79.255 189.065 ;
        RECT 79.530 188.935 80.285 189.185 ;
        RECT 80.455 189.010 80.785 189.255 ;
        RECT 79.530 188.900 80.300 188.935 ;
        RECT 79.530 188.890 80.315 188.900 ;
        RECT 79.425 188.875 80.320 188.890 ;
        RECT 79.425 188.860 80.340 188.875 ;
        RECT 79.425 188.850 80.360 188.860 ;
        RECT 79.425 188.840 80.385 188.850 ;
        RECT 79.425 188.810 80.455 188.840 ;
        RECT 79.425 188.780 80.475 188.810 ;
        RECT 79.425 188.750 80.495 188.780 ;
        RECT 79.425 188.725 80.525 188.750 ;
        RECT 79.425 188.690 80.560 188.725 ;
        RECT 79.425 188.685 80.590 188.690 ;
        RECT 79.425 188.290 79.655 188.685 ;
        RECT 80.200 188.680 80.590 188.685 ;
        RECT 80.225 188.670 80.590 188.680 ;
        RECT 80.240 188.665 80.590 188.670 ;
        RECT 80.255 188.660 80.590 188.665 ;
        RECT 80.955 188.660 81.215 189.110 ;
        RECT 81.385 188.845 82.595 189.935 ;
        RECT 80.255 188.655 81.215 188.660 ;
        RECT 80.265 188.645 81.215 188.655 ;
        RECT 80.275 188.640 81.215 188.645 ;
        RECT 80.285 188.630 81.215 188.640 ;
        RECT 80.290 188.620 81.215 188.630 ;
        RECT 80.295 188.615 81.215 188.620 ;
        RECT 80.305 188.600 81.215 188.615 ;
        RECT 80.310 188.585 81.215 188.600 ;
        RECT 80.320 188.560 81.215 188.585 ;
        RECT 79.825 188.090 80.155 188.515 ;
        RECT 79.085 187.555 79.345 188.035 ;
        RECT 79.515 187.385 79.765 187.925 ;
        RECT 79.935 187.605 80.155 188.090 ;
        RECT 80.325 188.490 81.215 188.560 ;
        RECT 80.325 187.765 80.495 188.490 ;
        RECT 80.665 187.935 81.215 188.320 ;
        RECT 81.385 188.135 81.905 188.675 ;
        RECT 82.075 188.305 82.595 188.845 ;
        RECT 82.765 188.770 83.055 189.935 ;
        RECT 83.225 188.795 83.565 189.765 ;
        RECT 83.735 188.795 83.905 189.935 ;
        RECT 84.175 189.135 84.425 189.935 ;
        RECT 85.070 188.965 85.400 189.765 ;
        RECT 85.700 189.135 86.030 189.935 ;
        RECT 86.200 188.965 86.530 189.765 ;
        RECT 84.095 188.795 86.530 188.965 ;
        RECT 86.905 188.845 90.415 189.935 ;
        RECT 83.225 188.185 83.400 188.795 ;
        RECT 84.095 188.545 84.265 188.795 ;
        RECT 83.570 188.375 84.265 188.545 ;
        RECT 84.440 188.375 84.860 188.575 ;
        RECT 85.030 188.375 85.360 188.575 ;
        RECT 85.530 188.375 85.860 188.575 ;
        RECT 80.325 187.595 81.215 187.765 ;
        RECT 81.385 187.385 82.595 188.135 ;
        RECT 82.765 187.385 83.055 188.110 ;
        RECT 83.225 187.555 83.565 188.185 ;
        RECT 83.735 187.385 83.985 188.185 ;
        RECT 84.175 188.035 85.400 188.205 ;
        RECT 84.175 187.555 84.505 188.035 ;
        RECT 84.675 187.385 84.900 187.845 ;
        RECT 85.070 187.555 85.400 188.035 ;
        RECT 86.030 188.165 86.200 188.795 ;
        RECT 86.385 188.375 86.735 188.625 ;
        RECT 86.030 187.555 86.530 188.165 ;
        RECT 86.905 188.155 88.555 188.675 ;
        RECT 88.725 188.325 90.415 188.845 ;
        RECT 91.045 188.845 92.255 189.935 ;
        RECT 91.045 188.305 91.565 188.845 ;
        RECT 86.905 187.385 90.415 188.155 ;
        RECT 91.735 188.135 92.255 188.675 ;
        RECT 91.045 187.385 92.255 188.135 ;
        RECT 18.280 187.215 92.340 187.385 ;
        RECT 18.365 186.465 19.575 187.215 ;
        RECT 19.745 186.670 25.090 187.215 ;
        RECT 25.265 186.670 30.610 187.215 ;
        RECT 18.365 185.925 18.885 186.465 ;
        RECT 19.055 185.755 19.575 186.295 ;
        RECT 21.330 185.840 21.670 186.670 ;
        RECT 18.365 184.665 19.575 185.755 ;
        RECT 23.150 185.100 23.500 186.350 ;
        RECT 26.850 185.840 27.190 186.670 ;
        RECT 30.785 186.445 34.295 187.215 ;
        RECT 34.490 186.565 34.800 187.035 ;
        RECT 34.970 186.735 35.705 187.215 ;
        RECT 35.875 186.645 36.045 186.995 ;
        RECT 36.215 186.815 36.595 187.215 ;
        RECT 28.670 185.100 29.020 186.350 ;
        RECT 30.785 185.925 32.435 186.445 ;
        RECT 34.490 186.395 35.225 186.565 ;
        RECT 35.875 186.475 36.615 186.645 ;
        RECT 36.785 186.540 37.055 186.885 ;
        RECT 34.975 186.305 35.225 186.395 ;
        RECT 36.445 186.305 36.615 186.475 ;
        RECT 32.605 185.755 34.295 186.275 ;
        RECT 34.470 185.975 34.805 186.225 ;
        RECT 34.975 185.975 35.715 186.305 ;
        RECT 36.445 185.975 36.675 186.305 ;
        RECT 19.745 184.665 25.090 185.100 ;
        RECT 25.265 184.665 30.610 185.100 ;
        RECT 30.785 184.665 34.295 185.755 ;
        RECT 34.470 184.665 34.725 185.805 ;
        RECT 34.975 185.415 35.145 185.975 ;
        RECT 36.445 185.805 36.615 185.975 ;
        RECT 36.885 185.805 37.055 186.540 ;
        RECT 37.250 186.565 37.560 187.035 ;
        RECT 37.730 186.735 38.465 187.215 ;
        RECT 38.635 186.645 38.805 186.995 ;
        RECT 38.975 186.815 39.355 187.215 ;
        RECT 37.250 186.395 37.985 186.565 ;
        RECT 38.635 186.475 39.375 186.645 ;
        RECT 39.545 186.540 39.815 186.885 ;
        RECT 37.735 186.305 37.985 186.395 ;
        RECT 39.205 186.305 39.375 186.475 ;
        RECT 37.230 185.975 37.565 186.225 ;
        RECT 37.735 185.975 38.475 186.305 ;
        RECT 39.205 185.975 39.435 186.305 ;
        RECT 35.370 185.635 36.615 185.805 ;
        RECT 35.370 185.385 35.790 185.635 ;
        RECT 34.920 184.885 36.115 185.215 ;
        RECT 36.295 184.665 36.575 185.465 ;
        RECT 36.785 184.835 37.055 185.805 ;
        RECT 37.230 184.665 37.485 185.805 ;
        RECT 37.735 185.415 37.905 185.975 ;
        RECT 39.205 185.805 39.375 185.975 ;
        RECT 39.645 185.805 39.815 186.540 ;
        RECT 39.985 186.395 40.245 187.215 ;
        RECT 40.415 186.395 40.745 186.815 ;
        RECT 40.925 186.645 41.185 187.045 ;
        RECT 41.355 186.815 41.685 187.215 ;
        RECT 41.855 186.645 42.025 186.995 ;
        RECT 42.195 186.815 42.570 187.215 ;
        RECT 40.925 186.475 42.590 186.645 ;
        RECT 42.760 186.540 43.035 186.885 ;
        RECT 40.495 186.305 40.745 186.395 ;
        RECT 42.420 186.305 42.590 186.475 ;
        RECT 39.990 185.975 40.325 186.225 ;
        RECT 40.495 185.975 41.210 186.305 ;
        RECT 41.425 185.975 42.250 186.305 ;
        RECT 42.420 185.975 42.695 186.305 ;
        RECT 38.130 185.635 39.375 185.805 ;
        RECT 38.130 185.385 38.550 185.635 ;
        RECT 37.680 184.885 38.875 185.215 ;
        RECT 39.055 184.665 39.335 185.465 ;
        RECT 39.545 184.835 39.815 185.805 ;
        RECT 39.985 184.665 40.245 185.805 ;
        RECT 40.495 185.415 40.665 185.975 ;
        RECT 40.925 185.515 41.255 185.805 ;
        RECT 41.425 185.685 41.670 185.975 ;
        RECT 42.420 185.805 42.590 185.975 ;
        RECT 42.865 185.805 43.035 186.540 ;
        RECT 44.125 186.490 44.415 187.215 ;
        RECT 44.585 186.475 45.075 187.045 ;
        RECT 45.245 186.645 45.475 187.045 ;
        RECT 45.645 186.815 46.065 187.215 ;
        RECT 46.235 186.645 46.405 187.045 ;
        RECT 45.245 186.475 46.405 186.645 ;
        RECT 46.575 186.475 47.025 187.215 ;
        RECT 47.195 186.475 47.635 187.035 ;
        RECT 41.930 185.635 42.590 185.805 ;
        RECT 41.930 185.515 42.100 185.635 ;
        RECT 40.925 185.345 42.100 185.515 ;
        RECT 40.485 184.845 42.100 185.175 ;
        RECT 42.270 184.665 42.550 185.465 ;
        RECT 42.760 184.835 43.035 185.805 ;
        RECT 44.125 184.665 44.415 185.830 ;
        RECT 44.585 185.805 44.755 186.475 ;
        RECT 44.925 185.975 45.330 186.305 ;
        RECT 44.585 185.635 45.355 185.805 ;
        RECT 44.595 184.665 44.925 185.465 ;
        RECT 45.105 185.005 45.355 185.635 ;
        RECT 45.545 185.175 45.795 186.305 ;
        RECT 45.995 185.975 46.240 186.305 ;
        RECT 46.425 186.025 46.815 186.305 ;
        RECT 45.995 185.175 46.195 185.975 ;
        RECT 46.985 185.855 47.155 186.305 ;
        RECT 46.365 185.685 47.155 185.855 ;
        RECT 46.365 185.005 46.535 185.685 ;
        RECT 45.105 184.835 46.535 185.005 ;
        RECT 46.705 184.665 47.020 185.515 ;
        RECT 47.325 185.465 47.635 186.475 ;
        RECT 47.195 184.835 47.635 185.465 ;
        RECT 47.805 184.835 48.085 186.935 ;
        RECT 48.315 186.755 48.485 187.215 ;
        RECT 48.755 186.825 50.005 187.005 ;
        RECT 49.140 186.585 49.505 186.655 ;
        RECT 48.255 186.405 49.505 186.585 ;
        RECT 49.675 186.605 50.005 186.825 ;
        RECT 50.175 186.775 50.345 187.215 ;
        RECT 50.515 186.605 50.855 187.020 ;
        RECT 49.675 186.435 50.855 186.605 ;
        RECT 48.255 185.805 48.530 186.405 ;
        RECT 48.700 185.975 49.055 186.225 ;
        RECT 49.250 186.195 49.715 186.225 ;
        RECT 49.245 186.025 49.715 186.195 ;
        RECT 49.250 185.975 49.715 186.025 ;
        RECT 49.885 185.975 50.215 186.225 ;
        RECT 50.390 186.025 50.855 186.225 ;
        RECT 50.035 185.855 50.215 185.975 ;
        RECT 48.255 185.595 49.865 185.805 ;
        RECT 50.035 185.685 50.365 185.855 ;
        RECT 49.455 185.495 49.865 185.595 ;
        RECT 48.275 184.665 49.060 185.425 ;
        RECT 49.455 184.835 49.840 185.495 ;
        RECT 50.165 184.895 50.365 185.685 ;
        RECT 50.535 184.665 50.855 185.845 ;
        RECT 51.075 185.680 51.405 187.045 ;
        RECT 51.575 186.830 52.250 187.215 ;
        RECT 52.525 186.650 52.855 187.040 ;
        RECT 53.025 186.815 53.370 187.215 ;
        RECT 51.635 186.645 52.855 186.650 ;
        RECT 53.540 186.645 53.745 187.040 ;
        RECT 51.635 186.475 53.745 186.645 ;
        RECT 51.635 185.835 51.855 186.475 ;
        RECT 53.925 186.455 54.480 187.015 ;
        RECT 54.655 186.540 54.895 187.215 ;
        RECT 53.925 186.305 54.230 186.455 ;
        RECT 52.230 186.010 52.660 186.250 ;
        RECT 51.075 184.840 51.330 185.680 ;
        RECT 51.635 185.655 52.285 185.835 ;
        RECT 51.505 184.665 51.835 185.485 ;
        RECT 52.075 184.840 52.285 185.655 ;
        RECT 52.455 184.835 52.660 186.010 ;
        RECT 52.830 184.835 53.160 186.250 ;
        RECT 53.340 184.835 53.620 186.305 ;
        RECT 53.845 185.975 54.230 186.305 ;
        RECT 55.165 186.445 57.755 187.215 ;
        RECT 57.950 186.565 58.260 187.035 ;
        RECT 58.430 186.735 59.165 187.215 ;
        RECT 59.335 186.645 59.505 186.995 ;
        RECT 59.675 186.815 60.055 187.215 ;
        RECT 54.450 186.010 54.950 186.275 ;
        RECT 55.165 185.925 56.375 186.445 ;
        RECT 57.950 186.395 58.685 186.565 ;
        RECT 59.335 186.475 60.075 186.645 ;
        RECT 60.245 186.540 60.515 186.885 ;
        RECT 58.435 186.305 58.685 186.395 ;
        RECT 59.905 186.305 60.075 186.475 ;
        RECT 53.800 185.635 54.930 185.805 ;
        RECT 56.545 185.755 57.755 186.275 ;
        RECT 57.930 185.975 58.265 186.225 ;
        RECT 58.435 185.975 59.175 186.305 ;
        RECT 59.905 185.975 60.135 186.305 ;
        RECT 53.800 184.840 54.085 185.635 ;
        RECT 54.265 184.665 54.480 185.465 ;
        RECT 54.660 184.840 54.930 185.635 ;
        RECT 55.165 184.665 57.755 185.755 ;
        RECT 57.930 184.665 58.185 185.805 ;
        RECT 58.435 185.415 58.605 185.975 ;
        RECT 59.905 185.805 60.075 185.975 ;
        RECT 60.345 185.805 60.515 186.540 ;
        RECT 60.685 186.445 63.275 187.215 ;
        RECT 60.685 185.925 61.895 186.445 ;
        RECT 58.830 185.635 60.075 185.805 ;
        RECT 58.830 185.385 59.250 185.635 ;
        RECT 58.380 184.885 59.575 185.215 ;
        RECT 59.755 184.665 60.035 185.465 ;
        RECT 60.245 184.835 60.515 185.805 ;
        RECT 62.065 185.755 63.275 186.275 ;
        RECT 60.685 184.665 63.275 185.755 ;
        RECT 63.905 186.230 64.175 187.045 ;
        RECT 64.345 186.475 65.015 187.215 ;
        RECT 65.185 186.645 65.480 186.990 ;
        RECT 65.660 186.815 66.035 187.215 ;
        RECT 66.250 186.645 66.580 186.990 ;
        RECT 65.185 186.475 66.580 186.645 ;
        RECT 66.830 186.475 67.415 187.045 ;
        RECT 63.905 184.835 64.255 186.230 ;
        RECT 64.425 185.805 64.595 186.305 ;
        RECT 64.765 185.975 65.100 186.305 ;
        RECT 65.270 185.975 65.610 186.305 ;
        RECT 64.425 185.635 65.170 185.805 ;
        RECT 64.425 184.665 64.830 185.465 ;
        RECT 65.000 185.005 65.170 185.635 ;
        RECT 65.340 185.230 65.610 185.975 ;
        RECT 65.800 185.975 66.090 186.305 ;
        RECT 66.260 185.975 66.660 186.305 ;
        RECT 65.800 185.230 66.035 185.975 ;
        RECT 66.830 185.805 67.000 186.475 ;
        RECT 67.645 186.395 67.855 187.215 ;
        RECT 68.025 186.415 68.355 187.045 ;
        RECT 67.170 185.975 67.415 186.305 ;
        RECT 68.025 185.815 68.275 186.415 ;
        RECT 68.525 186.395 68.755 187.215 ;
        RECT 69.885 186.490 70.175 187.215 ;
        RECT 70.345 186.445 72.935 187.215 ;
        RECT 68.445 185.975 68.775 186.225 ;
        RECT 70.345 185.925 71.555 186.445 ;
        RECT 73.380 186.405 73.625 187.010 ;
        RECT 73.845 186.680 74.355 187.215 ;
        RECT 66.205 185.635 67.415 185.805 ;
        RECT 66.205 185.005 66.535 185.635 ;
        RECT 65.000 184.835 66.535 185.005 ;
        RECT 66.720 184.665 66.955 185.465 ;
        RECT 67.125 184.835 67.415 185.635 ;
        RECT 67.645 184.665 67.855 185.805 ;
        RECT 68.025 184.835 68.355 185.815 ;
        RECT 68.525 184.665 68.755 185.805 ;
        RECT 69.885 184.665 70.175 185.830 ;
        RECT 71.725 185.755 72.935 186.275 ;
        RECT 70.345 184.665 72.935 185.755 ;
        RECT 73.105 186.235 74.335 186.405 ;
        RECT 73.105 185.425 73.445 186.235 ;
        RECT 73.615 185.670 74.365 185.860 ;
        RECT 73.105 185.015 73.620 185.425 ;
        RECT 73.855 184.665 74.025 185.425 ;
        RECT 74.195 185.005 74.365 185.670 ;
        RECT 74.535 185.685 74.725 187.045 ;
        RECT 74.895 186.875 75.170 187.045 ;
        RECT 74.895 186.705 75.175 186.875 ;
        RECT 74.895 185.885 75.170 186.705 ;
        RECT 75.360 186.680 75.890 187.045 ;
        RECT 76.315 186.815 76.645 187.215 ;
        RECT 75.715 186.645 75.890 186.680 ;
        RECT 75.375 185.685 75.545 186.485 ;
        RECT 74.535 185.515 75.545 185.685 ;
        RECT 75.715 186.475 76.645 186.645 ;
        RECT 76.815 186.475 77.070 187.045 ;
        RECT 75.715 185.345 75.885 186.475 ;
        RECT 76.475 186.305 76.645 186.475 ;
        RECT 74.760 185.175 75.885 185.345 ;
        RECT 76.055 185.975 76.250 186.305 ;
        RECT 76.475 185.975 76.730 186.305 ;
        RECT 76.055 185.005 76.225 185.975 ;
        RECT 76.900 185.805 77.070 186.475 ;
        RECT 77.335 186.565 77.505 187.045 ;
        RECT 77.675 186.735 78.005 187.215 ;
        RECT 78.230 186.795 79.765 187.045 ;
        RECT 78.230 186.565 78.400 186.795 ;
        RECT 77.335 186.395 78.400 186.565 ;
        RECT 78.580 186.225 78.860 186.625 ;
        RECT 77.250 186.015 77.600 186.225 ;
        RECT 77.770 186.025 78.215 186.225 ;
        RECT 78.385 186.025 78.860 186.225 ;
        RECT 79.130 186.225 79.415 186.625 ;
        RECT 79.595 186.565 79.765 186.795 ;
        RECT 79.935 186.735 80.265 187.215 ;
        RECT 80.480 186.715 80.735 187.045 ;
        RECT 80.525 186.705 80.735 186.715 ;
        RECT 80.550 186.635 80.735 186.705 ;
        RECT 79.595 186.395 80.395 186.565 ;
        RECT 79.130 186.025 79.460 186.225 ;
        RECT 79.630 186.025 79.995 186.225 ;
        RECT 80.225 185.845 80.395 186.395 ;
        RECT 74.195 184.835 76.225 185.005 ;
        RECT 76.395 184.665 76.565 185.805 ;
        RECT 76.735 184.835 77.070 185.805 ;
        RECT 77.335 185.675 80.395 185.845 ;
        RECT 77.335 184.835 77.505 185.675 ;
        RECT 80.565 185.505 80.735 186.635 ;
        RECT 80.925 186.465 82.135 187.215 ;
        RECT 82.395 186.665 82.565 186.955 ;
        RECT 82.735 186.835 83.065 187.215 ;
        RECT 82.395 186.495 83.060 186.665 ;
        RECT 80.925 185.925 81.445 186.465 ;
        RECT 81.615 185.755 82.135 186.295 ;
        RECT 77.675 185.005 78.005 185.505 ;
        RECT 78.175 185.265 79.810 185.505 ;
        RECT 78.175 185.175 78.405 185.265 ;
        RECT 78.515 185.005 78.845 185.045 ;
        RECT 77.675 184.835 78.845 185.005 ;
        RECT 79.035 184.665 79.390 185.085 ;
        RECT 79.560 184.835 79.810 185.265 ;
        RECT 79.980 184.665 80.310 185.425 ;
        RECT 80.480 184.835 80.735 185.505 ;
        RECT 80.925 184.665 82.135 185.755 ;
        RECT 82.310 185.675 82.660 186.325 ;
        RECT 82.830 185.505 83.060 186.495 ;
        RECT 82.395 185.335 83.060 185.505 ;
        RECT 82.395 184.835 82.565 185.335 ;
        RECT 82.735 184.665 83.065 185.165 ;
        RECT 83.235 184.835 83.460 186.955 ;
        RECT 83.675 186.755 83.925 187.215 ;
        RECT 84.110 186.765 84.440 186.935 ;
        RECT 84.620 186.765 85.370 186.935 ;
        RECT 83.660 185.635 83.940 186.235 ;
        RECT 84.110 185.235 84.280 186.765 ;
        RECT 84.450 186.265 85.030 186.595 ;
        RECT 84.450 185.395 84.690 186.265 ;
        RECT 85.200 185.985 85.370 186.765 ;
        RECT 85.620 186.715 85.990 187.215 ;
        RECT 86.170 186.765 86.630 186.935 ;
        RECT 86.860 186.765 87.530 186.935 ;
        RECT 86.170 186.535 86.340 186.765 ;
        RECT 85.540 186.235 86.340 186.535 ;
        RECT 86.510 186.265 87.060 186.595 ;
        RECT 85.540 186.205 85.710 186.235 ;
        RECT 85.830 185.985 86.000 186.055 ;
        RECT 85.200 185.815 86.000 185.985 ;
        RECT 85.490 185.725 86.000 185.815 ;
        RECT 84.880 185.290 85.320 185.645 ;
        RECT 83.660 184.665 83.925 185.125 ;
        RECT 84.110 184.860 84.345 185.235 ;
        RECT 85.490 185.110 85.660 185.725 ;
        RECT 84.590 184.940 85.660 185.110 ;
        RECT 85.830 184.665 86.000 185.465 ;
        RECT 86.170 185.165 86.340 186.235 ;
        RECT 86.510 185.335 86.700 186.055 ;
        RECT 86.870 185.725 87.060 186.265 ;
        RECT 87.360 186.225 87.530 186.765 ;
        RECT 87.845 186.685 88.015 187.215 ;
        RECT 88.310 186.565 88.670 187.005 ;
        RECT 88.845 186.735 89.015 187.215 ;
        RECT 89.205 186.570 89.540 186.995 ;
        RECT 89.715 186.740 89.885 187.215 ;
        RECT 90.060 186.570 90.395 186.995 ;
        RECT 90.565 186.740 90.735 187.215 ;
        RECT 88.310 186.395 88.810 186.565 ;
        RECT 89.205 186.400 90.875 186.570 ;
        RECT 91.045 186.465 92.255 187.215 ;
        RECT 88.640 186.225 88.810 186.395 ;
        RECT 87.360 186.055 88.450 186.225 ;
        RECT 88.640 186.055 90.460 186.225 ;
        RECT 86.870 185.395 87.190 185.725 ;
        RECT 86.170 184.835 86.420 185.165 ;
        RECT 87.360 185.135 87.530 186.055 ;
        RECT 88.640 185.800 88.810 186.055 ;
        RECT 90.630 185.835 90.875 186.400 ;
        RECT 87.700 185.630 88.810 185.800 ;
        RECT 89.205 185.665 90.875 185.835 ;
        RECT 91.045 185.755 91.565 186.295 ;
        RECT 91.735 185.925 92.255 186.465 ;
        RECT 87.700 185.470 88.560 185.630 ;
        RECT 86.645 184.965 87.530 185.135 ;
        RECT 87.710 184.665 87.925 185.165 ;
        RECT 88.390 184.845 88.560 185.470 ;
        RECT 88.845 184.665 89.025 185.445 ;
        RECT 89.205 184.905 89.540 185.665 ;
        RECT 89.720 184.665 89.890 185.495 ;
        RECT 90.060 184.905 90.390 185.665 ;
        RECT 90.560 184.665 90.730 185.495 ;
        RECT 91.045 184.665 92.255 185.755 ;
        RECT 18.280 184.495 92.340 184.665 ;
        RECT 18.365 183.405 19.575 184.495 ;
        RECT 19.745 184.060 25.090 184.495 ;
        RECT 25.265 184.060 30.610 184.495 ;
        RECT 18.365 182.695 18.885 183.235 ;
        RECT 19.055 182.865 19.575 183.405 ;
        RECT 18.365 181.945 19.575 182.695 ;
        RECT 21.330 182.490 21.670 183.320 ;
        RECT 23.150 182.810 23.500 184.060 ;
        RECT 26.850 182.490 27.190 183.320 ;
        RECT 28.670 182.810 29.020 184.060 ;
        RECT 31.245 183.330 31.535 184.495 ;
        RECT 31.705 184.060 37.050 184.495 ;
        RECT 19.745 181.945 25.090 182.490 ;
        RECT 25.265 181.945 30.610 182.490 ;
        RECT 31.245 181.945 31.535 182.670 ;
        RECT 33.290 182.490 33.630 183.320 ;
        RECT 35.110 182.810 35.460 184.060 ;
        RECT 38.235 183.875 38.405 184.305 ;
        RECT 38.575 184.045 38.905 184.495 ;
        RECT 38.235 183.645 38.910 183.875 ;
        RECT 38.205 182.625 38.505 183.475 ;
        RECT 38.675 182.995 38.910 183.645 ;
        RECT 39.080 183.335 39.365 184.280 ;
        RECT 39.545 184.025 40.230 184.495 ;
        RECT 39.540 183.505 40.235 183.815 ;
        RECT 40.410 183.440 40.715 184.225 ;
        RECT 41.915 183.750 42.185 184.495 ;
        RECT 42.815 184.490 49.090 184.495 ;
        RECT 42.355 183.580 42.645 184.320 ;
        RECT 42.815 183.765 43.070 184.490 ;
        RECT 43.255 183.595 43.515 184.320 ;
        RECT 43.685 183.765 43.930 184.490 ;
        RECT 44.115 183.595 44.375 184.320 ;
        RECT 44.545 183.765 44.790 184.490 ;
        RECT 44.975 183.595 45.235 184.320 ;
        RECT 45.405 183.765 45.650 184.490 ;
        RECT 45.820 183.595 46.080 184.320 ;
        RECT 46.250 183.765 46.510 184.490 ;
        RECT 46.680 183.595 46.940 184.320 ;
        RECT 47.110 183.765 47.370 184.490 ;
        RECT 47.540 183.595 47.800 184.320 ;
        RECT 47.970 183.765 48.230 184.490 ;
        RECT 48.400 183.595 48.660 184.320 ;
        RECT 48.830 183.695 49.090 184.490 ;
        RECT 43.255 183.580 48.660 183.595 ;
        RECT 39.080 183.185 39.940 183.335 ;
        RECT 39.080 183.165 40.365 183.185 ;
        RECT 38.675 182.665 39.210 182.995 ;
        RECT 39.380 182.805 40.365 183.165 ;
        RECT 38.675 182.515 38.895 182.665 ;
        RECT 31.705 181.945 37.050 182.490 ;
        RECT 38.150 181.945 38.485 182.450 ;
        RECT 38.655 182.140 38.895 182.515 ;
        RECT 39.380 182.470 39.550 182.805 ;
        RECT 40.540 182.635 40.715 183.440 ;
        RECT 39.175 182.275 39.550 182.470 ;
        RECT 39.175 182.130 39.345 182.275 ;
        RECT 39.910 181.945 40.305 182.440 ;
        RECT 40.475 182.115 40.715 182.635 ;
        RECT 41.915 183.355 48.660 183.580 ;
        RECT 41.915 182.765 43.080 183.355 ;
        RECT 49.260 183.185 49.510 184.320 ;
        RECT 49.690 183.685 49.950 184.495 ;
        RECT 50.125 183.185 50.370 184.325 ;
        RECT 50.550 183.685 50.845 184.495 ;
        RECT 51.025 184.060 56.370 184.495 ;
        RECT 43.250 182.935 50.370 183.185 ;
        RECT 41.915 182.595 48.660 182.765 ;
        RECT 41.915 181.945 42.215 182.425 ;
        RECT 42.385 182.140 42.645 182.595 ;
        RECT 42.815 181.945 43.075 182.425 ;
        RECT 43.255 182.140 43.515 182.595 ;
        RECT 43.685 181.945 43.935 182.425 ;
        RECT 44.115 182.140 44.375 182.595 ;
        RECT 44.545 181.945 44.795 182.425 ;
        RECT 44.975 182.140 45.235 182.595 ;
        RECT 45.405 181.945 45.650 182.425 ;
        RECT 45.820 182.140 46.095 182.595 ;
        RECT 46.265 181.945 46.510 182.425 ;
        RECT 46.680 182.140 46.940 182.595 ;
        RECT 47.110 181.945 47.370 182.425 ;
        RECT 47.540 182.140 47.800 182.595 ;
        RECT 47.970 181.945 48.230 182.425 ;
        RECT 48.400 182.140 48.660 182.595 ;
        RECT 48.830 181.945 49.090 182.505 ;
        RECT 49.260 182.125 49.510 182.935 ;
        RECT 49.690 181.945 49.950 182.470 ;
        RECT 50.120 182.125 50.370 182.935 ;
        RECT 50.540 182.625 50.855 183.185 ;
        RECT 52.610 182.490 52.950 183.320 ;
        RECT 54.430 182.810 54.780 184.060 ;
        RECT 57.005 183.330 57.295 184.495 ;
        RECT 57.465 184.060 62.810 184.495 ;
        RECT 50.550 181.945 50.855 182.455 ;
        RECT 51.025 181.945 56.370 182.490 ;
        RECT 57.005 181.945 57.295 182.670 ;
        RECT 59.050 182.490 59.390 183.320 ;
        RECT 60.870 182.810 61.220 184.060 ;
        RECT 62.985 183.405 64.195 184.495 ;
        RECT 64.665 183.855 64.995 184.285 ;
        RECT 62.985 182.695 63.505 183.235 ;
        RECT 63.675 182.865 64.195 183.405 ;
        RECT 64.540 183.685 64.995 183.855 ;
        RECT 65.175 183.855 65.425 184.275 ;
        RECT 65.655 184.025 65.985 184.495 ;
        RECT 66.215 183.855 66.465 184.275 ;
        RECT 65.175 183.685 66.465 183.855 ;
        RECT 57.465 181.945 62.810 182.490 ;
        RECT 62.985 181.945 64.195 182.695 ;
        RECT 64.540 182.685 64.710 183.685 ;
        RECT 64.880 182.855 65.125 183.515 ;
        RECT 65.340 182.855 65.605 183.515 ;
        RECT 65.800 182.855 66.085 183.515 ;
        RECT 66.260 183.185 66.475 183.515 ;
        RECT 66.655 183.355 66.905 184.495 ;
        RECT 67.075 183.435 67.405 184.285 ;
        RECT 67.595 183.685 67.890 184.495 ;
        RECT 66.260 182.855 66.565 183.185 ;
        RECT 66.735 182.855 67.045 183.185 ;
        RECT 66.735 182.685 66.905 182.855 ;
        RECT 64.540 182.515 66.905 182.685 ;
        RECT 67.215 182.670 67.405 183.435 ;
        RECT 68.070 183.185 68.315 184.325 ;
        RECT 68.490 183.685 68.750 184.495 ;
        RECT 69.350 184.490 75.625 184.495 ;
        RECT 68.930 183.185 69.180 184.320 ;
        RECT 69.350 183.695 69.610 184.490 ;
        RECT 69.780 183.595 70.040 184.320 ;
        RECT 70.210 183.765 70.470 184.490 ;
        RECT 70.640 183.595 70.900 184.320 ;
        RECT 71.070 183.765 71.330 184.490 ;
        RECT 71.500 183.595 71.760 184.320 ;
        RECT 71.930 183.765 72.190 184.490 ;
        RECT 72.360 183.595 72.620 184.320 ;
        RECT 72.790 183.765 73.035 184.490 ;
        RECT 73.205 183.595 73.465 184.320 ;
        RECT 73.650 183.765 73.895 184.490 ;
        RECT 74.065 183.595 74.325 184.320 ;
        RECT 74.510 183.765 74.755 184.490 ;
        RECT 74.925 183.595 75.185 184.320 ;
        RECT 75.370 183.765 75.625 184.490 ;
        RECT 69.780 183.580 75.185 183.595 ;
        RECT 75.795 183.580 76.085 184.320 ;
        RECT 76.255 183.750 76.525 184.495 ;
        RECT 69.780 183.355 76.525 183.580 ;
        RECT 76.785 183.405 78.455 184.495 ;
        RECT 64.695 181.945 65.025 182.345 ;
        RECT 65.195 182.175 65.525 182.515 ;
        RECT 66.575 181.945 66.905 182.345 ;
        RECT 67.075 182.160 67.405 182.670 ;
        RECT 67.585 182.625 67.900 183.185 ;
        RECT 68.070 182.935 75.190 183.185 ;
        RECT 67.585 181.945 67.890 182.455 ;
        RECT 68.070 182.125 68.320 182.935 ;
        RECT 68.490 181.945 68.750 182.470 ;
        RECT 68.930 182.125 69.180 182.935 ;
        RECT 75.360 182.795 76.525 183.355 ;
        RECT 75.360 182.765 76.555 182.795 ;
        RECT 69.780 182.625 76.555 182.765 ;
        RECT 76.785 182.715 77.535 183.235 ;
        RECT 77.705 182.885 78.455 183.405 ;
        RECT 69.780 182.595 76.525 182.625 ;
        RECT 69.350 181.945 69.610 182.505 ;
        RECT 69.780 182.140 70.040 182.595 ;
        RECT 70.210 181.945 70.470 182.425 ;
        RECT 70.640 182.140 70.900 182.595 ;
        RECT 71.070 181.945 71.330 182.425 ;
        RECT 71.500 182.140 71.760 182.595 ;
        RECT 71.930 181.945 72.175 182.425 ;
        RECT 72.345 182.140 72.620 182.595 ;
        RECT 72.790 181.945 73.035 182.425 ;
        RECT 73.205 182.140 73.465 182.595 ;
        RECT 73.645 181.945 73.895 182.425 ;
        RECT 74.065 182.140 74.325 182.595 ;
        RECT 74.505 181.945 74.755 182.425 ;
        RECT 74.925 182.140 75.185 182.595 ;
        RECT 75.365 181.945 75.625 182.425 ;
        RECT 75.795 182.140 76.055 182.595 ;
        RECT 76.225 181.945 76.525 182.425 ;
        RECT 76.785 181.945 78.455 182.715 ;
        RECT 78.635 182.125 78.895 184.315 ;
        RECT 79.065 183.765 79.405 184.495 ;
        RECT 79.585 183.585 79.855 184.315 ;
        RECT 79.085 183.365 79.855 183.585 ;
        RECT 80.035 183.605 80.265 184.315 ;
        RECT 80.435 183.785 80.765 184.495 ;
        RECT 80.935 183.605 81.195 184.315 ;
        RECT 80.035 183.365 81.195 183.605 ;
        RECT 79.085 182.695 79.375 183.365 ;
        RECT 81.385 183.355 81.645 184.495 ;
        RECT 81.815 183.345 82.145 184.325 ;
        RECT 82.315 183.355 82.595 184.495 ;
        RECT 79.555 182.875 80.020 183.185 ;
        RECT 80.200 182.875 80.725 183.185 ;
        RECT 79.085 182.495 80.315 182.695 ;
        RECT 79.155 181.945 79.825 182.315 ;
        RECT 80.005 182.125 80.315 182.495 ;
        RECT 80.495 182.235 80.725 182.875 ;
        RECT 80.905 182.855 81.205 183.185 ;
        RECT 81.405 182.935 81.740 183.185 ;
        RECT 81.910 182.745 82.080 183.345 ;
        RECT 82.765 183.330 83.055 184.495 ;
        RECT 83.225 184.060 88.570 184.495 ;
        RECT 82.250 182.915 82.585 183.185 ;
        RECT 80.905 181.945 81.195 182.675 ;
        RECT 81.385 182.115 82.080 182.745 ;
        RECT 82.285 181.945 82.595 182.745 ;
        RECT 82.765 181.945 83.055 182.670 ;
        RECT 84.810 182.490 85.150 183.320 ;
        RECT 86.630 182.810 86.980 184.060 ;
        RECT 88.745 183.405 90.415 184.495 ;
        RECT 88.745 182.715 89.495 183.235 ;
        RECT 89.665 182.885 90.415 183.405 ;
        RECT 91.045 183.405 92.255 184.495 ;
        RECT 91.045 182.865 91.565 183.405 ;
        RECT 83.225 181.945 88.570 182.490 ;
        RECT 88.745 181.945 90.415 182.715 ;
        RECT 91.735 182.695 92.255 183.235 ;
        RECT 91.045 181.945 92.255 182.695 ;
        RECT 18.280 181.775 92.340 181.945 ;
        RECT 18.365 181.025 19.575 181.775 ;
        RECT 19.745 181.230 25.090 181.775 ;
        RECT 25.265 181.230 30.610 181.775 ;
        RECT 30.785 181.230 36.130 181.775 ;
        RECT 18.365 180.485 18.885 181.025 ;
        RECT 19.055 180.315 19.575 180.855 ;
        RECT 21.330 180.400 21.670 181.230 ;
        RECT 18.365 179.225 19.575 180.315 ;
        RECT 23.150 179.660 23.500 180.910 ;
        RECT 26.850 180.400 27.190 181.230 ;
        RECT 28.670 179.660 29.020 180.910 ;
        RECT 32.370 180.400 32.710 181.230 ;
        RECT 36.305 181.005 39.815 181.775 ;
        RECT 39.985 181.025 41.195 181.775 ;
        RECT 34.190 179.660 34.540 180.910 ;
        RECT 36.305 180.485 37.955 181.005 ;
        RECT 38.125 180.315 39.815 180.835 ;
        RECT 39.985 180.485 40.505 181.025 ;
        RECT 41.375 180.965 41.645 181.775 ;
        RECT 41.815 180.965 42.145 181.605 ;
        RECT 42.315 180.965 42.555 181.775 ;
        RECT 42.745 181.025 43.955 181.775 ;
        RECT 44.125 181.050 44.415 181.775 ;
        RECT 44.585 181.275 44.885 181.605 ;
        RECT 45.055 181.295 45.330 181.775 ;
        RECT 40.675 180.315 41.195 180.855 ;
        RECT 41.365 180.535 41.715 180.785 ;
        RECT 41.885 180.365 42.055 180.965 ;
        RECT 42.225 180.535 42.575 180.785 ;
        RECT 42.745 180.485 43.265 181.025 ;
        RECT 19.745 179.225 25.090 179.660 ;
        RECT 25.265 179.225 30.610 179.660 ;
        RECT 30.785 179.225 36.130 179.660 ;
        RECT 36.305 179.225 39.815 180.315 ;
        RECT 39.985 179.225 41.195 180.315 ;
        RECT 41.375 179.225 41.705 180.365 ;
        RECT 41.885 180.195 42.565 180.365 ;
        RECT 43.435 180.315 43.955 180.855 ;
        RECT 42.235 179.410 42.565 180.195 ;
        RECT 42.745 179.225 43.955 180.315 ;
        RECT 44.125 179.225 44.415 180.390 ;
        RECT 44.585 180.365 44.755 181.275 ;
        RECT 45.510 181.125 45.805 181.515 ;
        RECT 45.975 181.295 46.230 181.775 ;
        RECT 46.405 181.125 46.665 181.515 ;
        RECT 46.835 181.295 47.115 181.775 ;
        RECT 44.925 180.535 45.275 181.105 ;
        RECT 45.510 180.955 47.160 181.125 ;
        RECT 47.405 180.955 47.615 181.775 ;
        RECT 47.785 180.975 48.115 181.605 ;
        RECT 45.445 180.615 46.585 180.785 ;
        RECT 45.445 180.365 45.615 180.615 ;
        RECT 46.755 180.445 47.160 180.955 ;
        RECT 44.585 180.195 45.615 180.365 ;
        RECT 46.405 180.275 47.160 180.445 ;
        RECT 47.785 180.375 48.035 180.975 ;
        RECT 48.285 180.955 48.515 181.775 ;
        RECT 48.725 181.005 51.315 181.775 ;
        RECT 48.205 180.535 48.535 180.785 ;
        RECT 48.725 180.485 49.935 181.005 ;
        RECT 52.005 180.955 52.215 181.775 ;
        RECT 52.385 180.975 52.715 181.605 ;
        RECT 44.585 179.395 44.895 180.195 ;
        RECT 46.405 180.025 46.665 180.275 ;
        RECT 45.065 179.225 45.375 180.025 ;
        RECT 45.545 179.855 46.665 180.025 ;
        RECT 45.545 179.395 45.805 179.855 ;
        RECT 45.975 179.225 46.230 179.685 ;
        RECT 46.405 179.395 46.665 179.855 ;
        RECT 46.835 179.225 47.120 180.095 ;
        RECT 47.405 179.225 47.615 180.365 ;
        RECT 47.785 179.395 48.115 180.375 ;
        RECT 48.285 179.225 48.515 180.365 ;
        RECT 50.105 180.315 51.315 180.835 ;
        RECT 52.385 180.375 52.635 180.975 ;
        RECT 52.885 180.955 53.115 181.775 ;
        RECT 53.385 180.955 53.595 181.775 ;
        RECT 53.765 180.975 54.095 181.605 ;
        RECT 52.805 180.535 53.135 180.785 ;
        RECT 53.765 180.375 54.015 180.975 ;
        RECT 54.265 180.955 54.495 181.775 ;
        RECT 54.705 181.005 57.295 181.775 ;
        RECT 57.945 181.045 58.235 181.775 ;
        RECT 54.185 180.535 54.515 180.785 ;
        RECT 54.705 180.485 55.915 181.005 ;
        RECT 48.725 179.225 51.315 180.315 ;
        RECT 52.005 179.225 52.215 180.365 ;
        RECT 52.385 179.395 52.715 180.375 ;
        RECT 52.885 179.225 53.115 180.365 ;
        RECT 53.385 179.225 53.595 180.365 ;
        RECT 53.765 179.395 54.095 180.375 ;
        RECT 54.265 179.225 54.495 180.365 ;
        RECT 56.085 180.315 57.295 180.835 ;
        RECT 57.935 180.535 58.235 180.865 ;
        RECT 58.415 180.845 58.645 181.485 ;
        RECT 58.825 181.225 59.135 181.595 ;
        RECT 59.315 181.405 59.985 181.775 ;
        RECT 58.825 181.025 60.055 181.225 ;
        RECT 58.415 180.535 58.940 180.845 ;
        RECT 59.120 180.535 59.585 180.845 ;
        RECT 59.765 180.355 60.055 181.025 ;
        RECT 54.705 179.225 57.295 180.315 ;
        RECT 57.945 180.115 59.105 180.355 ;
        RECT 57.945 179.405 58.205 180.115 ;
        RECT 58.375 179.225 58.705 179.935 ;
        RECT 58.875 179.405 59.105 180.115 ;
        RECT 59.285 180.135 60.055 180.355 ;
        RECT 59.285 179.405 59.555 180.135 ;
        RECT 59.735 179.225 60.075 179.955 ;
        RECT 60.245 179.405 60.505 181.595 ;
        RECT 60.890 180.995 61.390 181.605 ;
        RECT 60.685 180.535 61.035 180.785 ;
        RECT 61.220 180.365 61.390 180.995 ;
        RECT 62.020 181.125 62.350 181.605 ;
        RECT 62.520 181.315 62.745 181.775 ;
        RECT 62.915 181.125 63.245 181.605 ;
        RECT 62.020 180.955 63.245 181.125 ;
        RECT 63.435 180.975 63.685 181.775 ;
        RECT 63.855 180.975 64.195 181.605 ;
        RECT 64.375 181.045 64.675 181.775 ;
        RECT 61.560 180.585 61.890 180.785 ;
        RECT 62.060 180.585 62.390 180.785 ;
        RECT 62.560 180.585 62.980 180.785 ;
        RECT 63.155 180.615 63.850 180.785 ;
        RECT 63.155 180.365 63.325 180.615 ;
        RECT 64.020 180.365 64.195 180.975 ;
        RECT 64.855 180.865 65.085 181.485 ;
        RECT 65.285 181.215 65.510 181.595 ;
        RECT 65.680 181.385 66.010 181.775 ;
        RECT 65.285 181.035 65.615 181.215 ;
        RECT 64.380 180.535 64.675 180.865 ;
        RECT 64.855 180.535 65.270 180.865 ;
        RECT 60.890 180.195 63.325 180.365 ;
        RECT 60.890 179.395 61.220 180.195 ;
        RECT 61.390 179.225 61.720 180.025 ;
        RECT 62.020 179.395 62.350 180.195 ;
        RECT 62.995 179.225 63.245 180.025 ;
        RECT 63.515 179.225 63.685 180.365 ;
        RECT 63.855 179.395 64.195 180.365 ;
        RECT 65.440 180.365 65.615 181.035 ;
        RECT 65.785 180.535 66.025 181.185 ;
        RECT 66.205 181.005 69.715 181.775 ;
        RECT 69.885 181.050 70.175 181.775 ;
        RECT 70.345 181.025 71.555 181.775 ;
        RECT 71.725 181.275 72.025 181.605 ;
        RECT 72.195 181.295 72.470 181.775 ;
        RECT 66.205 180.485 67.855 181.005 ;
        RECT 64.375 180.005 65.270 180.335 ;
        RECT 65.440 180.175 66.025 180.365 ;
        RECT 68.025 180.315 69.715 180.835 ;
        RECT 70.345 180.485 70.865 181.025 ;
        RECT 64.375 179.835 65.580 180.005 ;
        RECT 64.375 179.405 64.705 179.835 ;
        RECT 64.885 179.225 65.080 179.665 ;
        RECT 65.250 179.405 65.580 179.835 ;
        RECT 65.750 179.405 66.025 180.175 ;
        RECT 66.205 179.225 69.715 180.315 ;
        RECT 69.885 179.225 70.175 180.390 ;
        RECT 71.035 180.315 71.555 180.855 ;
        RECT 70.345 179.225 71.555 180.315 ;
        RECT 71.725 180.365 71.895 181.275 ;
        RECT 72.650 181.125 72.945 181.515 ;
        RECT 73.115 181.295 73.370 181.775 ;
        RECT 73.545 181.125 73.805 181.515 ;
        RECT 73.975 181.295 74.255 181.775 ;
        RECT 72.065 180.535 72.415 181.105 ;
        RECT 72.650 180.955 74.300 181.125 ;
        RECT 72.585 180.615 73.725 180.785 ;
        RECT 72.585 180.365 72.755 180.615 ;
        RECT 73.895 180.445 74.300 180.955 ;
        RECT 74.485 181.005 76.155 181.775 ;
        RECT 76.945 181.215 77.275 181.605 ;
        RECT 77.445 181.385 78.630 181.555 ;
        RECT 78.890 181.305 79.060 181.775 ;
        RECT 76.945 181.035 77.455 181.215 ;
        RECT 74.485 180.485 75.235 181.005 ;
        RECT 71.725 180.195 72.755 180.365 ;
        RECT 73.545 180.275 74.300 180.445 ;
        RECT 75.405 180.315 76.155 180.835 ;
        RECT 76.785 180.575 77.115 180.865 ;
        RECT 77.285 180.405 77.455 181.035 ;
        RECT 77.860 181.125 78.245 181.215 ;
        RECT 79.230 181.125 79.560 181.590 ;
        RECT 77.860 180.955 79.560 181.125 ;
        RECT 79.730 180.955 79.900 181.775 ;
        RECT 80.070 180.955 80.755 181.595 ;
        RECT 80.935 180.965 81.205 181.775 ;
        RECT 81.375 180.965 81.705 181.605 ;
        RECT 81.875 180.965 82.115 181.775 ;
        RECT 82.395 181.225 82.565 181.515 ;
        RECT 82.735 181.395 83.065 181.775 ;
        RECT 82.395 181.055 83.060 181.225 ;
        RECT 77.625 180.575 77.955 180.785 ;
        RECT 78.135 180.535 78.515 180.785 ;
        RECT 71.725 179.395 72.035 180.195 ;
        RECT 73.545 180.025 73.805 180.275 ;
        RECT 72.205 179.225 72.515 180.025 ;
        RECT 72.685 179.855 73.805 180.025 ;
        RECT 72.685 179.395 72.945 179.855 ;
        RECT 73.115 179.225 73.370 179.685 ;
        RECT 73.545 179.395 73.805 179.855 ;
        RECT 73.975 179.225 74.260 180.095 ;
        RECT 74.485 179.225 76.155 180.315 ;
        RECT 76.940 180.235 78.025 180.405 ;
        RECT 76.940 179.395 77.240 180.235 ;
        RECT 77.435 179.225 77.685 180.065 ;
        RECT 77.855 179.985 78.025 180.235 ;
        RECT 78.195 180.155 78.515 180.535 ;
        RECT 78.705 180.575 79.190 180.785 ;
        RECT 79.380 180.575 79.830 180.785 ;
        RECT 80.000 180.575 80.335 180.785 ;
        RECT 78.705 180.415 79.080 180.575 ;
        RECT 78.685 180.245 79.080 180.415 ;
        RECT 80.000 180.405 80.170 180.575 ;
        RECT 78.705 180.155 79.080 180.245 ;
        RECT 79.250 180.235 80.170 180.405 ;
        RECT 79.250 179.985 79.420 180.235 ;
        RECT 77.855 179.815 79.420 179.985 ;
        RECT 78.275 179.395 79.080 179.815 ;
        RECT 79.590 179.225 79.920 180.065 ;
        RECT 80.505 179.985 80.755 180.955 ;
        RECT 80.925 180.535 81.275 180.785 ;
        RECT 81.445 180.365 81.615 180.965 ;
        RECT 81.785 180.535 82.135 180.785 ;
        RECT 80.090 179.395 80.755 179.985 ;
        RECT 80.935 179.225 81.265 180.365 ;
        RECT 81.445 180.195 82.125 180.365 ;
        RECT 82.310 180.235 82.660 180.885 ;
        RECT 81.795 179.410 82.125 180.195 ;
        RECT 82.830 180.065 83.060 181.055 ;
        RECT 82.395 179.895 83.060 180.065 ;
        RECT 82.395 179.395 82.565 179.895 ;
        RECT 82.735 179.225 83.065 179.725 ;
        RECT 83.235 179.395 83.460 181.515 ;
        RECT 83.675 181.315 83.925 181.775 ;
        RECT 84.110 181.325 84.440 181.495 ;
        RECT 84.620 181.325 85.370 181.495 ;
        RECT 83.660 180.195 83.940 180.795 ;
        RECT 84.110 179.795 84.280 181.325 ;
        RECT 84.450 180.825 85.030 181.155 ;
        RECT 84.450 179.955 84.690 180.825 ;
        RECT 85.200 180.545 85.370 181.325 ;
        RECT 85.620 181.275 85.990 181.775 ;
        RECT 86.170 181.325 86.630 181.495 ;
        RECT 86.860 181.325 87.530 181.495 ;
        RECT 86.170 181.095 86.340 181.325 ;
        RECT 85.540 180.795 86.340 181.095 ;
        RECT 86.510 180.825 87.060 181.155 ;
        RECT 85.540 180.765 85.710 180.795 ;
        RECT 85.830 180.545 86.000 180.615 ;
        RECT 85.200 180.375 86.000 180.545 ;
        RECT 85.490 180.285 86.000 180.375 ;
        RECT 84.880 179.850 85.320 180.205 ;
        RECT 83.660 179.225 83.925 179.685 ;
        RECT 84.110 179.420 84.345 179.795 ;
        RECT 85.490 179.670 85.660 180.285 ;
        RECT 84.590 179.500 85.660 179.670 ;
        RECT 85.830 179.225 86.000 180.025 ;
        RECT 86.170 179.725 86.340 180.795 ;
        RECT 86.510 179.895 86.700 180.615 ;
        RECT 86.870 180.285 87.060 180.825 ;
        RECT 87.360 180.785 87.530 181.325 ;
        RECT 87.845 181.245 88.015 181.775 ;
        RECT 88.310 181.125 88.670 181.565 ;
        RECT 88.845 181.295 89.015 181.775 ;
        RECT 89.205 181.130 89.540 181.555 ;
        RECT 89.715 181.300 89.885 181.775 ;
        RECT 90.060 181.130 90.395 181.555 ;
        RECT 90.565 181.300 90.735 181.775 ;
        RECT 88.310 180.955 88.810 181.125 ;
        RECT 89.205 180.960 90.875 181.130 ;
        RECT 91.045 181.025 92.255 181.775 ;
        RECT 88.640 180.785 88.810 180.955 ;
        RECT 87.360 180.615 88.450 180.785 ;
        RECT 88.640 180.615 90.460 180.785 ;
        RECT 86.870 179.955 87.190 180.285 ;
        RECT 86.170 179.395 86.420 179.725 ;
        RECT 87.360 179.695 87.530 180.615 ;
        RECT 88.640 180.360 88.810 180.615 ;
        RECT 90.630 180.395 90.875 180.960 ;
        RECT 87.700 180.190 88.810 180.360 ;
        RECT 89.205 180.225 90.875 180.395 ;
        RECT 91.045 180.315 91.565 180.855 ;
        RECT 91.735 180.485 92.255 181.025 ;
        RECT 87.700 180.030 88.560 180.190 ;
        RECT 86.645 179.525 87.530 179.695 ;
        RECT 87.710 179.225 87.925 179.725 ;
        RECT 88.390 179.405 88.560 180.030 ;
        RECT 88.845 179.225 89.025 180.005 ;
        RECT 89.205 179.465 89.540 180.225 ;
        RECT 89.720 179.225 89.890 180.055 ;
        RECT 90.060 179.465 90.390 180.225 ;
        RECT 90.560 179.225 90.730 180.055 ;
        RECT 91.045 179.225 92.255 180.315 ;
        RECT 18.280 179.055 92.340 179.225 ;
        RECT 18.365 177.965 19.575 179.055 ;
        RECT 19.745 178.620 25.090 179.055 ;
        RECT 25.265 178.620 30.610 179.055 ;
        RECT 18.365 177.255 18.885 177.795 ;
        RECT 19.055 177.425 19.575 177.965 ;
        RECT 18.365 176.505 19.575 177.255 ;
        RECT 21.330 177.050 21.670 177.880 ;
        RECT 23.150 177.370 23.500 178.620 ;
        RECT 26.850 177.050 27.190 177.880 ;
        RECT 28.670 177.370 29.020 178.620 ;
        RECT 31.245 177.890 31.535 179.055 ;
        RECT 31.705 178.620 37.050 179.055 ;
        RECT 19.745 176.505 25.090 177.050 ;
        RECT 25.265 176.505 30.610 177.050 ;
        RECT 31.245 176.505 31.535 177.230 ;
        RECT 33.290 177.050 33.630 177.880 ;
        RECT 35.110 177.370 35.460 178.620 ;
        RECT 37.225 177.965 39.815 179.055 ;
        RECT 40.075 178.385 40.245 178.885 ;
        RECT 40.415 178.555 40.745 179.055 ;
        RECT 40.075 178.215 40.740 178.385 ;
        RECT 37.225 177.275 38.435 177.795 ;
        RECT 38.605 177.445 39.815 177.965 ;
        RECT 39.990 177.395 40.340 178.045 ;
        RECT 31.705 176.505 37.050 177.050 ;
        RECT 37.225 176.505 39.815 177.275 ;
        RECT 40.510 177.225 40.740 178.215 ;
        RECT 40.075 177.055 40.740 177.225 ;
        RECT 40.075 176.765 40.245 177.055 ;
        RECT 40.415 176.505 40.745 176.885 ;
        RECT 40.915 176.765 41.100 178.885 ;
        RECT 41.340 178.595 41.605 179.055 ;
        RECT 41.775 178.460 42.025 178.885 ;
        RECT 42.235 178.610 43.340 178.780 ;
        RECT 41.720 178.330 42.025 178.460 ;
        RECT 41.270 177.135 41.550 178.085 ;
        RECT 41.720 177.225 41.890 178.330 ;
        RECT 42.060 177.545 42.300 178.140 ;
        RECT 42.470 178.075 43.000 178.440 ;
        RECT 42.470 177.375 42.640 178.075 ;
        RECT 43.170 177.995 43.340 178.610 ;
        RECT 43.510 178.255 43.680 179.055 ;
        RECT 43.850 178.555 44.100 178.885 ;
        RECT 44.325 178.585 45.210 178.755 ;
        RECT 43.170 177.905 43.680 177.995 ;
        RECT 41.720 177.095 41.945 177.225 ;
        RECT 42.115 177.155 42.640 177.375 ;
        RECT 42.810 177.735 43.680 177.905 ;
        RECT 41.355 176.505 41.605 176.965 ;
        RECT 41.775 176.955 41.945 177.095 ;
        RECT 42.810 176.955 42.980 177.735 ;
        RECT 43.510 177.665 43.680 177.735 ;
        RECT 43.190 177.485 43.390 177.515 ;
        RECT 43.850 177.485 44.020 178.555 ;
        RECT 44.190 177.665 44.380 178.385 ;
        RECT 43.190 177.185 44.020 177.485 ;
        RECT 44.550 177.455 44.870 178.415 ;
        RECT 41.775 176.785 42.110 176.955 ;
        RECT 42.305 176.785 42.980 176.955 ;
        RECT 43.300 176.505 43.670 177.005 ;
        RECT 43.850 176.955 44.020 177.185 ;
        RECT 44.405 177.125 44.870 177.455 ;
        RECT 45.040 177.745 45.210 178.585 ;
        RECT 45.390 178.555 45.705 179.055 ;
        RECT 45.935 178.325 46.275 178.885 ;
        RECT 45.380 177.950 46.275 178.325 ;
        RECT 46.445 178.045 46.615 179.055 ;
        RECT 46.085 177.745 46.275 177.950 ;
        RECT 46.785 177.995 47.115 178.840 ;
        RECT 46.785 177.915 47.175 177.995 ;
        RECT 47.345 177.965 49.015 179.055 ;
        RECT 46.960 177.865 47.175 177.915 ;
        RECT 45.040 177.415 45.915 177.745 ;
        RECT 46.085 177.415 46.835 177.745 ;
        RECT 45.040 176.955 45.210 177.415 ;
        RECT 46.085 177.245 46.285 177.415 ;
        RECT 47.005 177.285 47.175 177.865 ;
        RECT 46.950 177.245 47.175 177.285 ;
        RECT 43.850 176.785 44.255 176.955 ;
        RECT 44.425 176.785 45.210 176.955 ;
        RECT 45.485 176.505 45.695 177.035 ;
        RECT 45.955 176.720 46.285 177.245 ;
        RECT 46.795 177.160 47.175 177.245 ;
        RECT 47.345 177.275 48.095 177.795 ;
        RECT 48.265 177.445 49.015 177.965 ;
        RECT 49.185 177.915 49.570 178.875 ;
        RECT 49.785 178.255 50.075 179.055 ;
        RECT 50.245 178.715 51.610 178.885 ;
        RECT 50.245 178.085 50.415 178.715 ;
        RECT 49.740 177.915 50.415 178.085 ;
        RECT 46.455 176.505 46.625 177.115 ;
        RECT 46.795 176.725 47.125 177.160 ;
        RECT 47.345 176.505 49.015 177.275 ;
        RECT 49.185 177.245 49.360 177.915 ;
        RECT 49.740 177.745 49.910 177.915 ;
        RECT 50.585 177.745 50.910 178.545 ;
        RECT 51.280 178.505 51.610 178.715 ;
        RECT 51.280 178.255 52.235 178.505 ;
        RECT 49.545 177.495 49.910 177.745 ;
        RECT 50.105 177.495 50.355 177.745 ;
        RECT 49.545 177.415 49.735 177.495 ;
        RECT 50.105 177.415 50.275 177.495 ;
        RECT 50.565 177.415 50.910 177.745 ;
        RECT 51.080 177.415 51.355 178.080 ;
        RECT 51.540 177.415 51.895 178.080 ;
        RECT 52.065 177.245 52.235 178.255 ;
        RECT 52.405 177.915 52.695 179.055 ;
        RECT 53.325 178.185 53.600 178.885 ;
        RECT 53.770 178.510 54.025 179.055 ;
        RECT 54.195 178.545 54.675 178.885 ;
        RECT 54.850 178.500 55.455 179.055 ;
        RECT 54.840 178.400 55.455 178.500 ;
        RECT 54.840 178.375 55.025 178.400 ;
        RECT 52.420 177.415 52.695 177.745 ;
        RECT 49.185 176.675 49.695 177.245 ;
        RECT 50.240 177.075 51.640 177.245 ;
        RECT 49.865 176.505 50.035 177.065 ;
        RECT 50.240 176.675 50.570 177.075 ;
        RECT 50.745 176.505 51.075 176.905 ;
        RECT 51.310 176.885 51.640 177.075 ;
        RECT 51.810 177.055 52.235 177.245 ;
        RECT 53.325 177.155 53.495 178.185 ;
        RECT 53.770 178.055 54.525 178.305 ;
        RECT 54.695 178.130 55.025 178.375 ;
        RECT 53.770 178.020 54.540 178.055 ;
        RECT 53.770 178.010 54.555 178.020 ;
        RECT 53.665 177.995 54.560 178.010 ;
        RECT 53.665 177.980 54.580 177.995 ;
        RECT 53.665 177.970 54.600 177.980 ;
        RECT 53.665 177.960 54.625 177.970 ;
        RECT 53.665 177.930 54.695 177.960 ;
        RECT 53.665 177.900 54.715 177.930 ;
        RECT 53.665 177.870 54.735 177.900 ;
        RECT 53.665 177.845 54.765 177.870 ;
        RECT 53.665 177.810 54.800 177.845 ;
        RECT 53.665 177.805 54.830 177.810 ;
        RECT 53.665 177.410 53.895 177.805 ;
        RECT 54.440 177.800 54.830 177.805 ;
        RECT 54.465 177.790 54.830 177.800 ;
        RECT 54.480 177.785 54.830 177.790 ;
        RECT 54.495 177.780 54.830 177.785 ;
        RECT 55.195 177.780 55.455 178.230 ;
        RECT 55.625 177.965 56.835 179.055 ;
        RECT 54.495 177.775 55.455 177.780 ;
        RECT 54.505 177.765 55.455 177.775 ;
        RECT 54.515 177.760 55.455 177.765 ;
        RECT 54.525 177.750 55.455 177.760 ;
        RECT 54.530 177.740 55.455 177.750 ;
        RECT 54.535 177.735 55.455 177.740 ;
        RECT 54.545 177.720 55.455 177.735 ;
        RECT 54.550 177.705 55.455 177.720 ;
        RECT 54.560 177.680 55.455 177.705 ;
        RECT 54.065 177.210 54.395 177.635 ;
        RECT 52.405 176.885 52.695 177.155 ;
        RECT 51.310 176.675 52.695 176.885 ;
        RECT 53.325 176.675 53.585 177.155 ;
        RECT 53.755 176.505 54.005 177.045 ;
        RECT 54.175 176.725 54.395 177.210 ;
        RECT 54.565 177.610 55.455 177.680 ;
        RECT 54.565 176.885 54.735 177.610 ;
        RECT 54.905 177.055 55.455 177.440 ;
        RECT 55.625 177.255 56.145 177.795 ;
        RECT 56.315 177.425 56.835 177.965 ;
        RECT 57.005 177.890 57.295 179.055 ;
        RECT 57.465 178.500 58.070 179.055 ;
        RECT 58.245 178.545 58.725 178.885 ;
        RECT 58.895 178.510 59.150 179.055 ;
        RECT 57.465 178.400 58.080 178.500 ;
        RECT 57.895 178.375 58.080 178.400 ;
        RECT 57.465 177.780 57.725 178.230 ;
        RECT 57.895 178.130 58.225 178.375 ;
        RECT 58.395 178.055 59.150 178.305 ;
        RECT 59.320 178.185 59.595 178.885 ;
        RECT 58.380 178.020 59.150 178.055 ;
        RECT 58.365 178.010 59.150 178.020 ;
        RECT 58.360 177.995 59.255 178.010 ;
        RECT 58.340 177.980 59.255 177.995 ;
        RECT 58.320 177.970 59.255 177.980 ;
        RECT 58.295 177.960 59.255 177.970 ;
        RECT 58.225 177.930 59.255 177.960 ;
        RECT 58.205 177.900 59.255 177.930 ;
        RECT 58.185 177.870 59.255 177.900 ;
        RECT 58.155 177.845 59.255 177.870 ;
        RECT 58.120 177.810 59.255 177.845 ;
        RECT 58.090 177.805 59.255 177.810 ;
        RECT 58.090 177.800 58.480 177.805 ;
        RECT 58.090 177.790 58.455 177.800 ;
        RECT 58.090 177.785 58.440 177.790 ;
        RECT 58.090 177.780 58.425 177.785 ;
        RECT 57.465 177.775 58.425 177.780 ;
        RECT 57.465 177.765 58.415 177.775 ;
        RECT 57.465 177.760 58.405 177.765 ;
        RECT 57.465 177.750 58.395 177.760 ;
        RECT 57.465 177.740 58.390 177.750 ;
        RECT 57.465 177.735 58.385 177.740 ;
        RECT 57.465 177.720 58.375 177.735 ;
        RECT 57.465 177.705 58.370 177.720 ;
        RECT 57.465 177.680 58.360 177.705 ;
        RECT 57.465 177.610 58.355 177.680 ;
        RECT 54.565 176.715 55.455 176.885 ;
        RECT 55.625 176.505 56.835 177.255 ;
        RECT 57.005 176.505 57.295 177.230 ;
        RECT 57.465 177.055 58.015 177.440 ;
        RECT 58.185 176.885 58.355 177.610 ;
        RECT 57.465 176.715 58.355 176.885 ;
        RECT 58.525 177.210 58.855 177.635 ;
        RECT 59.025 177.410 59.255 177.805 ;
        RECT 58.525 176.725 58.745 177.210 ;
        RECT 59.425 177.155 59.595 178.185 ;
        RECT 59.765 177.965 61.435 179.055 ;
        RECT 62.125 177.995 62.455 178.840 ;
        RECT 62.625 178.045 62.795 179.055 ;
        RECT 62.965 178.325 63.305 178.885 ;
        RECT 63.535 178.555 63.850 179.055 ;
        RECT 64.030 178.585 64.915 178.755 ;
        RECT 58.915 176.505 59.165 177.045 ;
        RECT 59.335 176.675 59.595 177.155 ;
        RECT 59.765 177.275 60.515 177.795 ;
        RECT 60.685 177.445 61.435 177.965 ;
        RECT 62.065 177.915 62.455 177.995 ;
        RECT 62.965 177.950 63.860 178.325 ;
        RECT 62.065 177.865 62.280 177.915 ;
        RECT 62.065 177.285 62.235 177.865 ;
        RECT 62.965 177.745 63.155 177.950 ;
        RECT 64.030 177.745 64.200 178.585 ;
        RECT 65.140 178.555 65.390 178.885 ;
        RECT 62.405 177.415 63.155 177.745 ;
        RECT 63.325 177.415 64.200 177.745 ;
        RECT 59.765 176.505 61.435 177.275 ;
        RECT 62.065 177.245 62.290 177.285 ;
        RECT 62.955 177.245 63.155 177.415 ;
        RECT 62.065 177.160 62.445 177.245 ;
        RECT 62.115 176.725 62.445 177.160 ;
        RECT 62.615 176.505 62.785 177.115 ;
        RECT 62.955 176.720 63.285 177.245 ;
        RECT 63.545 176.505 63.755 177.035 ;
        RECT 64.030 176.955 64.200 177.415 ;
        RECT 64.370 177.455 64.690 178.415 ;
        RECT 64.860 177.665 65.050 178.385 ;
        RECT 65.220 177.485 65.390 178.555 ;
        RECT 65.560 178.255 65.730 179.055 ;
        RECT 65.900 178.610 67.005 178.780 ;
        RECT 65.900 177.995 66.070 178.610 ;
        RECT 67.215 178.460 67.465 178.885 ;
        RECT 67.635 178.595 67.900 179.055 ;
        RECT 66.240 178.075 66.770 178.440 ;
        RECT 67.215 178.330 67.520 178.460 ;
        RECT 65.560 177.905 66.070 177.995 ;
        RECT 65.560 177.735 66.430 177.905 ;
        RECT 65.560 177.665 65.730 177.735 ;
        RECT 65.850 177.485 66.050 177.515 ;
        RECT 64.370 177.125 64.835 177.455 ;
        RECT 65.220 177.185 66.050 177.485 ;
        RECT 65.220 176.955 65.390 177.185 ;
        RECT 64.030 176.785 64.815 176.955 ;
        RECT 64.985 176.785 65.390 176.955 ;
        RECT 65.570 176.505 65.940 177.005 ;
        RECT 66.260 176.955 66.430 177.735 ;
        RECT 66.600 177.375 66.770 178.075 ;
        RECT 66.940 177.545 67.180 178.140 ;
        RECT 66.600 177.155 67.125 177.375 ;
        RECT 67.350 177.225 67.520 178.330 ;
        RECT 67.295 177.095 67.520 177.225 ;
        RECT 67.690 177.135 67.970 178.085 ;
        RECT 67.295 176.955 67.465 177.095 ;
        RECT 66.260 176.785 66.935 176.955 ;
        RECT 67.130 176.785 67.465 176.955 ;
        RECT 67.635 176.505 67.885 176.965 ;
        RECT 68.140 176.765 68.325 178.885 ;
        RECT 68.495 178.555 68.825 179.055 ;
        RECT 68.995 178.385 69.165 178.885 ;
        RECT 68.500 178.215 69.165 178.385 ;
        RECT 68.500 177.225 68.730 178.215 ;
        RECT 68.900 177.395 69.250 178.045 ;
        RECT 69.425 177.915 69.705 179.055 ;
        RECT 69.875 177.905 70.205 178.885 ;
        RECT 70.375 177.915 70.635 179.055 ;
        RECT 71.355 178.125 71.525 178.885 ;
        RECT 71.740 178.295 72.070 179.055 ;
        RECT 71.355 177.955 72.070 178.125 ;
        RECT 72.240 177.980 72.495 178.885 ;
        RECT 69.435 177.475 69.770 177.745 ;
        RECT 69.940 177.305 70.110 177.905 ;
        RECT 70.280 177.495 70.615 177.745 ;
        RECT 71.265 177.405 71.620 177.775 ;
        RECT 71.900 177.745 72.070 177.955 ;
        RECT 71.900 177.415 72.155 177.745 ;
        RECT 68.500 177.055 69.165 177.225 ;
        RECT 68.495 176.505 68.825 176.885 ;
        RECT 68.995 176.765 69.165 177.055 ;
        RECT 69.425 176.505 69.735 177.305 ;
        RECT 69.940 176.675 70.635 177.305 ;
        RECT 71.900 177.225 72.070 177.415 ;
        RECT 72.325 177.250 72.495 177.980 ;
        RECT 72.670 177.905 72.930 179.055 ;
        RECT 73.105 177.965 76.615 179.055 ;
        RECT 71.355 177.055 72.070 177.225 ;
        RECT 71.355 176.675 71.525 177.055 ;
        RECT 71.740 176.505 72.070 176.885 ;
        RECT 72.240 176.675 72.495 177.250 ;
        RECT 72.670 176.505 72.930 177.345 ;
        RECT 73.105 177.275 74.755 177.795 ;
        RECT 74.925 177.445 76.615 177.965 ;
        RECT 77.795 178.045 77.965 178.885 ;
        RECT 78.135 178.715 79.305 178.885 ;
        RECT 78.135 178.215 78.465 178.715 ;
        RECT 78.975 178.675 79.305 178.715 ;
        RECT 79.495 178.635 79.850 179.055 ;
        RECT 78.635 178.455 78.865 178.545 ;
        RECT 80.020 178.455 80.270 178.885 ;
        RECT 78.635 178.215 80.270 178.455 ;
        RECT 80.440 178.295 80.770 179.055 ;
        RECT 80.940 178.215 81.195 178.885 ;
        RECT 80.985 178.205 81.195 178.215 ;
        RECT 77.795 177.875 80.855 178.045 ;
        RECT 77.710 177.495 78.060 177.705 ;
        RECT 78.230 177.495 78.675 177.695 ;
        RECT 78.845 177.495 79.320 177.695 ;
        RECT 73.105 176.505 76.615 177.275 ;
        RECT 77.795 177.155 78.860 177.325 ;
        RECT 77.795 176.675 77.965 177.155 ;
        RECT 78.135 176.505 78.465 176.985 ;
        RECT 78.690 176.925 78.860 177.155 ;
        RECT 79.040 177.095 79.320 177.495 ;
        RECT 79.590 177.495 79.920 177.695 ;
        RECT 80.090 177.495 80.455 177.695 ;
        RECT 79.590 177.095 79.875 177.495 ;
        RECT 80.685 177.325 80.855 177.875 ;
        RECT 80.055 177.155 80.855 177.325 ;
        RECT 80.055 176.925 80.225 177.155 ;
        RECT 81.025 177.085 81.195 178.205 ;
        RECT 81.395 177.915 81.725 179.055 ;
        RECT 82.255 178.085 82.585 178.870 ;
        RECT 81.905 177.915 82.585 178.085 ;
        RECT 81.385 177.495 81.735 177.745 ;
        RECT 81.905 177.315 82.075 177.915 ;
        RECT 82.765 177.890 83.055 179.055 ;
        RECT 83.225 177.915 83.565 178.885 ;
        RECT 83.735 177.915 83.905 179.055 ;
        RECT 84.175 178.255 84.425 179.055 ;
        RECT 85.070 178.085 85.400 178.885 ;
        RECT 85.700 178.255 86.030 179.055 ;
        RECT 86.200 178.085 86.530 178.885 ;
        RECT 84.095 177.915 86.530 178.085 ;
        RECT 86.905 177.965 90.415 179.055 ;
        RECT 82.245 177.495 82.595 177.745 ;
        RECT 81.010 177.005 81.195 177.085 ;
        RECT 78.690 176.675 80.225 176.925 ;
        RECT 80.395 176.505 80.725 176.985 ;
        RECT 80.940 176.675 81.195 177.005 ;
        RECT 81.395 176.505 81.665 177.315 ;
        RECT 81.835 176.675 82.165 177.315 ;
        RECT 82.335 176.505 82.575 177.315 ;
        RECT 83.225 177.305 83.400 177.915 ;
        RECT 84.095 177.665 84.265 177.915 ;
        RECT 83.570 177.495 84.265 177.665 ;
        RECT 84.440 177.495 84.860 177.695 ;
        RECT 85.030 177.495 85.360 177.695 ;
        RECT 85.530 177.495 85.860 177.695 ;
        RECT 82.765 176.505 83.055 177.230 ;
        RECT 83.225 176.675 83.565 177.305 ;
        RECT 83.735 176.505 83.985 177.305 ;
        RECT 84.175 177.155 85.400 177.325 ;
        RECT 84.175 176.675 84.505 177.155 ;
        RECT 84.675 176.505 84.900 176.965 ;
        RECT 85.070 176.675 85.400 177.155 ;
        RECT 86.030 177.285 86.200 177.915 ;
        RECT 86.385 177.495 86.735 177.745 ;
        RECT 86.030 176.675 86.530 177.285 ;
        RECT 86.905 177.275 88.555 177.795 ;
        RECT 88.725 177.445 90.415 177.965 ;
        RECT 91.045 177.965 92.255 179.055 ;
        RECT 91.045 177.425 91.565 177.965 ;
        RECT 86.905 176.505 90.415 177.275 ;
        RECT 91.735 177.255 92.255 177.795 ;
        RECT 91.045 176.505 92.255 177.255 ;
        RECT 18.280 176.335 92.340 176.505 ;
        RECT 18.365 175.585 19.575 176.335 ;
        RECT 19.745 175.790 25.090 176.335 ;
        RECT 25.265 175.790 30.610 176.335 ;
        RECT 18.365 175.045 18.885 175.585 ;
        RECT 19.055 174.875 19.575 175.415 ;
        RECT 21.330 174.960 21.670 175.790 ;
        RECT 18.365 173.785 19.575 174.875 ;
        RECT 23.150 174.220 23.500 175.470 ;
        RECT 26.850 174.960 27.190 175.790 ;
        RECT 30.785 175.565 34.295 176.335 ;
        RECT 34.515 175.680 34.845 176.115 ;
        RECT 35.015 175.725 35.185 176.335 ;
        RECT 34.465 175.595 34.845 175.680 ;
        RECT 35.355 175.595 35.685 176.120 ;
        RECT 35.945 175.805 36.155 176.335 ;
        RECT 36.430 175.885 37.215 176.055 ;
        RECT 37.385 175.885 37.790 176.055 ;
        RECT 28.670 174.220 29.020 175.470 ;
        RECT 30.785 175.045 32.435 175.565 ;
        RECT 34.465 175.555 34.690 175.595 ;
        RECT 32.605 174.875 34.295 175.395 ;
        RECT 19.745 173.785 25.090 174.220 ;
        RECT 25.265 173.785 30.610 174.220 ;
        RECT 30.785 173.785 34.295 174.875 ;
        RECT 34.465 174.975 34.635 175.555 ;
        RECT 35.355 175.425 35.555 175.595 ;
        RECT 36.430 175.425 36.600 175.885 ;
        RECT 34.805 175.095 35.555 175.425 ;
        RECT 35.725 175.095 36.600 175.425 ;
        RECT 34.465 174.925 34.680 174.975 ;
        RECT 34.465 174.845 34.855 174.925 ;
        RECT 34.525 174.000 34.855 174.845 ;
        RECT 35.365 174.890 35.555 175.095 ;
        RECT 35.025 173.785 35.195 174.795 ;
        RECT 35.365 174.515 36.260 174.890 ;
        RECT 35.365 173.955 35.705 174.515 ;
        RECT 35.935 173.785 36.250 174.285 ;
        RECT 36.430 174.255 36.600 175.095 ;
        RECT 36.770 175.385 37.235 175.715 ;
        RECT 37.620 175.655 37.790 175.885 ;
        RECT 37.970 175.835 38.340 176.335 ;
        RECT 38.660 175.885 39.335 176.055 ;
        RECT 39.530 175.885 39.865 176.055 ;
        RECT 36.770 174.425 37.090 175.385 ;
        RECT 37.620 175.355 38.450 175.655 ;
        RECT 37.260 174.455 37.450 175.175 ;
        RECT 37.620 174.285 37.790 175.355 ;
        RECT 38.250 175.325 38.450 175.355 ;
        RECT 37.960 175.105 38.130 175.175 ;
        RECT 38.660 175.105 38.830 175.885 ;
        RECT 39.695 175.745 39.865 175.885 ;
        RECT 40.035 175.875 40.285 176.335 ;
        RECT 37.960 174.935 38.830 175.105 ;
        RECT 39.000 175.465 39.525 175.685 ;
        RECT 39.695 175.615 39.920 175.745 ;
        RECT 37.960 174.845 38.470 174.935 ;
        RECT 36.430 174.085 37.315 174.255 ;
        RECT 37.540 173.955 37.790 174.285 ;
        RECT 37.960 173.785 38.130 174.585 ;
        RECT 38.300 174.230 38.470 174.845 ;
        RECT 39.000 174.765 39.170 175.465 ;
        RECT 38.640 174.400 39.170 174.765 ;
        RECT 39.340 174.700 39.580 175.295 ;
        RECT 39.750 174.510 39.920 175.615 ;
        RECT 40.090 174.755 40.370 175.705 ;
        RECT 39.615 174.380 39.920 174.510 ;
        RECT 38.300 174.060 39.405 174.230 ;
        RECT 39.615 173.955 39.865 174.380 ;
        RECT 40.035 173.785 40.300 174.245 ;
        RECT 40.540 173.955 40.725 176.075 ;
        RECT 40.895 175.955 41.225 176.335 ;
        RECT 41.395 175.785 41.565 176.075 ;
        RECT 40.900 175.615 41.565 175.785 ;
        RECT 40.900 174.625 41.130 175.615 ;
        RECT 41.835 175.525 42.105 176.335 ;
        RECT 42.275 175.525 42.605 176.165 ;
        RECT 42.775 175.525 43.015 176.335 ;
        RECT 44.125 175.610 44.415 176.335 ;
        RECT 45.505 175.595 46.015 176.165 ;
        RECT 46.185 175.775 46.355 176.335 ;
        RECT 46.560 175.765 46.890 176.165 ;
        RECT 47.065 175.935 47.395 176.335 ;
        RECT 47.630 175.955 49.015 176.165 ;
        RECT 47.630 175.765 47.960 175.955 ;
        RECT 46.560 175.595 47.960 175.765 ;
        RECT 48.130 175.595 48.555 175.785 ;
        RECT 48.725 175.685 49.015 175.955 ;
        RECT 41.300 174.795 41.650 175.445 ;
        RECT 41.825 175.095 42.175 175.345 ;
        RECT 42.345 174.925 42.515 175.525 ;
        RECT 42.685 175.095 43.035 175.345 ;
        RECT 45.505 174.975 45.680 175.595 ;
        RECT 45.865 175.345 46.055 175.425 ;
        RECT 46.425 175.345 46.595 175.425 ;
        RECT 45.865 175.095 46.230 175.345 ;
        RECT 46.425 175.095 46.675 175.345 ;
        RECT 46.885 175.095 47.230 175.425 ;
        RECT 40.900 174.455 41.565 174.625 ;
        RECT 40.895 173.785 41.225 174.285 ;
        RECT 41.395 173.955 41.565 174.455 ;
        RECT 41.835 173.785 42.165 174.925 ;
        RECT 42.345 174.755 43.025 174.925 ;
        RECT 42.695 173.970 43.025 174.755 ;
        RECT 44.125 173.785 44.415 174.950 ;
        RECT 45.505 174.925 45.735 174.975 ;
        RECT 46.060 174.925 46.230 175.095 ;
        RECT 45.505 173.965 45.890 174.925 ;
        RECT 46.060 174.755 46.735 174.925 ;
        RECT 46.105 173.785 46.395 174.585 ;
        RECT 46.565 174.125 46.735 174.755 ;
        RECT 46.905 174.295 47.230 175.095 ;
        RECT 47.400 174.760 47.675 175.425 ;
        RECT 47.860 174.760 48.215 175.425 ;
        RECT 48.385 174.585 48.555 175.595 ;
        RECT 49.225 175.515 49.455 176.335 ;
        RECT 49.625 175.535 49.955 176.165 ;
        RECT 48.740 175.095 49.015 175.425 ;
        RECT 49.205 175.095 49.535 175.345 ;
        RECT 49.705 174.935 49.955 175.535 ;
        RECT 50.125 175.515 50.335 176.335 ;
        RECT 51.050 175.945 51.380 176.335 ;
        RECT 51.550 175.775 51.775 176.155 ;
        RECT 51.035 175.095 51.275 175.745 ;
        RECT 51.445 175.595 51.775 175.775 ;
        RECT 47.600 174.335 48.555 174.585 ;
        RECT 47.600 174.125 47.930 174.335 ;
        RECT 46.565 173.955 47.930 174.125 ;
        RECT 48.725 173.785 49.015 174.925 ;
        RECT 49.225 173.785 49.455 174.925 ;
        RECT 49.625 173.955 49.955 174.935 ;
        RECT 51.445 174.925 51.620 175.595 ;
        RECT 51.975 175.425 52.205 176.045 ;
        RECT 52.385 175.605 52.685 176.335 ;
        RECT 53.365 175.515 53.595 176.335 ;
        RECT 53.765 175.535 54.095 176.165 ;
        RECT 51.790 175.095 52.205 175.425 ;
        RECT 52.385 175.095 52.680 175.425 ;
        RECT 53.345 175.095 53.675 175.345 ;
        RECT 53.845 174.935 54.095 175.535 ;
        RECT 54.265 175.515 54.475 176.335 ;
        RECT 54.705 175.565 57.295 176.335 ;
        RECT 58.015 175.855 58.315 176.335 ;
        RECT 58.485 175.685 58.745 176.140 ;
        RECT 58.915 175.855 59.175 176.335 ;
        RECT 59.355 175.685 59.615 176.140 ;
        RECT 59.785 175.855 60.035 176.335 ;
        RECT 60.215 175.685 60.475 176.140 ;
        RECT 60.645 175.855 60.895 176.335 ;
        RECT 61.075 175.685 61.335 176.140 ;
        RECT 61.505 175.855 61.750 176.335 ;
        RECT 61.920 175.685 62.195 176.140 ;
        RECT 62.365 175.855 62.610 176.335 ;
        RECT 62.780 175.685 63.040 176.140 ;
        RECT 63.210 175.855 63.470 176.335 ;
        RECT 63.640 175.685 63.900 176.140 ;
        RECT 64.070 175.855 64.330 176.335 ;
        RECT 64.500 175.685 64.760 176.140 ;
        RECT 64.930 175.775 65.190 176.335 ;
        RECT 54.705 175.045 55.915 175.565 ;
        RECT 58.015 175.515 64.760 175.685 ;
        RECT 50.125 173.785 50.335 174.925 ;
        RECT 51.035 174.735 51.620 174.925 ;
        RECT 51.035 173.965 51.310 174.735 ;
        RECT 51.790 174.565 52.685 174.895 ;
        RECT 51.480 174.395 52.685 174.565 ;
        RECT 51.480 173.965 51.810 174.395 ;
        RECT 51.980 173.785 52.175 174.225 ;
        RECT 52.355 173.965 52.685 174.395 ;
        RECT 53.365 173.785 53.595 174.925 ;
        RECT 53.765 173.955 54.095 174.935 ;
        RECT 54.265 173.785 54.475 174.925 ;
        RECT 56.085 174.875 57.295 175.395 ;
        RECT 54.705 173.785 57.295 174.875 ;
        RECT 58.015 174.925 59.180 175.515 ;
        RECT 65.360 175.345 65.610 176.155 ;
        RECT 65.790 175.810 66.050 176.335 ;
        RECT 66.220 175.345 66.470 176.155 ;
        RECT 66.650 175.825 66.955 176.335 ;
        RECT 59.350 175.095 66.470 175.345 ;
        RECT 66.640 175.095 66.955 175.655 ;
        RECT 67.125 175.565 69.715 176.335 ;
        RECT 69.885 175.610 70.175 176.335 ;
        RECT 70.675 175.935 71.005 176.335 ;
        RECT 71.175 175.765 71.505 176.105 ;
        RECT 72.555 175.935 72.885 176.335 ;
        RECT 70.520 175.595 72.885 175.765 ;
        RECT 73.055 175.610 73.385 176.120 ;
        RECT 58.015 174.700 64.760 174.925 ;
        RECT 58.015 173.785 58.285 174.530 ;
        RECT 58.455 173.960 58.745 174.700 ;
        RECT 59.355 174.685 64.760 174.700 ;
        RECT 58.915 173.790 59.170 174.515 ;
        RECT 59.355 173.960 59.615 174.685 ;
        RECT 59.785 173.790 60.030 174.515 ;
        RECT 60.215 173.960 60.475 174.685 ;
        RECT 60.645 173.790 60.890 174.515 ;
        RECT 61.075 173.960 61.335 174.685 ;
        RECT 61.505 173.790 61.750 174.515 ;
        RECT 61.920 173.960 62.180 174.685 ;
        RECT 62.350 173.790 62.610 174.515 ;
        RECT 62.780 173.960 63.040 174.685 ;
        RECT 63.210 173.790 63.470 174.515 ;
        RECT 63.640 173.960 63.900 174.685 ;
        RECT 64.070 173.790 64.330 174.515 ;
        RECT 64.500 173.960 64.760 174.685 ;
        RECT 64.930 173.790 65.190 174.585 ;
        RECT 65.360 173.960 65.610 175.095 ;
        RECT 58.915 173.785 65.190 173.790 ;
        RECT 65.790 173.785 66.050 174.595 ;
        RECT 66.225 173.955 66.470 175.095 ;
        RECT 67.125 175.045 68.335 175.565 ;
        RECT 68.505 174.875 69.715 175.395 ;
        RECT 66.650 173.785 66.945 174.595 ;
        RECT 67.125 173.785 69.715 174.875 ;
        RECT 69.885 173.785 70.175 174.950 ;
        RECT 70.520 174.595 70.690 175.595 ;
        RECT 72.715 175.425 72.885 175.595 ;
        RECT 70.860 174.765 71.105 175.425 ;
        RECT 71.320 174.765 71.585 175.425 ;
        RECT 71.780 174.765 72.065 175.425 ;
        RECT 72.240 175.095 72.545 175.425 ;
        RECT 72.715 175.095 73.025 175.425 ;
        RECT 72.240 174.765 72.455 175.095 ;
        RECT 70.520 174.425 70.975 174.595 ;
        RECT 70.645 173.995 70.975 174.425 ;
        RECT 71.155 174.425 72.445 174.595 ;
        RECT 71.155 174.005 71.405 174.425 ;
        RECT 71.635 173.785 71.965 174.255 ;
        RECT 72.195 174.005 72.445 174.425 ;
        RECT 72.635 173.785 72.885 174.925 ;
        RECT 73.195 174.845 73.385 175.610 ;
        RECT 73.055 173.995 73.385 174.845 ;
        RECT 73.570 175.660 73.845 176.005 ;
        RECT 74.035 175.935 74.415 176.335 ;
        RECT 74.585 175.765 74.755 176.115 ;
        RECT 74.925 175.935 75.255 176.335 ;
        RECT 75.425 175.765 75.680 176.115 ;
        RECT 73.570 174.925 73.740 175.660 ;
        RECT 74.015 175.595 75.680 175.765 ;
        RECT 74.015 175.425 74.185 175.595 ;
        RECT 75.865 175.585 77.075 176.335 ;
        RECT 77.410 175.825 77.650 176.335 ;
        RECT 77.830 175.825 78.110 176.155 ;
        RECT 78.340 175.825 78.555 176.335 ;
        RECT 73.910 175.095 74.185 175.425 ;
        RECT 74.355 175.095 75.180 175.425 ;
        RECT 75.350 175.095 75.695 175.425 ;
        RECT 74.015 174.925 74.185 175.095 ;
        RECT 73.570 173.955 73.845 174.925 ;
        RECT 74.015 174.755 74.675 174.925 ;
        RECT 74.985 174.805 75.180 175.095 ;
        RECT 75.865 175.045 76.385 175.585 ;
        RECT 74.505 174.635 74.675 174.755 ;
        RECT 75.350 174.635 75.675 174.925 ;
        RECT 76.555 174.875 77.075 175.415 ;
        RECT 77.305 175.095 77.660 175.655 ;
        RECT 77.830 174.925 78.000 175.825 ;
        RECT 78.170 175.095 78.435 175.655 ;
        RECT 78.725 175.595 79.340 176.165 ;
        RECT 78.685 174.925 78.855 175.425 ;
        RECT 74.055 173.785 74.335 174.585 ;
        RECT 74.505 174.465 75.675 174.635 ;
        RECT 74.505 174.005 75.695 174.295 ;
        RECT 75.865 173.785 77.075 174.875 ;
        RECT 77.430 174.755 78.855 174.925 ;
        RECT 77.430 174.580 77.820 174.755 ;
        RECT 78.305 173.785 78.635 174.585 ;
        RECT 79.025 174.575 79.340 175.595 ;
        RECT 79.545 175.565 82.135 176.335 ;
        RECT 82.395 175.785 82.565 176.075 ;
        RECT 82.735 175.955 83.065 176.335 ;
        RECT 82.395 175.615 83.060 175.785 ;
        RECT 79.545 175.045 80.755 175.565 ;
        RECT 80.925 174.875 82.135 175.395 ;
        RECT 78.805 173.955 79.340 174.575 ;
        RECT 79.545 173.785 82.135 174.875 ;
        RECT 82.310 174.795 82.660 175.445 ;
        RECT 82.830 174.625 83.060 175.615 ;
        RECT 82.395 174.455 83.060 174.625 ;
        RECT 82.395 173.955 82.565 174.455 ;
        RECT 82.735 173.785 83.065 174.285 ;
        RECT 83.235 173.955 83.460 176.075 ;
        RECT 83.675 175.875 83.925 176.335 ;
        RECT 84.110 175.885 84.440 176.055 ;
        RECT 84.620 175.885 85.370 176.055 ;
        RECT 83.660 174.755 83.940 175.355 ;
        RECT 84.110 174.355 84.280 175.885 ;
        RECT 84.450 175.385 85.030 175.715 ;
        RECT 84.450 174.515 84.690 175.385 ;
        RECT 85.200 175.105 85.370 175.885 ;
        RECT 85.620 175.835 85.990 176.335 ;
        RECT 86.170 175.885 86.630 176.055 ;
        RECT 86.860 175.885 87.530 176.055 ;
        RECT 86.170 175.655 86.340 175.885 ;
        RECT 85.540 175.355 86.340 175.655 ;
        RECT 86.510 175.385 87.060 175.715 ;
        RECT 85.540 175.325 85.710 175.355 ;
        RECT 85.830 175.105 86.000 175.175 ;
        RECT 85.200 174.935 86.000 175.105 ;
        RECT 85.490 174.845 86.000 174.935 ;
        RECT 84.880 174.410 85.320 174.765 ;
        RECT 83.660 173.785 83.925 174.245 ;
        RECT 84.110 173.980 84.345 174.355 ;
        RECT 85.490 174.230 85.660 174.845 ;
        RECT 84.590 174.060 85.660 174.230 ;
        RECT 85.830 173.785 86.000 174.585 ;
        RECT 86.170 174.285 86.340 175.355 ;
        RECT 86.510 174.455 86.700 175.175 ;
        RECT 86.870 174.845 87.060 175.385 ;
        RECT 87.360 175.345 87.530 175.885 ;
        RECT 87.845 175.805 88.015 176.335 ;
        RECT 88.310 175.685 88.670 176.125 ;
        RECT 88.845 175.855 89.015 176.335 ;
        RECT 89.205 175.690 89.540 176.115 ;
        RECT 89.715 175.860 89.885 176.335 ;
        RECT 90.060 175.690 90.395 176.115 ;
        RECT 90.565 175.860 90.735 176.335 ;
        RECT 88.310 175.515 88.810 175.685 ;
        RECT 89.205 175.520 90.875 175.690 ;
        RECT 91.045 175.585 92.255 176.335 ;
        RECT 88.640 175.345 88.810 175.515 ;
        RECT 87.360 175.175 88.450 175.345 ;
        RECT 88.640 175.175 90.460 175.345 ;
        RECT 86.870 174.515 87.190 174.845 ;
        RECT 86.170 173.955 86.420 174.285 ;
        RECT 87.360 174.255 87.530 175.175 ;
        RECT 88.640 174.920 88.810 175.175 ;
        RECT 90.630 174.955 90.875 175.520 ;
        RECT 87.700 174.750 88.810 174.920 ;
        RECT 89.205 174.785 90.875 174.955 ;
        RECT 91.045 174.875 91.565 175.415 ;
        RECT 91.735 175.045 92.255 175.585 ;
        RECT 87.700 174.590 88.560 174.750 ;
        RECT 86.645 174.085 87.530 174.255 ;
        RECT 87.710 173.785 87.925 174.285 ;
        RECT 88.390 173.965 88.560 174.590 ;
        RECT 88.845 173.785 89.025 174.565 ;
        RECT 89.205 174.025 89.540 174.785 ;
        RECT 89.720 173.785 89.890 174.615 ;
        RECT 90.060 174.025 90.390 174.785 ;
        RECT 90.560 173.785 90.730 174.615 ;
        RECT 91.045 173.785 92.255 174.875 ;
        RECT 18.280 173.615 92.340 173.785 ;
        RECT 18.365 172.525 19.575 173.615 ;
        RECT 19.745 173.180 25.090 173.615 ;
        RECT 25.265 173.180 30.610 173.615 ;
        RECT 18.365 171.815 18.885 172.355 ;
        RECT 19.055 171.985 19.575 172.525 ;
        RECT 18.365 171.065 19.575 171.815 ;
        RECT 21.330 171.610 21.670 172.440 ;
        RECT 23.150 171.930 23.500 173.180 ;
        RECT 26.850 171.610 27.190 172.440 ;
        RECT 28.670 171.930 29.020 173.180 ;
        RECT 31.245 172.450 31.535 173.615 ;
        RECT 31.705 173.180 37.050 173.615 ;
        RECT 19.745 171.065 25.090 171.610 ;
        RECT 25.265 171.065 30.610 171.610 ;
        RECT 31.245 171.065 31.535 171.790 ;
        RECT 33.290 171.610 33.630 172.440 ;
        RECT 35.110 171.930 35.460 173.180 ;
        RECT 38.260 172.985 38.545 173.445 ;
        RECT 38.715 173.155 38.985 173.615 ;
        RECT 38.260 172.765 39.215 172.985 ;
        RECT 38.145 172.035 38.835 172.595 ;
        RECT 39.005 171.865 39.215 172.765 ;
        RECT 38.260 171.695 39.215 171.865 ;
        RECT 39.385 172.595 39.785 173.445 ;
        RECT 39.975 172.985 40.255 173.445 ;
        RECT 40.775 173.155 41.100 173.615 ;
        RECT 39.975 172.765 41.100 172.985 ;
        RECT 39.385 172.035 40.480 172.595 ;
        RECT 40.650 172.305 41.100 172.765 ;
        RECT 41.270 172.475 41.655 173.445 ;
        RECT 41.825 172.525 44.415 173.615 ;
        RECT 31.705 171.065 37.050 171.610 ;
        RECT 38.260 171.235 38.545 171.695 ;
        RECT 38.715 171.065 38.985 171.525 ;
        RECT 39.385 171.235 39.785 172.035 ;
        RECT 40.650 171.975 41.205 172.305 ;
        RECT 40.650 171.865 41.100 171.975 ;
        RECT 39.975 171.695 41.100 171.865 ;
        RECT 41.375 171.805 41.655 172.475 ;
        RECT 39.975 171.235 40.255 171.695 ;
        RECT 40.775 171.065 41.100 171.525 ;
        RECT 41.270 171.235 41.655 171.805 ;
        RECT 41.825 171.835 43.035 172.355 ;
        RECT 43.205 172.005 44.415 172.525 ;
        RECT 45.055 173.005 45.385 173.435 ;
        RECT 45.565 173.175 45.760 173.615 ;
        RECT 45.930 173.005 46.260 173.435 ;
        RECT 45.055 172.835 46.260 173.005 ;
        RECT 45.055 172.505 45.950 172.835 ;
        RECT 46.430 172.665 46.705 173.435 ;
        RECT 46.120 172.475 46.705 172.665 ;
        RECT 46.885 172.525 50.395 173.615 ;
        RECT 45.060 171.975 45.355 172.305 ;
        RECT 45.535 171.975 45.950 172.305 ;
        RECT 41.825 171.065 44.415 171.835 ;
        RECT 45.055 171.065 45.355 171.795 ;
        RECT 45.535 171.355 45.765 171.975 ;
        RECT 46.120 171.805 46.295 172.475 ;
        RECT 45.965 171.625 46.295 171.805 ;
        RECT 46.465 171.655 46.705 172.305 ;
        RECT 46.885 171.835 48.535 172.355 ;
        RECT 48.705 172.005 50.395 172.525 ;
        RECT 51.025 172.475 51.305 173.615 ;
        RECT 51.475 172.465 51.805 173.445 ;
        RECT 51.975 172.475 52.235 173.615 ;
        RECT 52.605 172.945 52.885 173.615 ;
        RECT 53.055 172.725 53.355 173.275 ;
        RECT 53.555 172.895 53.885 173.615 ;
        RECT 54.075 172.895 54.535 173.445 ;
        RECT 51.035 172.035 51.370 172.305 ;
        RECT 51.540 171.865 51.710 172.465 ;
        RECT 52.420 172.305 52.685 172.665 ;
        RECT 53.055 172.555 53.995 172.725 ;
        RECT 53.825 172.305 53.995 172.555 ;
        RECT 51.880 172.055 52.215 172.305 ;
        RECT 52.420 172.055 53.095 172.305 ;
        RECT 53.315 172.055 53.655 172.305 ;
        RECT 53.825 171.975 54.115 172.305 ;
        RECT 53.825 171.885 53.995 171.975 ;
        RECT 45.965 171.245 46.190 171.625 ;
        RECT 46.360 171.065 46.690 171.455 ;
        RECT 46.885 171.065 50.395 171.835 ;
        RECT 51.025 171.065 51.335 171.865 ;
        RECT 51.540 171.235 52.235 171.865 ;
        RECT 52.605 171.695 53.995 171.885 ;
        RECT 52.605 171.335 52.935 171.695 ;
        RECT 54.285 171.525 54.535 172.895 ;
        RECT 54.890 172.645 55.280 172.820 ;
        RECT 55.765 172.815 56.095 173.615 ;
        RECT 56.265 172.825 56.800 173.445 ;
        RECT 54.890 172.475 56.315 172.645 ;
        RECT 54.765 171.745 55.120 172.305 ;
        RECT 55.290 171.575 55.460 172.475 ;
        RECT 55.630 171.745 55.895 172.305 ;
        RECT 56.145 171.975 56.315 172.475 ;
        RECT 56.485 171.805 56.800 172.825 ;
        RECT 57.005 172.450 57.295 173.615 ;
        RECT 57.555 173.275 58.715 173.445 ;
        RECT 57.555 172.775 57.725 173.275 ;
        RECT 57.985 172.645 58.155 173.105 ;
        RECT 58.385 173.025 58.715 173.275 ;
        RECT 58.940 173.195 59.270 173.615 ;
        RECT 59.525 173.025 59.810 173.445 ;
        RECT 58.385 172.855 59.810 173.025 ;
        RECT 60.055 172.815 60.385 173.615 ;
        RECT 60.635 172.895 60.970 173.405 ;
        RECT 57.530 172.305 57.735 172.595 ;
        RECT 57.985 172.475 60.355 172.645 ;
        RECT 60.185 172.305 60.355 172.475 ;
        RECT 57.530 172.255 57.880 172.305 ;
        RECT 57.525 172.085 57.880 172.255 ;
        RECT 57.530 171.975 57.880 172.085 ;
        RECT 53.555 171.065 53.805 171.525 ;
        RECT 53.975 171.235 54.535 171.525 ;
        RECT 54.870 171.065 55.110 171.575 ;
        RECT 55.290 171.245 55.570 171.575 ;
        RECT 55.800 171.065 56.015 171.575 ;
        RECT 56.185 171.235 56.800 171.805 ;
        RECT 57.005 171.065 57.295 171.790 ;
        RECT 57.475 171.065 57.805 171.785 ;
        RECT 58.190 171.640 58.610 172.305 ;
        RECT 58.780 171.915 59.070 172.305 ;
        RECT 59.260 171.915 59.530 172.305 ;
        RECT 59.740 172.255 59.990 172.305 ;
        RECT 59.740 172.085 59.995 172.255 ;
        RECT 59.740 171.975 59.990 172.085 ;
        RECT 60.185 171.975 60.490 172.305 ;
        RECT 58.780 171.745 59.075 171.915 ;
        RECT 59.260 171.745 59.535 171.915 ;
        RECT 60.185 171.805 60.355 171.975 ;
        RECT 58.780 171.645 59.070 171.745 ;
        RECT 59.260 171.645 59.530 171.745 ;
        RECT 59.795 171.635 60.355 171.805 ;
        RECT 59.795 171.465 59.965 171.635 ;
        RECT 60.715 171.540 60.970 172.895 ;
        RECT 61.145 172.475 61.425 173.615 ;
        RECT 61.595 172.465 61.925 173.445 ;
        RECT 62.095 172.475 62.355 173.615 ;
        RECT 62.585 172.555 62.915 173.400 ;
        RECT 63.085 172.605 63.255 173.615 ;
        RECT 63.425 172.885 63.765 173.445 ;
        RECT 63.995 173.115 64.310 173.615 ;
        RECT 64.490 173.145 65.375 173.315 ;
        RECT 62.525 172.475 62.915 172.555 ;
        RECT 63.425 172.510 64.320 172.885 ;
        RECT 61.155 172.035 61.490 172.305 ;
        RECT 61.660 171.915 61.830 172.465 ;
        RECT 62.525 172.425 62.740 172.475 ;
        RECT 62.000 172.055 62.335 172.305 ;
        RECT 61.660 171.865 61.835 171.915 ;
        RECT 58.350 171.295 59.965 171.465 ;
        RECT 60.135 171.065 60.465 171.465 ;
        RECT 60.635 171.280 60.970 171.540 ;
        RECT 61.145 171.065 61.455 171.865 ;
        RECT 61.660 171.235 62.355 171.865 ;
        RECT 62.525 171.845 62.695 172.425 ;
        RECT 63.425 172.305 63.615 172.510 ;
        RECT 64.490 172.305 64.660 173.145 ;
        RECT 65.600 173.115 65.850 173.445 ;
        RECT 62.865 171.975 63.615 172.305 ;
        RECT 63.785 171.975 64.660 172.305 ;
        RECT 62.525 171.805 62.750 171.845 ;
        RECT 63.415 171.805 63.615 171.975 ;
        RECT 62.525 171.720 62.905 171.805 ;
        RECT 62.575 171.285 62.905 171.720 ;
        RECT 63.075 171.065 63.245 171.675 ;
        RECT 63.415 171.280 63.745 171.805 ;
        RECT 64.005 171.065 64.215 171.595 ;
        RECT 64.490 171.515 64.660 171.975 ;
        RECT 64.830 172.015 65.150 172.975 ;
        RECT 65.320 172.225 65.510 172.945 ;
        RECT 65.680 172.045 65.850 173.115 ;
        RECT 66.020 172.815 66.190 173.615 ;
        RECT 66.360 173.170 67.465 173.340 ;
        RECT 66.360 172.555 66.530 173.170 ;
        RECT 67.675 173.020 67.925 173.445 ;
        RECT 68.095 173.155 68.360 173.615 ;
        RECT 66.700 172.635 67.230 173.000 ;
        RECT 67.675 172.890 67.980 173.020 ;
        RECT 66.020 172.465 66.530 172.555 ;
        RECT 66.020 172.295 66.890 172.465 ;
        RECT 66.020 172.225 66.190 172.295 ;
        RECT 66.310 172.045 66.510 172.075 ;
        RECT 64.830 171.685 65.295 172.015 ;
        RECT 65.680 171.745 66.510 172.045 ;
        RECT 65.680 171.515 65.850 171.745 ;
        RECT 64.490 171.345 65.275 171.515 ;
        RECT 65.445 171.345 65.850 171.515 ;
        RECT 66.030 171.065 66.400 171.565 ;
        RECT 66.720 171.515 66.890 172.295 ;
        RECT 67.060 171.935 67.230 172.635 ;
        RECT 67.400 172.105 67.640 172.700 ;
        RECT 67.060 171.715 67.585 171.935 ;
        RECT 67.810 171.785 67.980 172.890 ;
        RECT 67.755 171.655 67.980 171.785 ;
        RECT 68.150 171.695 68.430 172.645 ;
        RECT 67.755 171.515 67.925 171.655 ;
        RECT 66.720 171.345 67.395 171.515 ;
        RECT 67.590 171.345 67.925 171.515 ;
        RECT 68.095 171.065 68.345 171.525 ;
        RECT 68.600 171.325 68.785 173.445 ;
        RECT 68.955 173.115 69.285 173.615 ;
        RECT 69.455 172.945 69.625 173.445 ;
        RECT 68.960 172.775 69.625 172.945 ;
        RECT 68.960 171.785 69.190 172.775 ;
        RECT 69.360 171.955 69.710 172.605 ;
        RECT 69.885 172.525 72.475 173.615 ;
        RECT 69.885 171.835 71.095 172.355 ;
        RECT 71.265 172.005 72.475 172.525 ;
        RECT 73.115 173.005 73.445 173.435 ;
        RECT 73.625 173.175 73.820 173.615 ;
        RECT 73.990 173.005 74.320 173.435 ;
        RECT 73.115 172.835 74.320 173.005 ;
        RECT 73.115 172.505 74.010 172.835 ;
        RECT 74.490 172.665 74.765 173.435 ;
        RECT 74.180 172.475 74.765 172.665 ;
        RECT 75.405 172.745 75.680 173.445 ;
        RECT 75.850 173.070 76.105 173.615 ;
        RECT 76.275 173.105 76.755 173.445 ;
        RECT 76.930 173.060 77.535 173.615 ;
        RECT 76.920 172.960 77.535 173.060 ;
        RECT 76.920 172.935 77.105 172.960 ;
        RECT 73.120 171.975 73.415 172.305 ;
        RECT 73.595 171.975 74.010 172.305 ;
        RECT 68.960 171.615 69.625 171.785 ;
        RECT 68.955 171.065 69.285 171.445 ;
        RECT 69.455 171.325 69.625 171.615 ;
        RECT 69.885 171.065 72.475 171.835 ;
        RECT 73.115 171.065 73.415 171.795 ;
        RECT 73.595 171.355 73.825 171.975 ;
        RECT 74.180 171.805 74.355 172.475 ;
        RECT 74.025 171.625 74.355 171.805 ;
        RECT 74.525 171.655 74.765 172.305 ;
        RECT 75.405 171.715 75.575 172.745 ;
        RECT 75.850 172.615 76.605 172.865 ;
        RECT 76.775 172.690 77.105 172.935 ;
        RECT 75.850 172.580 76.620 172.615 ;
        RECT 75.850 172.570 76.635 172.580 ;
        RECT 75.745 172.555 76.640 172.570 ;
        RECT 75.745 172.540 76.660 172.555 ;
        RECT 75.745 172.530 76.680 172.540 ;
        RECT 75.745 172.520 76.705 172.530 ;
        RECT 75.745 172.490 76.775 172.520 ;
        RECT 75.745 172.460 76.795 172.490 ;
        RECT 75.745 172.430 76.815 172.460 ;
        RECT 75.745 172.405 76.845 172.430 ;
        RECT 75.745 172.370 76.880 172.405 ;
        RECT 75.745 172.365 76.910 172.370 ;
        RECT 75.745 171.970 75.975 172.365 ;
        RECT 76.520 172.360 76.910 172.365 ;
        RECT 76.545 172.350 76.910 172.360 ;
        RECT 76.560 172.345 76.910 172.350 ;
        RECT 76.575 172.340 76.910 172.345 ;
        RECT 77.275 172.340 77.535 172.790 ;
        RECT 77.705 172.525 78.915 173.615 ;
        RECT 79.090 173.235 79.425 173.615 ;
        RECT 76.575 172.335 77.535 172.340 ;
        RECT 76.585 172.325 77.535 172.335 ;
        RECT 76.595 172.320 77.535 172.325 ;
        RECT 76.605 172.310 77.535 172.320 ;
        RECT 76.610 172.300 77.535 172.310 ;
        RECT 76.615 172.295 77.535 172.300 ;
        RECT 76.625 172.280 77.535 172.295 ;
        RECT 76.630 172.265 77.535 172.280 ;
        RECT 76.640 172.240 77.535 172.265 ;
        RECT 76.145 171.770 76.475 172.195 ;
        RECT 74.025 171.245 74.250 171.625 ;
        RECT 74.420 171.065 74.750 171.455 ;
        RECT 75.405 171.235 75.665 171.715 ;
        RECT 75.835 171.065 76.085 171.605 ;
        RECT 76.255 171.285 76.475 171.770 ;
        RECT 76.645 172.170 77.535 172.240 ;
        RECT 76.645 171.445 76.815 172.170 ;
        RECT 76.985 171.615 77.535 172.000 ;
        RECT 77.705 171.815 78.225 172.355 ;
        RECT 78.395 171.985 78.915 172.525 ;
        RECT 76.645 171.275 77.535 171.445 ;
        RECT 77.705 171.065 78.915 171.815 ;
        RECT 79.085 171.745 79.325 173.055 ;
        RECT 79.595 172.645 79.845 173.445 ;
        RECT 80.065 172.895 80.395 173.615 ;
        RECT 80.580 172.645 80.830 173.445 ;
        RECT 81.295 172.815 81.625 173.615 ;
        RECT 81.795 173.185 82.135 173.445 ;
        RECT 79.495 172.475 81.685 172.645 ;
        RECT 79.495 171.565 79.665 172.475 ;
        RECT 81.370 172.305 81.685 172.475 ;
        RECT 79.170 171.235 79.665 171.565 ;
        RECT 79.885 171.340 80.235 172.305 ;
        RECT 80.415 171.335 80.715 172.305 ;
        RECT 80.895 171.335 81.175 172.305 ;
        RECT 81.370 172.055 81.700 172.305 ;
        RECT 81.355 171.065 81.625 171.865 ;
        RECT 81.875 171.785 82.135 173.185 ;
        RECT 82.765 172.450 83.055 173.615 ;
        RECT 83.225 172.460 83.565 173.445 ;
        RECT 83.735 173.185 84.145 173.615 ;
        RECT 84.890 173.195 85.220 173.615 ;
        RECT 85.390 173.015 85.715 173.445 ;
        RECT 83.735 172.845 85.715 173.015 ;
        RECT 83.225 171.805 83.480 172.460 ;
        RECT 83.735 172.305 84.000 172.845 ;
        RECT 84.215 172.505 84.840 172.675 ;
        RECT 83.650 171.975 84.000 172.305 ;
        RECT 84.170 171.975 84.500 172.305 ;
        RECT 84.670 171.805 84.840 172.505 ;
        RECT 81.795 171.275 82.135 171.785 ;
        RECT 82.765 171.065 83.055 171.790 ;
        RECT 83.225 171.430 83.585 171.805 ;
        RECT 83.285 171.405 83.455 171.430 ;
        RECT 83.850 171.065 84.020 171.805 ;
        RECT 84.300 171.635 84.840 171.805 ;
        RECT 85.010 172.435 85.715 172.845 ;
        RECT 86.190 172.515 86.520 173.615 ;
        RECT 87.365 172.475 87.750 173.445 ;
        RECT 87.920 173.155 88.245 173.615 ;
        RECT 88.765 172.985 89.045 173.445 ;
        RECT 87.920 172.765 89.045 172.985 ;
        RECT 84.300 171.430 84.470 171.635 ;
        RECT 85.010 171.235 85.180 172.435 ;
        RECT 85.350 172.055 85.920 172.265 ;
        RECT 86.090 172.055 86.735 172.265 ;
        RECT 85.410 171.715 86.580 171.885 ;
        RECT 85.410 171.235 85.740 171.715 ;
        RECT 85.910 171.065 86.080 171.535 ;
        RECT 86.250 171.250 86.580 171.715 ;
        RECT 87.365 171.805 87.645 172.475 ;
        RECT 87.920 172.305 88.370 172.765 ;
        RECT 89.235 172.595 89.635 173.445 ;
        RECT 90.035 173.155 90.305 173.615 ;
        RECT 90.475 172.985 90.760 173.445 ;
        RECT 87.815 171.975 88.370 172.305 ;
        RECT 88.540 172.035 89.635 172.595 ;
        RECT 87.920 171.865 88.370 171.975 ;
        RECT 87.365 171.235 87.750 171.805 ;
        RECT 87.920 171.695 89.045 171.865 ;
        RECT 87.920 171.065 88.245 171.525 ;
        RECT 88.765 171.235 89.045 171.695 ;
        RECT 89.235 171.235 89.635 172.035 ;
        RECT 89.805 172.765 90.760 172.985 ;
        RECT 89.805 171.865 90.015 172.765 ;
        RECT 90.185 172.035 90.875 172.595 ;
        RECT 91.045 172.525 92.255 173.615 ;
        RECT 91.045 171.985 91.565 172.525 ;
        RECT 89.805 171.695 90.760 171.865 ;
        RECT 91.735 171.815 92.255 172.355 ;
        RECT 90.035 171.065 90.305 171.525 ;
        RECT 90.475 171.235 90.760 171.695 ;
        RECT 91.045 171.065 92.255 171.815 ;
        RECT 18.280 170.895 92.340 171.065 ;
        RECT 18.365 170.145 19.575 170.895 ;
        RECT 19.745 170.350 25.090 170.895 ;
        RECT 25.265 170.350 30.610 170.895 ;
        RECT 18.365 169.605 18.885 170.145 ;
        RECT 19.055 169.435 19.575 169.975 ;
        RECT 21.330 169.520 21.670 170.350 ;
        RECT 18.365 168.345 19.575 169.435 ;
        RECT 23.150 168.780 23.500 170.030 ;
        RECT 26.850 169.520 27.190 170.350 ;
        RECT 30.785 170.125 32.455 170.895 ;
        RECT 33.135 170.240 33.465 170.675 ;
        RECT 33.635 170.285 33.805 170.895 ;
        RECT 33.085 170.155 33.465 170.240 ;
        RECT 33.975 170.155 34.305 170.680 ;
        RECT 34.565 170.365 34.775 170.895 ;
        RECT 35.050 170.445 35.835 170.615 ;
        RECT 36.005 170.445 36.410 170.615 ;
        RECT 28.670 168.780 29.020 170.030 ;
        RECT 30.785 169.605 31.535 170.125 ;
        RECT 33.085 170.115 33.310 170.155 ;
        RECT 31.705 169.435 32.455 169.955 ;
        RECT 19.745 168.345 25.090 168.780 ;
        RECT 25.265 168.345 30.610 168.780 ;
        RECT 30.785 168.345 32.455 169.435 ;
        RECT 33.085 169.535 33.255 170.115 ;
        RECT 33.975 169.985 34.175 170.155 ;
        RECT 35.050 169.985 35.220 170.445 ;
        RECT 33.425 169.655 34.175 169.985 ;
        RECT 34.345 169.655 35.220 169.985 ;
        RECT 33.085 169.485 33.300 169.535 ;
        RECT 33.085 169.405 33.475 169.485 ;
        RECT 33.145 168.560 33.475 169.405 ;
        RECT 33.985 169.450 34.175 169.655 ;
        RECT 33.645 168.345 33.815 169.355 ;
        RECT 33.985 169.075 34.880 169.450 ;
        RECT 33.985 168.515 34.325 169.075 ;
        RECT 34.555 168.345 34.870 168.845 ;
        RECT 35.050 168.815 35.220 169.655 ;
        RECT 35.390 169.945 35.855 170.275 ;
        RECT 36.240 170.215 36.410 170.445 ;
        RECT 36.590 170.395 36.960 170.895 ;
        RECT 37.280 170.445 37.955 170.615 ;
        RECT 38.150 170.445 38.485 170.615 ;
        RECT 35.390 168.985 35.710 169.945 ;
        RECT 36.240 169.915 37.070 170.215 ;
        RECT 35.880 169.015 36.070 169.735 ;
        RECT 36.240 168.845 36.410 169.915 ;
        RECT 36.870 169.885 37.070 169.915 ;
        RECT 36.580 169.665 36.750 169.735 ;
        RECT 37.280 169.665 37.450 170.445 ;
        RECT 38.315 170.305 38.485 170.445 ;
        RECT 38.655 170.435 38.905 170.895 ;
        RECT 36.580 169.495 37.450 169.665 ;
        RECT 37.620 170.025 38.145 170.245 ;
        RECT 38.315 170.175 38.540 170.305 ;
        RECT 36.580 169.405 37.090 169.495 ;
        RECT 35.050 168.645 35.935 168.815 ;
        RECT 36.160 168.515 36.410 168.845 ;
        RECT 36.580 168.345 36.750 169.145 ;
        RECT 36.920 168.790 37.090 169.405 ;
        RECT 37.620 169.325 37.790 170.025 ;
        RECT 37.260 168.960 37.790 169.325 ;
        RECT 37.960 169.260 38.200 169.855 ;
        RECT 38.370 169.070 38.540 170.175 ;
        RECT 38.710 169.315 38.990 170.265 ;
        RECT 38.235 168.940 38.540 169.070 ;
        RECT 36.920 168.620 38.025 168.790 ;
        RECT 38.235 168.515 38.485 168.940 ;
        RECT 38.655 168.345 38.920 168.805 ;
        RECT 39.160 168.515 39.345 170.635 ;
        RECT 39.515 170.515 39.845 170.895 ;
        RECT 40.015 170.345 40.185 170.635 ;
        RECT 40.470 170.505 40.800 170.895 ;
        RECT 39.520 170.175 40.185 170.345 ;
        RECT 40.970 170.335 41.195 170.715 ;
        RECT 39.520 169.185 39.750 170.175 ;
        RECT 39.920 169.355 40.270 170.005 ;
        RECT 40.455 169.655 40.695 170.305 ;
        RECT 40.865 170.155 41.195 170.335 ;
        RECT 40.865 169.485 41.040 170.155 ;
        RECT 41.395 169.985 41.625 170.605 ;
        RECT 41.805 170.165 42.105 170.895 ;
        RECT 42.285 170.095 42.595 170.895 ;
        RECT 42.800 170.095 43.495 170.725 ;
        RECT 44.125 170.170 44.415 170.895 ;
        RECT 42.800 170.045 42.975 170.095 ;
        RECT 41.210 169.655 41.625 169.985 ;
        RECT 41.805 169.655 42.100 169.985 ;
        RECT 42.295 169.655 42.630 169.925 ;
        RECT 42.800 169.495 42.970 170.045 ;
        RECT 43.140 169.655 43.475 169.905 ;
        RECT 40.455 169.295 41.040 169.485 ;
        RECT 39.520 169.015 40.185 169.185 ;
        RECT 39.515 168.345 39.845 168.845 ;
        RECT 40.015 168.515 40.185 169.015 ;
        RECT 40.455 168.525 40.730 169.295 ;
        RECT 41.210 169.125 42.105 169.455 ;
        RECT 40.900 168.955 42.105 169.125 ;
        RECT 40.900 168.525 41.230 168.955 ;
        RECT 41.400 168.345 41.595 168.785 ;
        RECT 41.775 168.525 42.105 168.955 ;
        RECT 42.285 168.345 42.565 169.485 ;
        RECT 42.735 168.515 43.065 169.495 ;
        RECT 43.235 168.345 43.495 169.485 ;
        RECT 44.125 168.345 44.415 169.510 ;
        RECT 44.590 169.295 44.925 170.715 ;
        RECT 45.105 170.525 45.850 170.895 ;
        RECT 46.415 170.355 46.670 170.715 ;
        RECT 46.850 170.525 47.180 170.895 ;
        RECT 47.360 170.355 47.585 170.715 ;
        RECT 45.100 170.165 47.585 170.355 ;
        RECT 45.100 169.475 45.325 170.165 ;
        RECT 47.825 170.085 48.065 170.895 ;
        RECT 48.235 170.085 48.565 170.725 ;
        RECT 48.735 170.085 49.005 170.895 ;
        RECT 49.270 170.395 49.765 170.725 ;
        RECT 45.525 169.655 45.805 169.985 ;
        RECT 45.985 169.655 46.560 169.985 ;
        RECT 46.740 169.655 47.175 169.985 ;
        RECT 47.355 169.655 47.625 169.985 ;
        RECT 47.805 169.655 48.155 169.905 ;
        RECT 48.325 169.485 48.495 170.085 ;
        RECT 48.665 169.655 49.015 169.905 ;
        RECT 45.100 169.295 47.595 169.475 ;
        RECT 44.590 168.525 44.855 169.295 ;
        RECT 45.025 168.345 45.355 169.065 ;
        RECT 45.545 168.885 46.735 169.115 ;
        RECT 45.545 168.525 45.805 168.885 ;
        RECT 45.975 168.345 46.305 168.715 ;
        RECT 46.475 168.525 46.735 168.885 ;
        RECT 47.305 168.525 47.595 169.295 ;
        RECT 47.815 169.315 48.495 169.485 ;
        RECT 47.815 168.530 48.145 169.315 ;
        RECT 48.675 168.345 49.005 169.485 ;
        RECT 49.185 168.905 49.425 170.215 ;
        RECT 49.595 169.485 49.765 170.395 ;
        RECT 49.985 169.655 50.335 170.620 ;
        RECT 50.515 169.655 50.815 170.625 ;
        RECT 50.995 169.655 51.275 170.625 ;
        RECT 51.455 170.095 51.725 170.895 ;
        RECT 51.895 170.175 52.235 170.685 ;
        RECT 52.405 170.350 57.750 170.895 ;
        RECT 51.470 169.655 51.800 169.905 ;
        RECT 51.470 169.485 51.785 169.655 ;
        RECT 49.595 169.315 51.785 169.485 ;
        RECT 49.190 168.345 49.525 168.725 ;
        RECT 49.695 168.515 49.945 169.315 ;
        RECT 50.165 168.345 50.495 169.065 ;
        RECT 50.680 168.515 50.930 169.315 ;
        RECT 51.395 168.345 51.725 169.145 ;
        RECT 51.975 168.775 52.235 170.175 ;
        RECT 53.990 169.520 54.330 170.350 ;
        RECT 57.925 170.125 60.515 170.895 ;
        RECT 60.885 170.265 61.215 170.625 ;
        RECT 61.835 170.435 62.085 170.895 ;
        RECT 62.255 170.435 62.815 170.725 ;
        RECT 55.810 168.780 56.160 170.030 ;
        RECT 57.925 169.605 59.135 170.125 ;
        RECT 60.885 170.075 62.275 170.265 ;
        RECT 62.105 169.985 62.275 170.075 ;
        RECT 59.305 169.435 60.515 169.955 ;
        RECT 51.895 168.515 52.235 168.775 ;
        RECT 52.405 168.345 57.750 168.780 ;
        RECT 57.925 168.345 60.515 169.435 ;
        RECT 60.700 169.655 61.375 169.905 ;
        RECT 61.595 169.655 61.935 169.905 ;
        RECT 62.105 169.655 62.395 169.985 ;
        RECT 60.700 169.295 60.965 169.655 ;
        RECT 62.105 169.405 62.275 169.655 ;
        RECT 61.335 169.235 62.275 169.405 ;
        RECT 60.885 168.345 61.165 169.015 ;
        RECT 61.335 168.685 61.635 169.235 ;
        RECT 62.565 169.065 62.815 170.435 ;
        RECT 63.075 170.345 63.245 170.725 ;
        RECT 63.425 170.515 63.755 170.895 ;
        RECT 63.075 170.175 63.740 170.345 ;
        RECT 63.935 170.220 64.195 170.725 ;
        RECT 64.365 170.350 69.710 170.895 ;
        RECT 63.005 169.625 63.335 169.995 ;
        RECT 63.570 169.920 63.740 170.175 ;
        RECT 63.570 169.590 63.855 169.920 ;
        RECT 63.570 169.445 63.740 169.590 ;
        RECT 61.835 168.345 62.165 169.065 ;
        RECT 62.355 168.515 62.815 169.065 ;
        RECT 63.075 169.275 63.740 169.445 ;
        RECT 64.025 169.420 64.195 170.220 ;
        RECT 65.950 169.520 66.290 170.350 ;
        RECT 69.885 170.170 70.175 170.895 ;
        RECT 70.345 170.125 72.015 170.895 ;
        RECT 72.650 170.130 73.105 170.895 ;
        RECT 73.380 170.515 74.680 170.725 ;
        RECT 74.935 170.535 75.265 170.895 ;
        RECT 74.510 170.365 74.680 170.515 ;
        RECT 75.435 170.395 75.695 170.725 ;
        RECT 63.075 168.515 63.245 169.275 ;
        RECT 63.425 168.345 63.755 169.105 ;
        RECT 63.925 168.515 64.195 169.420 ;
        RECT 67.770 168.780 68.120 170.030 ;
        RECT 70.345 169.605 71.095 170.125 ;
        RECT 64.365 168.345 69.710 168.780 ;
        RECT 69.885 168.345 70.175 169.510 ;
        RECT 71.265 169.435 72.015 169.955 ;
        RECT 73.580 169.905 73.800 170.305 ;
        RECT 72.645 169.705 73.135 169.905 ;
        RECT 73.325 169.695 73.800 169.905 ;
        RECT 74.045 169.905 74.255 170.305 ;
        RECT 74.510 170.240 75.265 170.365 ;
        RECT 74.510 170.195 75.355 170.240 ;
        RECT 75.085 170.075 75.355 170.195 ;
        RECT 74.045 169.695 74.375 169.905 ;
        RECT 74.545 169.635 74.955 169.940 ;
        RECT 70.345 168.345 72.015 169.435 ;
        RECT 72.650 169.465 73.825 169.525 ;
        RECT 75.185 169.500 75.355 170.075 ;
        RECT 75.155 169.465 75.355 169.500 ;
        RECT 72.650 169.355 75.355 169.465 ;
        RECT 72.650 168.735 72.905 169.355 ;
        RECT 73.495 169.295 75.295 169.355 ;
        RECT 73.495 169.265 73.825 169.295 ;
        RECT 75.525 169.195 75.695 170.395 ;
        RECT 75.885 170.085 76.125 170.895 ;
        RECT 76.295 170.085 76.625 170.725 ;
        RECT 76.795 170.085 77.065 170.895 ;
        RECT 77.245 170.125 80.755 170.895 ;
        RECT 80.925 170.145 82.135 170.895 ;
        RECT 82.395 170.345 82.565 170.635 ;
        RECT 82.735 170.515 83.065 170.895 ;
        RECT 82.395 170.175 83.060 170.345 ;
        RECT 75.865 169.655 76.215 169.905 ;
        RECT 76.385 169.485 76.555 170.085 ;
        RECT 76.725 169.655 77.075 169.905 ;
        RECT 77.245 169.605 78.895 170.125 ;
        RECT 73.155 169.095 73.340 169.185 ;
        RECT 73.930 169.095 74.765 169.105 ;
        RECT 73.155 168.895 74.765 169.095 ;
        RECT 73.155 168.855 73.385 168.895 ;
        RECT 72.650 168.515 72.985 168.735 ;
        RECT 73.990 168.345 74.345 168.725 ;
        RECT 74.515 168.515 74.765 168.895 ;
        RECT 75.015 168.345 75.265 169.125 ;
        RECT 75.435 168.515 75.695 169.195 ;
        RECT 75.875 169.315 76.555 169.485 ;
        RECT 75.875 168.530 76.205 169.315 ;
        RECT 76.735 168.345 77.065 169.485 ;
        RECT 79.065 169.435 80.755 169.955 ;
        RECT 80.925 169.605 81.445 170.145 ;
        RECT 81.615 169.435 82.135 169.975 ;
        RECT 77.245 168.345 80.755 169.435 ;
        RECT 80.925 168.345 82.135 169.435 ;
        RECT 82.310 169.355 82.660 170.005 ;
        RECT 82.830 169.185 83.060 170.175 ;
        RECT 82.395 169.015 83.060 169.185 ;
        RECT 82.395 168.515 82.565 169.015 ;
        RECT 82.735 168.345 83.065 168.845 ;
        RECT 83.235 168.515 83.460 170.635 ;
        RECT 83.675 170.435 83.925 170.895 ;
        RECT 84.110 170.445 84.440 170.615 ;
        RECT 84.620 170.445 85.370 170.615 ;
        RECT 83.660 169.315 83.940 169.915 ;
        RECT 84.110 168.915 84.280 170.445 ;
        RECT 84.450 169.945 85.030 170.275 ;
        RECT 84.450 169.075 84.690 169.945 ;
        RECT 85.200 169.665 85.370 170.445 ;
        RECT 85.620 170.395 85.990 170.895 ;
        RECT 86.170 170.445 86.630 170.615 ;
        RECT 86.860 170.445 87.530 170.615 ;
        RECT 86.170 170.215 86.340 170.445 ;
        RECT 85.540 169.915 86.340 170.215 ;
        RECT 86.510 169.945 87.060 170.275 ;
        RECT 85.540 169.885 85.710 169.915 ;
        RECT 85.830 169.665 86.000 169.735 ;
        RECT 85.200 169.495 86.000 169.665 ;
        RECT 85.490 169.405 86.000 169.495 ;
        RECT 84.880 168.970 85.320 169.325 ;
        RECT 83.660 168.345 83.925 168.805 ;
        RECT 84.110 168.540 84.345 168.915 ;
        RECT 85.490 168.790 85.660 169.405 ;
        RECT 84.590 168.620 85.660 168.790 ;
        RECT 85.830 168.345 86.000 169.145 ;
        RECT 86.170 168.845 86.340 169.915 ;
        RECT 86.510 169.015 86.700 169.735 ;
        RECT 86.870 169.405 87.060 169.945 ;
        RECT 87.360 169.905 87.530 170.445 ;
        RECT 87.845 170.365 88.015 170.895 ;
        RECT 88.310 170.245 88.670 170.685 ;
        RECT 88.845 170.415 89.015 170.895 ;
        RECT 89.205 170.250 89.540 170.675 ;
        RECT 89.715 170.420 89.885 170.895 ;
        RECT 90.060 170.250 90.395 170.675 ;
        RECT 90.565 170.420 90.735 170.895 ;
        RECT 88.310 170.075 88.810 170.245 ;
        RECT 89.205 170.080 90.875 170.250 ;
        RECT 91.045 170.145 92.255 170.895 ;
        RECT 88.640 169.905 88.810 170.075 ;
        RECT 87.360 169.735 88.450 169.905 ;
        RECT 88.640 169.735 90.460 169.905 ;
        RECT 86.870 169.075 87.190 169.405 ;
        RECT 86.170 168.515 86.420 168.845 ;
        RECT 87.360 168.815 87.530 169.735 ;
        RECT 88.640 169.480 88.810 169.735 ;
        RECT 90.630 169.515 90.875 170.080 ;
        RECT 87.700 169.310 88.810 169.480 ;
        RECT 89.205 169.345 90.875 169.515 ;
        RECT 91.045 169.435 91.565 169.975 ;
        RECT 91.735 169.605 92.255 170.145 ;
        RECT 87.700 169.150 88.560 169.310 ;
        RECT 86.645 168.645 87.530 168.815 ;
        RECT 87.710 168.345 87.925 168.845 ;
        RECT 88.390 168.525 88.560 169.150 ;
        RECT 88.845 168.345 89.025 169.125 ;
        RECT 89.205 168.585 89.540 169.345 ;
        RECT 89.720 168.345 89.890 169.175 ;
        RECT 90.060 168.585 90.390 169.345 ;
        RECT 90.560 168.345 90.730 169.175 ;
        RECT 91.045 168.345 92.255 169.435 ;
        RECT 18.280 168.175 92.340 168.345 ;
        RECT 18.365 167.085 19.575 168.175 ;
        RECT 19.745 167.740 25.090 168.175 ;
        RECT 25.265 167.740 30.610 168.175 ;
        RECT 18.365 166.375 18.885 166.915 ;
        RECT 19.055 166.545 19.575 167.085 ;
        RECT 18.365 165.625 19.575 166.375 ;
        RECT 21.330 166.170 21.670 167.000 ;
        RECT 23.150 166.490 23.500 167.740 ;
        RECT 26.850 166.170 27.190 167.000 ;
        RECT 28.670 166.490 29.020 167.740 ;
        RECT 31.245 167.010 31.535 168.175 ;
        RECT 31.705 167.740 37.050 168.175 ;
        RECT 37.225 167.740 42.570 168.175 ;
        RECT 42.745 167.740 48.090 168.175 ;
        RECT 19.745 165.625 25.090 166.170 ;
        RECT 25.265 165.625 30.610 166.170 ;
        RECT 31.245 165.625 31.535 166.350 ;
        RECT 33.290 166.170 33.630 167.000 ;
        RECT 35.110 166.490 35.460 167.740 ;
        RECT 38.810 166.170 39.150 167.000 ;
        RECT 40.630 166.490 40.980 167.740 ;
        RECT 44.330 166.170 44.670 167.000 ;
        RECT 46.150 166.490 46.500 167.740 ;
        RECT 48.265 167.085 51.775 168.175 ;
        RECT 51.945 167.085 53.155 168.175 ;
        RECT 53.525 167.505 53.805 168.175 ;
        RECT 53.975 167.285 54.275 167.835 ;
        RECT 54.475 167.455 54.805 168.175 ;
        RECT 54.995 167.455 55.455 168.005 ;
        RECT 48.265 166.395 49.915 166.915 ;
        RECT 50.085 166.565 51.775 167.085 ;
        RECT 31.705 165.625 37.050 166.170 ;
        RECT 37.225 165.625 42.570 166.170 ;
        RECT 42.745 165.625 48.090 166.170 ;
        RECT 48.265 165.625 51.775 166.395 ;
        RECT 51.945 166.375 52.465 166.915 ;
        RECT 52.635 166.545 53.155 167.085 ;
        RECT 53.340 166.865 53.605 167.225 ;
        RECT 53.975 167.115 54.915 167.285 ;
        RECT 54.745 166.865 54.915 167.115 ;
        RECT 53.340 166.615 54.015 166.865 ;
        RECT 54.235 166.615 54.575 166.865 ;
        RECT 54.745 166.535 55.035 166.865 ;
        RECT 54.745 166.445 54.915 166.535 ;
        RECT 51.945 165.625 53.155 166.375 ;
        RECT 53.525 166.255 54.915 166.445 ;
        RECT 53.525 165.895 53.855 166.255 ;
        RECT 55.205 166.085 55.455 167.455 ;
        RECT 55.625 167.085 56.835 168.175 ;
        RECT 54.475 165.625 54.725 166.085 ;
        RECT 54.895 165.795 55.455 166.085 ;
        RECT 55.625 166.375 56.145 166.915 ;
        RECT 56.315 166.545 56.835 167.085 ;
        RECT 57.005 167.010 57.295 168.175 ;
        RECT 57.470 167.455 57.805 167.965 ;
        RECT 55.625 165.625 56.835 166.375 ;
        RECT 57.005 165.625 57.295 166.350 ;
        RECT 57.470 166.100 57.725 167.455 ;
        RECT 58.055 167.375 58.385 168.175 ;
        RECT 58.630 167.585 58.915 168.005 ;
        RECT 59.170 167.755 59.500 168.175 ;
        RECT 59.725 167.835 60.885 168.005 ;
        RECT 59.725 167.585 60.055 167.835 ;
        RECT 58.630 167.415 60.055 167.585 ;
        RECT 60.285 167.205 60.455 167.665 ;
        RECT 60.715 167.335 60.885 167.835 ;
        RECT 58.085 167.035 60.455 167.205 ;
        RECT 61.145 167.205 61.455 168.005 ;
        RECT 61.625 167.375 61.935 168.175 ;
        RECT 62.105 167.545 62.365 168.005 ;
        RECT 62.535 167.715 62.790 168.175 ;
        RECT 62.965 167.545 63.225 168.005 ;
        RECT 62.105 167.375 63.225 167.545 ;
        RECT 58.085 166.865 58.255 167.035 ;
        RECT 60.705 166.985 60.915 167.155 ;
        RECT 61.145 167.035 62.175 167.205 ;
        RECT 60.705 166.865 60.910 166.985 ;
        RECT 57.950 166.535 58.255 166.865 ;
        RECT 58.450 166.815 58.700 166.865 ;
        RECT 58.445 166.645 58.700 166.815 ;
        RECT 58.450 166.535 58.700 166.645 ;
        RECT 58.085 166.365 58.255 166.535 ;
        RECT 58.910 166.475 59.180 166.865 ;
        RECT 59.370 166.475 59.660 166.865 ;
        RECT 58.085 166.195 58.645 166.365 ;
        RECT 58.905 166.305 59.180 166.475 ;
        RECT 59.365 166.305 59.660 166.475 ;
        RECT 58.910 166.205 59.180 166.305 ;
        RECT 59.370 166.205 59.660 166.305 ;
        RECT 59.830 166.200 60.250 166.865 ;
        RECT 60.560 166.535 60.910 166.865 ;
        RECT 57.470 165.840 57.805 166.100 ;
        RECT 58.475 166.025 58.645 166.195 ;
        RECT 57.975 165.625 58.305 166.025 ;
        RECT 58.475 165.855 60.090 166.025 ;
        RECT 60.635 165.625 60.965 166.345 ;
        RECT 61.145 166.125 61.315 167.035 ;
        RECT 61.485 166.295 61.835 166.865 ;
        RECT 62.005 166.785 62.175 167.035 ;
        RECT 62.965 167.125 63.225 167.375 ;
        RECT 63.395 167.305 63.680 168.175 ;
        RECT 63.905 167.740 69.250 168.175 ;
        RECT 62.965 166.955 63.720 167.125 ;
        RECT 62.005 166.615 63.145 166.785 ;
        RECT 63.315 166.445 63.720 166.955 ;
        RECT 62.070 166.275 63.720 166.445 ;
        RECT 61.145 165.795 61.445 166.125 ;
        RECT 61.615 165.625 61.890 166.105 ;
        RECT 62.070 165.885 62.365 166.275 ;
        RECT 62.535 165.625 62.790 166.105 ;
        RECT 62.965 165.885 63.225 166.275 ;
        RECT 65.490 166.170 65.830 167.000 ;
        RECT 67.310 166.490 67.660 167.740 ;
        RECT 69.425 167.085 72.015 168.175 ;
        RECT 69.425 166.395 70.635 166.915 ;
        RECT 70.805 166.565 72.015 167.085 ;
        RECT 72.185 167.035 72.570 168.005 ;
        RECT 72.740 167.715 73.065 168.175 ;
        RECT 73.585 167.545 73.865 168.005 ;
        RECT 72.740 167.325 73.865 167.545 ;
        RECT 63.395 165.625 63.675 166.105 ;
        RECT 63.905 165.625 69.250 166.170 ;
        RECT 69.425 165.625 72.015 166.395 ;
        RECT 72.185 166.365 72.465 167.035 ;
        RECT 72.740 166.865 73.190 167.325 ;
        RECT 74.055 167.155 74.455 168.005 ;
        RECT 74.855 167.715 75.125 168.175 ;
        RECT 75.295 167.545 75.580 168.005 ;
        RECT 72.635 166.535 73.190 166.865 ;
        RECT 73.360 166.595 74.455 167.155 ;
        RECT 72.740 166.425 73.190 166.535 ;
        RECT 72.185 165.795 72.570 166.365 ;
        RECT 72.740 166.255 73.865 166.425 ;
        RECT 72.740 165.625 73.065 166.085 ;
        RECT 73.585 165.795 73.865 166.255 ;
        RECT 74.055 165.795 74.455 166.595 ;
        RECT 74.625 167.325 75.580 167.545 ;
        RECT 76.335 167.565 76.665 167.995 ;
        RECT 76.845 167.735 77.040 168.175 ;
        RECT 77.210 167.565 77.540 167.995 ;
        RECT 76.335 167.395 77.540 167.565 ;
        RECT 74.625 166.425 74.835 167.325 ;
        RECT 75.005 166.595 75.695 167.155 ;
        RECT 76.335 167.065 77.230 167.395 ;
        RECT 77.710 167.225 77.985 167.995 ;
        RECT 77.400 167.035 77.985 167.225 ;
        RECT 78.175 167.205 78.505 167.990 ;
        RECT 78.175 167.035 78.855 167.205 ;
        RECT 79.035 167.035 79.365 168.175 ;
        RECT 79.545 167.085 82.135 168.175 ;
        RECT 76.340 166.535 76.635 166.865 ;
        RECT 76.815 166.535 77.230 166.865 ;
        RECT 74.625 166.255 75.580 166.425 ;
        RECT 74.855 165.625 75.125 166.085 ;
        RECT 75.295 165.795 75.580 166.255 ;
        RECT 76.335 165.625 76.635 166.355 ;
        RECT 76.815 165.915 77.045 166.535 ;
        RECT 77.400 166.365 77.575 167.035 ;
        RECT 77.245 166.185 77.575 166.365 ;
        RECT 77.745 166.215 77.985 166.865 ;
        RECT 78.165 166.615 78.515 166.865 ;
        RECT 78.685 166.435 78.855 167.035 ;
        RECT 79.025 166.615 79.375 166.865 ;
        RECT 77.245 165.805 77.470 166.185 ;
        RECT 77.640 165.625 77.970 166.015 ;
        RECT 78.185 165.625 78.425 166.435 ;
        RECT 78.595 165.795 78.925 166.435 ;
        RECT 79.095 165.625 79.365 166.435 ;
        RECT 79.545 166.395 80.755 166.915 ;
        RECT 80.925 166.565 82.135 167.085 ;
        RECT 82.765 167.010 83.055 168.175 ;
        RECT 83.225 167.740 88.570 168.175 ;
        RECT 79.545 165.625 82.135 166.395 ;
        RECT 82.765 165.625 83.055 166.350 ;
        RECT 84.810 166.170 85.150 167.000 ;
        RECT 86.630 166.490 86.980 167.740 ;
        RECT 88.745 167.085 90.415 168.175 ;
        RECT 88.745 166.395 89.495 166.915 ;
        RECT 89.665 166.565 90.415 167.085 ;
        RECT 91.045 167.085 92.255 168.175 ;
        RECT 91.045 166.545 91.565 167.085 ;
        RECT 83.225 165.625 88.570 166.170 ;
        RECT 88.745 165.625 90.415 166.395 ;
        RECT 91.735 166.375 92.255 166.915 ;
        RECT 91.045 165.625 92.255 166.375 ;
        RECT 18.280 165.455 92.340 165.625 ;
        RECT 18.365 164.705 19.575 165.455 ;
        RECT 19.745 164.910 25.090 165.455 ;
        RECT 25.265 164.910 30.610 165.455 ;
        RECT 30.785 164.910 36.130 165.455 ;
        RECT 18.365 164.165 18.885 164.705 ;
        RECT 19.055 163.995 19.575 164.535 ;
        RECT 21.330 164.080 21.670 164.910 ;
        RECT 18.365 162.905 19.575 163.995 ;
        RECT 23.150 163.340 23.500 164.590 ;
        RECT 26.850 164.080 27.190 164.910 ;
        RECT 28.670 163.340 29.020 164.590 ;
        RECT 32.370 164.080 32.710 164.910 ;
        RECT 36.305 164.685 37.975 165.455 ;
        RECT 34.190 163.340 34.540 164.590 ;
        RECT 36.305 164.165 37.055 164.685 ;
        RECT 38.625 164.645 38.865 165.455 ;
        RECT 39.035 164.645 39.365 165.285 ;
        RECT 39.535 164.645 39.805 165.455 ;
        RECT 39.985 164.685 43.495 165.455 ;
        RECT 44.125 164.730 44.415 165.455 ;
        RECT 44.585 164.715 45.095 165.285 ;
        RECT 45.265 164.895 45.435 165.455 ;
        RECT 45.640 164.885 45.970 165.285 ;
        RECT 46.145 165.055 46.475 165.455 ;
        RECT 46.710 165.075 48.095 165.285 ;
        RECT 46.710 164.885 47.040 165.075 ;
        RECT 45.640 164.715 47.040 164.885 ;
        RECT 47.210 164.715 47.635 164.905 ;
        RECT 47.805 164.805 48.095 165.075 ;
        RECT 48.265 164.805 48.525 165.285 ;
        RECT 48.695 164.915 48.945 165.455 ;
        RECT 37.225 163.995 37.975 164.515 ;
        RECT 38.605 164.215 38.955 164.465 ;
        RECT 39.125 164.045 39.295 164.645 ;
        RECT 39.465 164.215 39.815 164.465 ;
        RECT 39.985 164.165 41.635 164.685 ;
        RECT 19.745 162.905 25.090 163.340 ;
        RECT 25.265 162.905 30.610 163.340 ;
        RECT 30.785 162.905 36.130 163.340 ;
        RECT 36.305 162.905 37.975 163.995 ;
        RECT 38.615 163.875 39.295 164.045 ;
        RECT 38.615 163.090 38.945 163.875 ;
        RECT 39.475 162.905 39.805 164.045 ;
        RECT 41.805 163.995 43.495 164.515 ;
        RECT 44.585 164.095 44.760 164.715 ;
        RECT 44.945 164.465 45.135 164.545 ;
        RECT 45.505 164.465 45.675 164.545 ;
        RECT 44.945 164.215 45.310 164.465 ;
        RECT 45.505 164.215 45.755 164.465 ;
        RECT 45.965 164.215 46.310 164.545 ;
        RECT 39.985 162.905 43.495 163.995 ;
        RECT 44.125 162.905 44.415 164.070 ;
        RECT 44.585 164.045 44.815 164.095 ;
        RECT 45.140 164.045 45.310 164.215 ;
        RECT 44.585 163.085 44.970 164.045 ;
        RECT 45.140 163.875 45.815 164.045 ;
        RECT 45.185 162.905 45.475 163.705 ;
        RECT 45.645 163.245 45.815 163.875 ;
        RECT 45.985 163.415 46.310 164.215 ;
        RECT 46.480 163.880 46.755 164.545 ;
        RECT 46.940 163.880 47.295 164.545 ;
        RECT 47.465 163.705 47.635 164.715 ;
        RECT 47.820 164.215 48.095 164.545 ;
        RECT 46.680 163.455 47.635 163.705 ;
        RECT 46.680 163.245 47.010 163.455 ;
        RECT 45.645 163.075 47.010 163.245 ;
        RECT 47.805 162.905 48.095 164.045 ;
        RECT 48.265 163.775 48.435 164.805 ;
        RECT 49.115 164.750 49.335 165.235 ;
        RECT 48.605 164.155 48.835 164.550 ;
        RECT 49.005 164.325 49.335 164.750 ;
        RECT 49.505 165.075 50.395 165.245 ;
        RECT 49.505 164.350 49.675 165.075 ;
        RECT 50.565 164.995 51.125 165.285 ;
        RECT 51.295 164.995 51.545 165.455 ;
        RECT 49.845 164.520 50.395 164.905 ;
        RECT 49.505 164.280 50.395 164.350 ;
        RECT 49.500 164.255 50.395 164.280 ;
        RECT 49.490 164.240 50.395 164.255 ;
        RECT 49.485 164.225 50.395 164.240 ;
        RECT 49.475 164.220 50.395 164.225 ;
        RECT 49.470 164.210 50.395 164.220 ;
        RECT 49.465 164.200 50.395 164.210 ;
        RECT 49.455 164.195 50.395 164.200 ;
        RECT 49.445 164.185 50.395 164.195 ;
        RECT 49.435 164.180 50.395 164.185 ;
        RECT 49.435 164.175 49.770 164.180 ;
        RECT 49.420 164.170 49.770 164.175 ;
        RECT 49.405 164.160 49.770 164.170 ;
        RECT 49.380 164.155 49.770 164.160 ;
        RECT 48.605 164.150 49.770 164.155 ;
        RECT 48.605 164.115 49.740 164.150 ;
        RECT 48.605 164.090 49.705 164.115 ;
        RECT 48.605 164.060 49.675 164.090 ;
        RECT 48.605 164.030 49.655 164.060 ;
        RECT 48.605 164.000 49.635 164.030 ;
        RECT 48.605 163.990 49.565 164.000 ;
        RECT 48.605 163.980 49.540 163.990 ;
        RECT 48.605 163.965 49.520 163.980 ;
        RECT 48.605 163.950 49.500 163.965 ;
        RECT 48.710 163.940 49.495 163.950 ;
        RECT 48.710 163.905 49.480 163.940 ;
        RECT 48.265 163.075 48.540 163.775 ;
        RECT 48.710 163.655 49.465 163.905 ;
        RECT 49.635 163.585 49.965 163.830 ;
        RECT 50.135 163.730 50.395 164.180 ;
        RECT 49.780 163.560 49.965 163.585 ;
        RECT 50.565 163.625 50.815 164.995 ;
        RECT 52.165 164.825 52.495 165.185 ;
        RECT 51.105 164.635 52.495 164.825 ;
        RECT 52.865 164.655 53.560 165.285 ;
        RECT 53.765 164.655 54.075 165.455 ;
        RECT 54.410 164.945 54.650 165.455 ;
        RECT 54.830 164.945 55.110 165.275 ;
        RECT 55.340 164.945 55.555 165.455 ;
        RECT 51.105 164.545 51.275 164.635 ;
        RECT 53.385 164.605 53.560 164.655 ;
        RECT 50.985 164.215 51.275 164.545 ;
        RECT 51.445 164.215 51.785 164.465 ;
        RECT 52.005 164.215 52.680 164.465 ;
        RECT 52.885 164.215 53.220 164.465 ;
        RECT 51.105 163.965 51.275 164.215 ;
        RECT 51.105 163.795 52.045 163.965 ;
        RECT 52.415 163.855 52.680 164.215 ;
        RECT 53.390 164.055 53.560 164.605 ;
        RECT 53.730 164.215 54.065 164.485 ;
        RECT 54.305 164.215 54.660 164.775 ;
        RECT 49.780 163.460 50.395 163.560 ;
        RECT 48.710 162.905 48.965 163.450 ;
        RECT 49.135 163.075 49.615 163.415 ;
        RECT 49.790 162.905 50.395 163.460 ;
        RECT 50.565 163.075 51.025 163.625 ;
        RECT 51.215 162.905 51.545 163.625 ;
        RECT 51.745 163.245 52.045 163.795 ;
        RECT 52.215 162.905 52.495 163.575 ;
        RECT 52.865 162.905 53.125 164.045 ;
        RECT 53.295 163.075 53.625 164.055 ;
        RECT 54.830 164.045 55.000 164.945 ;
        RECT 55.170 164.215 55.435 164.775 ;
        RECT 55.725 164.715 56.340 165.285 ;
        RECT 55.685 164.045 55.855 164.545 ;
        RECT 53.795 162.905 54.075 164.045 ;
        RECT 54.430 163.875 55.855 164.045 ;
        RECT 54.430 163.700 54.820 163.875 ;
        RECT 55.305 162.905 55.635 163.705 ;
        RECT 56.025 163.695 56.340 164.715 ;
        RECT 56.745 164.825 57.075 165.185 ;
        RECT 57.695 164.995 57.945 165.455 ;
        RECT 58.115 164.995 58.675 165.285 ;
        RECT 56.745 164.635 58.135 164.825 ;
        RECT 57.965 164.545 58.135 164.635 ;
        RECT 56.560 164.215 57.235 164.465 ;
        RECT 57.455 164.215 57.795 164.465 ;
        RECT 57.965 164.215 58.255 164.545 ;
        RECT 56.560 163.855 56.825 164.215 ;
        RECT 57.965 163.965 58.135 164.215 ;
        RECT 55.805 163.075 56.340 163.695 ;
        RECT 57.195 163.795 58.135 163.965 ;
        RECT 56.745 162.905 57.025 163.575 ;
        RECT 57.195 163.245 57.495 163.795 ;
        RECT 58.425 163.625 58.675 164.995 ;
        RECT 58.895 164.800 59.225 165.235 ;
        RECT 59.395 164.845 59.565 165.455 ;
        RECT 58.845 164.715 59.225 164.800 ;
        RECT 59.735 164.715 60.065 165.240 ;
        RECT 60.325 164.925 60.535 165.455 ;
        RECT 60.810 165.005 61.595 165.175 ;
        RECT 61.765 165.005 62.170 165.175 ;
        RECT 58.845 164.675 59.070 164.715 ;
        RECT 58.845 164.095 59.015 164.675 ;
        RECT 59.735 164.545 59.935 164.715 ;
        RECT 60.810 164.545 60.980 165.005 ;
        RECT 59.185 164.215 59.935 164.545 ;
        RECT 60.105 164.215 60.980 164.545 ;
        RECT 58.845 164.045 59.060 164.095 ;
        RECT 58.845 163.965 59.235 164.045 ;
        RECT 57.695 162.905 58.025 163.625 ;
        RECT 58.215 163.075 58.675 163.625 ;
        RECT 58.905 163.120 59.235 163.965 ;
        RECT 59.745 164.010 59.935 164.215 ;
        RECT 59.405 162.905 59.575 163.915 ;
        RECT 59.745 163.635 60.640 164.010 ;
        RECT 59.745 163.075 60.085 163.635 ;
        RECT 60.315 162.905 60.630 163.405 ;
        RECT 60.810 163.375 60.980 164.215 ;
        RECT 61.150 164.505 61.615 164.835 ;
        RECT 62.000 164.775 62.170 165.005 ;
        RECT 62.350 164.955 62.720 165.455 ;
        RECT 63.040 165.005 63.715 165.175 ;
        RECT 63.910 165.005 64.245 165.175 ;
        RECT 61.150 163.545 61.470 164.505 ;
        RECT 62.000 164.475 62.830 164.775 ;
        RECT 61.640 163.575 61.830 164.295 ;
        RECT 62.000 163.405 62.170 164.475 ;
        RECT 62.630 164.445 62.830 164.475 ;
        RECT 62.340 164.225 62.510 164.295 ;
        RECT 63.040 164.225 63.210 165.005 ;
        RECT 64.075 164.865 64.245 165.005 ;
        RECT 64.415 164.995 64.665 165.455 ;
        RECT 62.340 164.055 63.210 164.225 ;
        RECT 63.380 164.585 63.905 164.805 ;
        RECT 64.075 164.735 64.300 164.865 ;
        RECT 62.340 163.965 62.850 164.055 ;
        RECT 60.810 163.205 61.695 163.375 ;
        RECT 61.920 163.075 62.170 163.405 ;
        RECT 62.340 162.905 62.510 163.705 ;
        RECT 62.680 163.350 62.850 163.965 ;
        RECT 63.380 163.885 63.550 164.585 ;
        RECT 63.020 163.520 63.550 163.885 ;
        RECT 63.720 163.820 63.960 164.415 ;
        RECT 64.130 163.630 64.300 164.735 ;
        RECT 64.470 163.875 64.750 164.825 ;
        RECT 63.995 163.500 64.300 163.630 ;
        RECT 62.680 163.180 63.785 163.350 ;
        RECT 63.995 163.075 64.245 163.500 ;
        RECT 64.415 162.905 64.680 163.365 ;
        RECT 64.920 163.075 65.105 165.195 ;
        RECT 65.275 165.075 65.605 165.455 ;
        RECT 65.775 164.905 65.945 165.195 ;
        RECT 65.280 164.735 65.945 164.905 ;
        RECT 67.125 164.825 67.465 165.285 ;
        RECT 67.635 164.995 67.805 165.455 ;
        RECT 68.435 165.020 68.795 165.285 ;
        RECT 68.440 165.015 68.795 165.020 ;
        RECT 68.445 165.005 68.795 165.015 ;
        RECT 68.450 165.000 68.795 165.005 ;
        RECT 68.455 164.990 68.795 165.000 ;
        RECT 69.035 164.995 69.205 165.455 ;
        RECT 68.460 164.985 68.795 164.990 ;
        RECT 68.470 164.975 68.795 164.985 ;
        RECT 68.480 164.965 68.795 164.975 ;
        RECT 67.975 164.825 68.305 164.905 ;
        RECT 65.280 163.745 65.510 164.735 ;
        RECT 67.125 164.635 68.305 164.825 ;
        RECT 68.495 164.825 68.795 164.965 ;
        RECT 68.495 164.635 69.205 164.825 ;
        RECT 65.680 163.915 66.030 164.565 ;
        RECT 67.125 164.265 67.455 164.465 ;
        RECT 67.765 164.445 68.095 164.465 ;
        RECT 67.645 164.265 68.095 164.445 ;
        RECT 67.125 163.925 67.355 164.265 ;
        RECT 65.280 163.575 65.945 163.745 ;
        RECT 65.275 162.905 65.605 163.405 ;
        RECT 65.775 163.075 65.945 163.575 ;
        RECT 67.135 162.905 67.465 163.625 ;
        RECT 67.645 163.150 67.860 164.265 ;
        RECT 68.265 164.235 68.735 164.465 ;
        RECT 68.920 164.065 69.205 164.635 ;
        RECT 69.375 164.510 69.715 165.285 ;
        RECT 69.885 164.730 70.175 165.455 ;
        RECT 70.435 164.905 70.605 165.195 ;
        RECT 70.775 165.075 71.105 165.455 ;
        RECT 70.435 164.735 71.100 164.905 ;
        RECT 68.055 163.850 69.205 164.065 ;
        RECT 68.055 163.075 68.385 163.850 ;
        RECT 68.555 162.905 69.265 163.680 ;
        RECT 69.435 163.075 69.715 164.510 ;
        RECT 69.885 162.905 70.175 164.070 ;
        RECT 70.350 163.915 70.700 164.565 ;
        RECT 70.870 163.745 71.100 164.735 ;
        RECT 70.435 163.575 71.100 163.745 ;
        RECT 70.435 163.075 70.605 163.575 ;
        RECT 70.775 162.905 71.105 163.405 ;
        RECT 71.275 163.075 71.460 165.195 ;
        RECT 71.715 164.995 71.965 165.455 ;
        RECT 72.135 165.005 72.470 165.175 ;
        RECT 72.665 165.005 73.340 165.175 ;
        RECT 72.135 164.865 72.305 165.005 ;
        RECT 71.630 163.875 71.910 164.825 ;
        RECT 72.080 164.735 72.305 164.865 ;
        RECT 72.080 163.630 72.250 164.735 ;
        RECT 72.475 164.585 73.000 164.805 ;
        RECT 72.420 163.820 72.660 164.415 ;
        RECT 72.830 163.885 73.000 164.585 ;
        RECT 73.170 164.225 73.340 165.005 ;
        RECT 73.660 164.955 74.030 165.455 ;
        RECT 74.210 165.005 74.615 165.175 ;
        RECT 74.785 165.005 75.570 165.175 ;
        RECT 74.210 164.775 74.380 165.005 ;
        RECT 73.550 164.475 74.380 164.775 ;
        RECT 74.765 164.505 75.230 164.835 ;
        RECT 73.550 164.445 73.750 164.475 ;
        RECT 73.870 164.225 74.040 164.295 ;
        RECT 73.170 164.055 74.040 164.225 ;
        RECT 73.530 163.965 74.040 164.055 ;
        RECT 72.080 163.500 72.385 163.630 ;
        RECT 72.830 163.520 73.360 163.885 ;
        RECT 71.700 162.905 71.965 163.365 ;
        RECT 72.135 163.075 72.385 163.500 ;
        RECT 73.530 163.350 73.700 163.965 ;
        RECT 72.595 163.180 73.700 163.350 ;
        RECT 73.870 162.905 74.040 163.705 ;
        RECT 74.210 163.405 74.380 164.475 ;
        RECT 74.550 163.575 74.740 164.295 ;
        RECT 74.910 163.545 75.230 164.505 ;
        RECT 75.400 164.545 75.570 165.005 ;
        RECT 75.845 164.925 76.055 165.455 ;
        RECT 76.315 164.715 76.645 165.240 ;
        RECT 76.815 164.845 76.985 165.455 ;
        RECT 77.155 164.800 77.485 165.235 ;
        RECT 77.155 164.715 77.535 164.800 ;
        RECT 76.445 164.545 76.645 164.715 ;
        RECT 77.310 164.675 77.535 164.715 ;
        RECT 75.400 164.215 76.275 164.545 ;
        RECT 76.445 164.215 77.195 164.545 ;
        RECT 74.210 163.075 74.460 163.405 ;
        RECT 75.400 163.375 75.570 164.215 ;
        RECT 76.445 164.010 76.635 164.215 ;
        RECT 77.365 164.095 77.535 164.675 ;
        RECT 77.795 164.585 77.965 165.150 ;
        RECT 78.155 164.925 78.385 165.230 ;
        RECT 78.555 165.095 78.885 165.455 ;
        RECT 79.080 164.925 79.370 165.275 ;
        RECT 78.155 164.755 79.370 164.925 ;
        RECT 80.470 164.925 80.760 165.275 ;
        RECT 80.955 165.095 81.285 165.455 ;
        RECT 81.455 164.925 81.685 165.230 ;
        RECT 80.470 164.755 81.685 164.925 ;
        RECT 81.875 164.585 82.045 165.150 ;
        RECT 82.395 164.905 82.565 165.195 ;
        RECT 82.735 165.075 83.065 165.455 ;
        RECT 82.395 164.735 83.060 164.905 ;
        RECT 77.795 164.415 78.315 164.585 ;
        RECT 77.320 164.045 77.535 164.095 ;
        RECT 75.740 163.635 76.635 164.010 ;
        RECT 77.145 163.965 77.535 164.045 ;
        RECT 74.685 163.205 75.570 163.375 ;
        RECT 75.750 162.905 76.065 163.405 ;
        RECT 76.295 163.075 76.635 163.635 ;
        RECT 76.805 162.905 76.975 163.915 ;
        RECT 77.145 163.120 77.475 163.965 ;
        RECT 77.710 163.885 77.955 164.245 ;
        RECT 78.145 164.035 78.315 164.415 ;
        RECT 78.485 164.215 78.870 164.545 ;
        RECT 79.050 164.435 79.310 164.545 ;
        RECT 80.530 164.435 80.790 164.545 ;
        RECT 79.050 164.265 79.315 164.435 ;
        RECT 80.525 164.265 80.790 164.435 ;
        RECT 79.050 164.215 79.310 164.265 ;
        RECT 80.530 164.215 80.790 164.265 ;
        RECT 80.970 164.215 81.355 164.545 ;
        RECT 81.525 164.415 82.045 164.585 ;
        RECT 78.145 163.755 78.495 164.035 ;
        RECT 77.710 162.905 77.965 163.705 ;
        RECT 78.165 163.075 78.495 163.755 ;
        RECT 78.675 163.165 78.870 164.215 ;
        RECT 79.050 162.905 79.370 164.045 ;
        RECT 80.470 162.905 80.790 164.045 ;
        RECT 80.970 163.165 81.165 164.215 ;
        RECT 81.525 164.035 81.695 164.415 ;
        RECT 81.345 163.755 81.695 164.035 ;
        RECT 81.885 163.885 82.130 164.245 ;
        RECT 82.310 163.915 82.660 164.565 ;
        RECT 81.345 163.075 81.675 163.755 ;
        RECT 82.830 163.745 83.060 164.735 ;
        RECT 81.875 162.905 82.130 163.705 ;
        RECT 82.395 163.575 83.060 163.745 ;
        RECT 82.395 163.075 82.565 163.575 ;
        RECT 82.735 162.905 83.065 163.405 ;
        RECT 83.235 163.075 83.460 165.195 ;
        RECT 83.675 164.995 83.925 165.455 ;
        RECT 84.110 165.005 84.440 165.175 ;
        RECT 84.620 165.005 85.370 165.175 ;
        RECT 83.660 163.875 83.940 164.475 ;
        RECT 84.110 163.475 84.280 165.005 ;
        RECT 84.450 164.505 85.030 164.835 ;
        RECT 84.450 163.635 84.690 164.505 ;
        RECT 85.200 164.225 85.370 165.005 ;
        RECT 85.620 164.955 85.990 165.455 ;
        RECT 86.170 165.005 86.630 165.175 ;
        RECT 86.860 165.005 87.530 165.175 ;
        RECT 86.170 164.775 86.340 165.005 ;
        RECT 85.540 164.475 86.340 164.775 ;
        RECT 86.510 164.505 87.060 164.835 ;
        RECT 85.540 164.445 85.710 164.475 ;
        RECT 85.830 164.225 86.000 164.295 ;
        RECT 85.200 164.055 86.000 164.225 ;
        RECT 85.490 163.965 86.000 164.055 ;
        RECT 84.880 163.530 85.320 163.885 ;
        RECT 83.660 162.905 83.925 163.365 ;
        RECT 84.110 163.100 84.345 163.475 ;
        RECT 85.490 163.350 85.660 163.965 ;
        RECT 84.590 163.180 85.660 163.350 ;
        RECT 85.830 162.905 86.000 163.705 ;
        RECT 86.170 163.405 86.340 164.475 ;
        RECT 86.510 163.575 86.700 164.295 ;
        RECT 86.870 163.965 87.060 164.505 ;
        RECT 87.360 164.465 87.530 165.005 ;
        RECT 87.845 164.925 88.015 165.455 ;
        RECT 88.310 164.805 88.670 165.245 ;
        RECT 88.845 164.975 89.015 165.455 ;
        RECT 89.205 164.810 89.540 165.235 ;
        RECT 89.715 164.980 89.885 165.455 ;
        RECT 90.060 164.810 90.395 165.235 ;
        RECT 90.565 164.980 90.735 165.455 ;
        RECT 88.310 164.635 88.810 164.805 ;
        RECT 89.205 164.640 90.875 164.810 ;
        RECT 91.045 164.705 92.255 165.455 ;
        RECT 88.640 164.465 88.810 164.635 ;
        RECT 87.360 164.295 88.450 164.465 ;
        RECT 88.640 164.295 90.460 164.465 ;
        RECT 86.870 163.635 87.190 163.965 ;
        RECT 86.170 163.075 86.420 163.405 ;
        RECT 87.360 163.375 87.530 164.295 ;
        RECT 88.640 164.040 88.810 164.295 ;
        RECT 90.630 164.075 90.875 164.640 ;
        RECT 87.700 163.870 88.810 164.040 ;
        RECT 89.205 163.905 90.875 164.075 ;
        RECT 91.045 163.995 91.565 164.535 ;
        RECT 91.735 164.165 92.255 164.705 ;
        RECT 87.700 163.710 88.560 163.870 ;
        RECT 86.645 163.205 87.530 163.375 ;
        RECT 87.710 162.905 87.925 163.405 ;
        RECT 88.390 163.085 88.560 163.710 ;
        RECT 88.845 162.905 89.025 163.685 ;
        RECT 89.205 163.145 89.540 163.905 ;
        RECT 89.720 162.905 89.890 163.735 ;
        RECT 90.060 163.145 90.390 163.905 ;
        RECT 90.560 162.905 90.730 163.735 ;
        RECT 91.045 162.905 92.255 163.995 ;
        RECT 18.280 162.735 92.340 162.905 ;
        RECT 18.365 161.645 19.575 162.735 ;
        RECT 19.745 162.300 25.090 162.735 ;
        RECT 25.265 162.300 30.610 162.735 ;
        RECT 18.365 160.935 18.885 161.475 ;
        RECT 19.055 161.105 19.575 161.645 ;
        RECT 18.365 160.185 19.575 160.935 ;
        RECT 21.330 160.730 21.670 161.560 ;
        RECT 23.150 161.050 23.500 162.300 ;
        RECT 26.850 160.730 27.190 161.560 ;
        RECT 28.670 161.050 29.020 162.300 ;
        RECT 31.245 161.570 31.535 162.735 ;
        RECT 31.705 161.645 35.215 162.735 ;
        RECT 36.395 162.065 36.565 162.565 ;
        RECT 36.735 162.235 37.065 162.735 ;
        RECT 36.395 161.895 37.060 162.065 ;
        RECT 31.705 160.955 33.355 161.475 ;
        RECT 33.525 161.125 35.215 161.645 ;
        RECT 36.310 161.075 36.660 161.725 ;
        RECT 19.745 160.185 25.090 160.730 ;
        RECT 25.265 160.185 30.610 160.730 ;
        RECT 31.245 160.185 31.535 160.910 ;
        RECT 31.705 160.185 35.215 160.955 ;
        RECT 36.830 160.905 37.060 161.895 ;
        RECT 36.395 160.735 37.060 160.905 ;
        RECT 36.395 160.445 36.565 160.735 ;
        RECT 36.735 160.185 37.065 160.565 ;
        RECT 37.235 160.445 37.420 162.565 ;
        RECT 37.660 162.275 37.925 162.735 ;
        RECT 38.095 162.140 38.345 162.565 ;
        RECT 38.555 162.290 39.660 162.460 ;
        RECT 38.040 162.010 38.345 162.140 ;
        RECT 37.590 160.815 37.870 161.765 ;
        RECT 38.040 160.905 38.210 162.010 ;
        RECT 38.380 161.225 38.620 161.820 ;
        RECT 38.790 161.755 39.320 162.120 ;
        RECT 38.790 161.055 38.960 161.755 ;
        RECT 39.490 161.675 39.660 162.290 ;
        RECT 39.830 161.935 40.000 162.735 ;
        RECT 40.170 162.235 40.420 162.565 ;
        RECT 40.645 162.265 41.530 162.435 ;
        RECT 39.490 161.585 40.000 161.675 ;
        RECT 38.040 160.775 38.265 160.905 ;
        RECT 38.435 160.835 38.960 161.055 ;
        RECT 39.130 161.415 40.000 161.585 ;
        RECT 37.675 160.185 37.925 160.645 ;
        RECT 38.095 160.635 38.265 160.775 ;
        RECT 39.130 160.635 39.300 161.415 ;
        RECT 39.830 161.345 40.000 161.415 ;
        RECT 39.510 161.165 39.710 161.195 ;
        RECT 40.170 161.165 40.340 162.235 ;
        RECT 40.510 161.345 40.700 162.065 ;
        RECT 39.510 160.865 40.340 161.165 ;
        RECT 40.870 161.135 41.190 162.095 ;
        RECT 38.095 160.465 38.430 160.635 ;
        RECT 38.625 160.465 39.300 160.635 ;
        RECT 39.620 160.185 39.990 160.685 ;
        RECT 40.170 160.635 40.340 160.865 ;
        RECT 40.725 160.805 41.190 161.135 ;
        RECT 41.360 161.425 41.530 162.265 ;
        RECT 41.710 162.235 42.025 162.735 ;
        RECT 42.255 162.005 42.595 162.565 ;
        RECT 41.700 161.630 42.595 162.005 ;
        RECT 42.765 161.725 42.935 162.735 ;
        RECT 42.405 161.425 42.595 161.630 ;
        RECT 43.105 161.675 43.435 162.520 ;
        RECT 43.105 161.595 43.495 161.675 ;
        RECT 43.665 161.645 46.255 162.735 ;
        RECT 43.280 161.545 43.495 161.595 ;
        RECT 41.360 161.095 42.235 161.425 ;
        RECT 42.405 161.095 43.155 161.425 ;
        RECT 41.360 160.635 41.530 161.095 ;
        RECT 42.405 160.925 42.605 161.095 ;
        RECT 43.325 160.965 43.495 161.545 ;
        RECT 43.270 160.925 43.495 160.965 ;
        RECT 40.170 160.465 40.575 160.635 ;
        RECT 40.745 160.465 41.530 160.635 ;
        RECT 41.805 160.185 42.015 160.715 ;
        RECT 42.275 160.400 42.605 160.925 ;
        RECT 43.115 160.840 43.495 160.925 ;
        RECT 43.665 160.955 44.875 161.475 ;
        RECT 45.045 161.125 46.255 161.645 ;
        RECT 46.925 161.595 47.155 162.735 ;
        RECT 47.325 161.585 47.655 162.565 ;
        RECT 47.825 161.595 48.035 162.735 ;
        RECT 48.265 161.645 50.855 162.735 ;
        RECT 46.905 161.175 47.235 161.425 ;
        RECT 42.775 160.185 42.945 160.795 ;
        RECT 43.115 160.405 43.445 160.840 ;
        RECT 43.665 160.185 46.255 160.955 ;
        RECT 46.925 160.185 47.155 161.005 ;
        RECT 47.405 160.985 47.655 161.585 ;
        RECT 47.325 160.355 47.655 160.985 ;
        RECT 47.825 160.185 48.035 161.005 ;
        RECT 48.265 160.955 49.475 161.475 ;
        RECT 49.645 161.125 50.855 161.645 ;
        RECT 51.485 161.865 51.760 162.565 ;
        RECT 51.930 162.190 52.185 162.735 ;
        RECT 52.355 162.225 52.835 162.565 ;
        RECT 53.010 162.180 53.615 162.735 ;
        RECT 53.000 162.080 53.615 162.180 ;
        RECT 53.000 162.055 53.185 162.080 ;
        RECT 48.265 160.185 50.855 160.955 ;
        RECT 51.485 160.835 51.655 161.865 ;
        RECT 51.930 161.735 52.685 161.985 ;
        RECT 52.855 161.810 53.185 162.055 ;
        RECT 51.930 161.700 52.700 161.735 ;
        RECT 51.930 161.690 52.715 161.700 ;
        RECT 51.825 161.675 52.720 161.690 ;
        RECT 51.825 161.660 52.740 161.675 ;
        RECT 51.825 161.650 52.760 161.660 ;
        RECT 51.825 161.640 52.785 161.650 ;
        RECT 51.825 161.610 52.855 161.640 ;
        RECT 51.825 161.580 52.875 161.610 ;
        RECT 51.825 161.550 52.895 161.580 ;
        RECT 51.825 161.525 52.925 161.550 ;
        RECT 51.825 161.490 52.960 161.525 ;
        RECT 51.825 161.485 52.990 161.490 ;
        RECT 51.825 161.090 52.055 161.485 ;
        RECT 52.600 161.480 52.990 161.485 ;
        RECT 52.625 161.470 52.990 161.480 ;
        RECT 52.640 161.465 52.990 161.470 ;
        RECT 52.655 161.460 52.990 161.465 ;
        RECT 53.355 161.460 53.615 161.910 ;
        RECT 53.795 161.765 54.125 162.550 ;
        RECT 53.795 161.595 54.475 161.765 ;
        RECT 54.655 161.595 54.985 162.735 ;
        RECT 55.165 161.645 56.835 162.735 ;
        RECT 52.655 161.455 53.615 161.460 ;
        RECT 52.665 161.445 53.615 161.455 ;
        RECT 52.675 161.440 53.615 161.445 ;
        RECT 52.685 161.430 53.615 161.440 ;
        RECT 52.690 161.420 53.615 161.430 ;
        RECT 52.695 161.415 53.615 161.420 ;
        RECT 52.705 161.400 53.615 161.415 ;
        RECT 52.710 161.385 53.615 161.400 ;
        RECT 52.720 161.360 53.615 161.385 ;
        RECT 52.225 160.890 52.555 161.315 ;
        RECT 51.485 160.355 51.745 160.835 ;
        RECT 51.915 160.185 52.165 160.725 ;
        RECT 52.335 160.405 52.555 160.890 ;
        RECT 52.725 161.290 53.615 161.360 ;
        RECT 52.725 160.565 52.895 161.290 ;
        RECT 53.785 161.175 54.135 161.425 ;
        RECT 53.065 160.735 53.615 161.120 ;
        RECT 54.305 160.995 54.475 161.595 ;
        RECT 54.645 161.175 54.995 161.425 ;
        RECT 52.725 160.395 53.615 160.565 ;
        RECT 53.805 160.185 54.045 160.995 ;
        RECT 54.215 160.355 54.545 160.995 ;
        RECT 54.715 160.185 54.985 160.995 ;
        RECT 55.165 160.955 55.915 161.475 ;
        RECT 56.085 161.125 56.835 161.645 ;
        RECT 57.005 161.570 57.295 162.735 ;
        RECT 57.465 161.765 57.775 162.565 ;
        RECT 57.945 161.935 58.255 162.735 ;
        RECT 58.425 162.105 58.685 162.565 ;
        RECT 58.855 162.275 59.110 162.735 ;
        RECT 59.285 162.105 59.545 162.565 ;
        RECT 58.425 161.935 59.545 162.105 ;
        RECT 57.465 161.595 58.495 161.765 ;
        RECT 55.165 160.185 56.835 160.955 ;
        RECT 57.005 160.185 57.295 160.910 ;
        RECT 57.465 160.685 57.635 161.595 ;
        RECT 57.805 160.855 58.155 161.425 ;
        RECT 58.325 161.345 58.495 161.595 ;
        RECT 59.285 161.685 59.545 161.935 ;
        RECT 59.715 161.865 60.000 162.735 ;
        RECT 60.315 161.805 60.485 162.565 ;
        RECT 60.665 161.975 60.995 162.735 ;
        RECT 59.285 161.515 60.040 161.685 ;
        RECT 60.315 161.635 60.980 161.805 ;
        RECT 61.165 161.660 61.435 162.565 ;
        RECT 61.605 162.300 66.950 162.735 ;
        RECT 58.325 161.175 59.465 161.345 ;
        RECT 59.635 161.005 60.040 161.515 ;
        RECT 60.810 161.490 60.980 161.635 ;
        RECT 60.245 161.085 60.575 161.455 ;
        RECT 60.810 161.160 61.095 161.490 ;
        RECT 58.390 160.835 60.040 161.005 ;
        RECT 60.810 160.905 60.980 161.160 ;
        RECT 57.465 160.355 57.765 160.685 ;
        RECT 57.935 160.185 58.210 160.665 ;
        RECT 58.390 160.445 58.685 160.835 ;
        RECT 58.855 160.185 59.110 160.665 ;
        RECT 59.285 160.445 59.545 160.835 ;
        RECT 60.315 160.735 60.980 160.905 ;
        RECT 61.265 160.860 61.435 161.660 ;
        RECT 59.715 160.185 59.995 160.665 ;
        RECT 60.315 160.355 60.485 160.735 ;
        RECT 60.665 160.185 60.995 160.565 ;
        RECT 61.175 160.355 61.435 160.860 ;
        RECT 63.190 160.730 63.530 161.560 ;
        RECT 65.010 161.050 65.360 162.300 ;
        RECT 67.125 161.645 68.335 162.735 ;
        RECT 67.125 160.935 67.645 161.475 ;
        RECT 67.815 161.105 68.335 161.645 ;
        RECT 68.515 161.785 68.790 162.555 ;
        RECT 68.960 162.125 69.290 162.555 ;
        RECT 69.460 162.295 69.655 162.735 ;
        RECT 69.835 162.125 70.165 162.555 ;
        RECT 70.345 162.300 75.690 162.735 ;
        RECT 68.960 161.955 70.165 162.125 ;
        RECT 68.515 161.595 69.100 161.785 ;
        RECT 69.270 161.625 70.165 161.955 ;
        RECT 61.605 160.185 66.950 160.730 ;
        RECT 67.125 160.185 68.335 160.935 ;
        RECT 68.515 160.775 68.755 161.425 ;
        RECT 68.925 160.925 69.100 161.595 ;
        RECT 69.270 161.095 69.685 161.425 ;
        RECT 69.865 161.095 70.160 161.425 ;
        RECT 68.925 160.745 69.255 160.925 ;
        RECT 68.530 160.185 68.860 160.575 ;
        RECT 69.030 160.365 69.255 160.745 ;
        RECT 69.455 160.475 69.685 161.095 ;
        RECT 69.865 160.185 70.165 160.915 ;
        RECT 71.930 160.730 72.270 161.560 ;
        RECT 73.750 161.050 74.100 162.300 ;
        RECT 76.325 161.595 76.605 162.735 ;
        RECT 76.775 161.585 77.105 162.565 ;
        RECT 77.275 161.595 77.535 162.735 ;
        RECT 77.715 162.125 78.045 162.555 ;
        RECT 78.225 162.295 78.420 162.735 ;
        RECT 78.590 162.125 78.920 162.555 ;
        RECT 77.715 161.955 78.920 162.125 ;
        RECT 77.715 161.625 78.610 161.955 ;
        RECT 79.090 161.785 79.365 162.555 ;
        RECT 78.780 161.595 79.365 161.785 ;
        RECT 79.545 161.645 82.135 162.735 ;
        RECT 76.335 161.155 76.670 161.425 ;
        RECT 76.840 160.985 77.010 161.585 ;
        RECT 77.180 161.175 77.515 161.425 ;
        RECT 77.720 161.095 78.015 161.425 ;
        RECT 78.195 161.095 78.610 161.425 ;
        RECT 70.345 160.185 75.690 160.730 ;
        RECT 76.325 160.185 76.635 160.985 ;
        RECT 76.840 160.355 77.535 160.985 ;
        RECT 77.715 160.185 78.015 160.915 ;
        RECT 78.195 160.475 78.425 161.095 ;
        RECT 78.780 160.925 78.955 161.595 ;
        RECT 78.625 160.745 78.955 160.925 ;
        RECT 79.125 160.775 79.365 161.425 ;
        RECT 79.545 160.955 80.755 161.475 ;
        RECT 80.925 161.125 82.135 161.645 ;
        RECT 82.765 161.570 83.055 162.735 ;
        RECT 83.235 161.785 83.510 162.555 ;
        RECT 83.680 162.125 84.010 162.555 ;
        RECT 84.180 162.295 84.375 162.735 ;
        RECT 84.555 162.125 84.885 162.555 ;
        RECT 85.065 162.300 90.410 162.735 ;
        RECT 83.680 161.955 84.885 162.125 ;
        RECT 83.235 161.595 83.820 161.785 ;
        RECT 83.990 161.625 84.885 161.955 ;
        RECT 78.625 160.365 78.850 160.745 ;
        RECT 79.020 160.185 79.350 160.575 ;
        RECT 79.545 160.185 82.135 160.955 ;
        RECT 82.765 160.185 83.055 160.910 ;
        RECT 83.235 160.775 83.475 161.425 ;
        RECT 83.645 160.925 83.820 161.595 ;
        RECT 83.990 161.095 84.405 161.425 ;
        RECT 84.585 161.095 84.880 161.425 ;
        RECT 83.645 160.745 83.975 160.925 ;
        RECT 83.250 160.185 83.580 160.575 ;
        RECT 83.750 160.365 83.975 160.745 ;
        RECT 84.175 160.475 84.405 161.095 ;
        RECT 84.585 160.185 84.885 160.915 ;
        RECT 86.650 160.730 86.990 161.560 ;
        RECT 88.470 161.050 88.820 162.300 ;
        RECT 91.045 161.645 92.255 162.735 ;
        RECT 91.045 161.105 91.565 161.645 ;
        RECT 91.735 160.935 92.255 161.475 ;
        RECT 85.065 160.185 90.410 160.730 ;
        RECT 91.045 160.185 92.255 160.935 ;
        RECT 18.280 160.015 92.340 160.185 ;
        RECT 18.365 159.265 19.575 160.015 ;
        RECT 19.745 159.470 25.090 160.015 ;
        RECT 25.265 159.470 30.610 160.015 ;
        RECT 30.785 159.470 36.130 160.015 ;
        RECT 18.365 158.725 18.885 159.265 ;
        RECT 19.055 158.555 19.575 159.095 ;
        RECT 21.330 158.640 21.670 159.470 ;
        RECT 18.365 157.465 19.575 158.555 ;
        RECT 23.150 157.900 23.500 159.150 ;
        RECT 26.850 158.640 27.190 159.470 ;
        RECT 28.670 157.900 29.020 159.150 ;
        RECT 32.370 158.640 32.710 159.470 ;
        RECT 36.855 159.465 37.025 159.755 ;
        RECT 37.195 159.635 37.525 160.015 ;
        RECT 36.855 159.295 37.520 159.465 ;
        RECT 34.190 157.900 34.540 159.150 ;
        RECT 36.770 158.475 37.120 159.125 ;
        RECT 37.290 158.305 37.520 159.295 ;
        RECT 36.855 158.135 37.520 158.305 ;
        RECT 19.745 157.465 25.090 157.900 ;
        RECT 25.265 157.465 30.610 157.900 ;
        RECT 30.785 157.465 36.130 157.900 ;
        RECT 36.855 157.635 37.025 158.135 ;
        RECT 37.195 157.465 37.525 157.965 ;
        RECT 37.695 157.635 37.880 159.755 ;
        RECT 38.135 159.555 38.385 160.015 ;
        RECT 38.555 159.565 38.890 159.735 ;
        RECT 39.085 159.565 39.760 159.735 ;
        RECT 38.555 159.425 38.725 159.565 ;
        RECT 38.050 158.435 38.330 159.385 ;
        RECT 38.500 159.295 38.725 159.425 ;
        RECT 38.500 158.190 38.670 159.295 ;
        RECT 38.895 159.145 39.420 159.365 ;
        RECT 38.840 158.380 39.080 158.975 ;
        RECT 39.250 158.445 39.420 159.145 ;
        RECT 39.590 158.785 39.760 159.565 ;
        RECT 40.080 159.515 40.450 160.015 ;
        RECT 40.630 159.565 41.035 159.735 ;
        RECT 41.205 159.565 41.990 159.735 ;
        RECT 40.630 159.335 40.800 159.565 ;
        RECT 39.970 159.035 40.800 159.335 ;
        RECT 41.185 159.065 41.650 159.395 ;
        RECT 39.970 159.005 40.170 159.035 ;
        RECT 40.290 158.785 40.460 158.855 ;
        RECT 39.590 158.615 40.460 158.785 ;
        RECT 39.950 158.525 40.460 158.615 ;
        RECT 38.500 158.060 38.805 158.190 ;
        RECT 39.250 158.080 39.780 158.445 ;
        RECT 38.120 157.465 38.385 157.925 ;
        RECT 38.555 157.635 38.805 158.060 ;
        RECT 39.950 157.910 40.120 158.525 ;
        RECT 39.015 157.740 40.120 157.910 ;
        RECT 40.290 157.465 40.460 158.265 ;
        RECT 40.630 157.965 40.800 159.035 ;
        RECT 40.970 158.135 41.160 158.855 ;
        RECT 41.330 158.105 41.650 159.065 ;
        RECT 41.820 159.105 41.990 159.565 ;
        RECT 42.265 159.485 42.475 160.015 ;
        RECT 42.735 159.275 43.065 159.800 ;
        RECT 43.235 159.405 43.405 160.015 ;
        RECT 43.575 159.360 43.905 159.795 ;
        RECT 43.575 159.275 43.955 159.360 ;
        RECT 44.125 159.290 44.415 160.015 ;
        RECT 44.675 159.535 44.975 160.015 ;
        RECT 45.145 159.365 45.405 159.820 ;
        RECT 45.575 159.535 45.835 160.015 ;
        RECT 46.015 159.365 46.275 159.820 ;
        RECT 46.445 159.535 46.695 160.015 ;
        RECT 46.875 159.365 47.135 159.820 ;
        RECT 47.305 159.535 47.555 160.015 ;
        RECT 47.735 159.365 47.995 159.820 ;
        RECT 48.165 159.535 48.410 160.015 ;
        RECT 48.580 159.365 48.855 159.820 ;
        RECT 49.025 159.535 49.270 160.015 ;
        RECT 49.440 159.365 49.700 159.820 ;
        RECT 49.870 159.535 50.130 160.015 ;
        RECT 50.300 159.365 50.560 159.820 ;
        RECT 50.730 159.535 50.990 160.015 ;
        RECT 51.160 159.365 51.420 159.820 ;
        RECT 51.590 159.455 51.850 160.015 ;
        RECT 42.865 159.105 43.065 159.275 ;
        RECT 43.730 159.235 43.955 159.275 ;
        RECT 41.820 158.775 42.695 159.105 ;
        RECT 42.865 158.775 43.615 159.105 ;
        RECT 40.630 157.635 40.880 157.965 ;
        RECT 41.820 157.935 41.990 158.775 ;
        RECT 42.865 158.570 43.055 158.775 ;
        RECT 43.785 158.655 43.955 159.235 ;
        RECT 43.740 158.605 43.955 158.655 ;
        RECT 44.675 159.195 51.420 159.365 ;
        RECT 42.160 158.195 43.055 158.570 ;
        RECT 43.565 158.525 43.955 158.605 ;
        RECT 41.105 157.765 41.990 157.935 ;
        RECT 42.170 157.465 42.485 157.965 ;
        RECT 42.715 157.635 43.055 158.195 ;
        RECT 43.225 157.465 43.395 158.475 ;
        RECT 43.565 157.680 43.895 158.525 ;
        RECT 44.125 157.465 44.415 158.630 ;
        RECT 44.675 158.605 45.840 159.195 ;
        RECT 52.020 159.025 52.270 159.835 ;
        RECT 52.450 159.490 52.710 160.015 ;
        RECT 52.880 159.025 53.130 159.835 ;
        RECT 53.310 159.505 53.615 160.015 ;
        RECT 54.795 159.465 54.965 159.845 ;
        RECT 55.180 159.635 55.510 160.015 ;
        RECT 46.010 158.775 53.130 159.025 ;
        RECT 53.300 158.775 53.615 159.335 ;
        RECT 54.795 159.295 55.510 159.465 ;
        RECT 44.675 158.380 51.420 158.605 ;
        RECT 44.675 157.465 44.945 158.210 ;
        RECT 45.115 157.640 45.405 158.380 ;
        RECT 46.015 158.365 51.420 158.380 ;
        RECT 45.575 157.470 45.830 158.195 ;
        RECT 46.015 157.640 46.275 158.365 ;
        RECT 46.445 157.470 46.690 158.195 ;
        RECT 46.875 157.640 47.135 158.365 ;
        RECT 47.305 157.470 47.550 158.195 ;
        RECT 47.735 157.640 47.995 158.365 ;
        RECT 48.165 157.470 48.410 158.195 ;
        RECT 48.580 157.640 48.840 158.365 ;
        RECT 49.010 157.470 49.270 158.195 ;
        RECT 49.440 157.640 49.700 158.365 ;
        RECT 49.870 157.470 50.130 158.195 ;
        RECT 50.300 157.640 50.560 158.365 ;
        RECT 50.730 157.470 50.990 158.195 ;
        RECT 51.160 157.640 51.420 158.365 ;
        RECT 51.590 157.470 51.850 158.265 ;
        RECT 52.020 157.640 52.270 158.775 ;
        RECT 45.575 157.465 51.850 157.470 ;
        RECT 52.450 157.465 52.710 158.275 ;
        RECT 52.885 157.635 53.130 158.775 ;
        RECT 54.705 158.745 55.060 159.115 ;
        RECT 55.340 159.105 55.510 159.295 ;
        RECT 55.680 159.270 55.935 159.845 ;
        RECT 55.340 158.775 55.595 159.105 ;
        RECT 55.340 158.565 55.510 158.775 ;
        RECT 54.795 158.395 55.510 158.565 ;
        RECT 55.765 158.540 55.935 159.270 ;
        RECT 56.110 159.175 56.370 160.015 ;
        RECT 56.545 159.470 61.890 160.015 ;
        RECT 62.065 159.470 67.410 160.015 ;
        RECT 58.130 158.640 58.470 159.470 ;
        RECT 53.310 157.465 53.605 158.275 ;
        RECT 54.795 157.635 54.965 158.395 ;
        RECT 55.180 157.465 55.510 158.225 ;
        RECT 55.680 157.635 55.935 158.540 ;
        RECT 56.110 157.465 56.370 158.615 ;
        RECT 59.950 157.900 60.300 159.150 ;
        RECT 63.650 158.640 63.990 159.470 ;
        RECT 67.585 159.245 69.255 160.015 ;
        RECT 69.885 159.290 70.175 160.015 ;
        RECT 70.345 159.505 70.650 160.015 ;
        RECT 65.470 157.900 65.820 159.150 ;
        RECT 67.585 158.725 68.335 159.245 ;
        RECT 68.505 158.555 69.255 159.075 ;
        RECT 70.345 158.775 70.660 159.335 ;
        RECT 70.830 159.025 71.080 159.835 ;
        RECT 71.250 159.490 71.510 160.015 ;
        RECT 71.690 159.025 71.940 159.835 ;
        RECT 72.110 159.455 72.370 160.015 ;
        RECT 72.540 159.365 72.800 159.820 ;
        RECT 72.970 159.535 73.230 160.015 ;
        RECT 73.400 159.365 73.660 159.820 ;
        RECT 73.830 159.535 74.090 160.015 ;
        RECT 74.260 159.365 74.520 159.820 ;
        RECT 74.690 159.535 74.935 160.015 ;
        RECT 75.105 159.365 75.380 159.820 ;
        RECT 75.550 159.535 75.795 160.015 ;
        RECT 75.965 159.365 76.225 159.820 ;
        RECT 76.405 159.535 76.655 160.015 ;
        RECT 76.825 159.365 77.085 159.820 ;
        RECT 77.265 159.535 77.515 160.015 ;
        RECT 77.685 159.365 77.945 159.820 ;
        RECT 78.125 159.535 78.385 160.015 ;
        RECT 78.555 159.365 78.815 159.820 ;
        RECT 78.985 159.535 79.285 160.015 ;
        RECT 79.635 159.465 79.805 159.755 ;
        RECT 79.975 159.635 80.305 160.015 ;
        RECT 72.540 159.195 79.285 159.365 ;
        RECT 79.635 159.295 80.300 159.465 ;
        RECT 70.830 158.775 77.950 159.025 ;
        RECT 78.120 158.995 79.285 159.195 ;
        RECT 78.120 158.825 79.315 158.995 ;
        RECT 56.545 157.465 61.890 157.900 ;
        RECT 62.065 157.465 67.410 157.900 ;
        RECT 67.585 157.465 69.255 158.555 ;
        RECT 69.885 157.465 70.175 158.630 ;
        RECT 70.355 157.465 70.650 158.275 ;
        RECT 70.830 157.635 71.075 158.775 ;
        RECT 71.250 157.465 71.510 158.275 ;
        RECT 71.690 157.640 71.940 158.775 ;
        RECT 78.120 158.605 79.285 158.825 ;
        RECT 72.540 158.380 79.285 158.605 ;
        RECT 79.550 158.475 79.900 159.125 ;
        RECT 72.540 158.365 77.945 158.380 ;
        RECT 72.110 157.470 72.370 158.265 ;
        RECT 72.540 157.640 72.800 158.365 ;
        RECT 72.970 157.470 73.230 158.195 ;
        RECT 73.400 157.640 73.660 158.365 ;
        RECT 73.830 157.470 74.090 158.195 ;
        RECT 74.260 157.640 74.520 158.365 ;
        RECT 74.690 157.470 74.950 158.195 ;
        RECT 75.120 157.640 75.380 158.365 ;
        RECT 75.550 157.470 75.795 158.195 ;
        RECT 75.965 157.640 76.225 158.365 ;
        RECT 76.410 157.470 76.655 158.195 ;
        RECT 76.825 157.640 77.085 158.365 ;
        RECT 77.270 157.470 77.515 158.195 ;
        RECT 77.685 157.640 77.945 158.365 ;
        RECT 78.130 157.470 78.385 158.195 ;
        RECT 78.555 157.640 78.845 158.380 ;
        RECT 80.070 158.305 80.300 159.295 ;
        RECT 72.110 157.465 78.385 157.470 ;
        RECT 79.015 157.465 79.285 158.210 ;
        RECT 79.635 158.135 80.300 158.305 ;
        RECT 79.635 157.635 79.805 158.135 ;
        RECT 79.975 157.465 80.305 157.965 ;
        RECT 80.475 157.635 80.700 159.755 ;
        RECT 80.915 159.555 81.165 160.015 ;
        RECT 81.350 159.565 81.680 159.735 ;
        RECT 81.860 159.565 82.610 159.735 ;
        RECT 80.900 158.435 81.180 159.035 ;
        RECT 81.350 158.035 81.520 159.565 ;
        RECT 81.690 159.065 82.270 159.395 ;
        RECT 81.690 158.195 81.930 159.065 ;
        RECT 82.440 158.785 82.610 159.565 ;
        RECT 82.860 159.515 83.230 160.015 ;
        RECT 83.410 159.565 83.870 159.735 ;
        RECT 84.100 159.565 84.770 159.735 ;
        RECT 83.410 159.335 83.580 159.565 ;
        RECT 82.780 159.035 83.580 159.335 ;
        RECT 83.750 159.065 84.300 159.395 ;
        RECT 82.780 159.005 82.950 159.035 ;
        RECT 83.070 158.785 83.240 158.855 ;
        RECT 82.440 158.615 83.240 158.785 ;
        RECT 82.730 158.525 83.240 158.615 ;
        RECT 82.120 158.090 82.560 158.445 ;
        RECT 80.900 157.465 81.165 157.925 ;
        RECT 81.350 157.660 81.585 158.035 ;
        RECT 82.730 157.910 82.900 158.525 ;
        RECT 81.830 157.740 82.900 157.910 ;
        RECT 83.070 157.465 83.240 158.265 ;
        RECT 83.410 157.965 83.580 159.035 ;
        RECT 83.750 158.135 83.940 158.855 ;
        RECT 84.110 158.525 84.300 159.065 ;
        RECT 84.600 159.025 84.770 159.565 ;
        RECT 85.085 159.485 85.255 160.015 ;
        RECT 85.550 159.365 85.910 159.805 ;
        RECT 86.085 159.535 86.255 160.015 ;
        RECT 86.445 159.370 86.780 159.795 ;
        RECT 86.955 159.540 87.125 160.015 ;
        RECT 87.300 159.370 87.635 159.795 ;
        RECT 87.805 159.540 87.975 160.015 ;
        RECT 85.550 159.195 86.050 159.365 ;
        RECT 86.445 159.200 88.115 159.370 ;
        RECT 85.880 159.025 86.050 159.195 ;
        RECT 84.600 158.855 85.690 159.025 ;
        RECT 85.880 158.855 87.700 159.025 ;
        RECT 84.110 158.195 84.430 158.525 ;
        RECT 83.410 157.635 83.660 157.965 ;
        RECT 84.600 157.935 84.770 158.855 ;
        RECT 85.880 158.600 86.050 158.855 ;
        RECT 87.870 158.635 88.115 159.200 ;
        RECT 88.285 159.245 90.875 160.015 ;
        RECT 91.045 159.265 92.255 160.015 ;
        RECT 88.285 158.725 89.495 159.245 ;
        RECT 84.940 158.430 86.050 158.600 ;
        RECT 86.445 158.465 88.115 158.635 ;
        RECT 89.665 158.555 90.875 159.075 ;
        RECT 84.940 158.270 85.800 158.430 ;
        RECT 83.885 157.765 84.770 157.935 ;
        RECT 84.950 157.465 85.165 157.965 ;
        RECT 85.630 157.645 85.800 158.270 ;
        RECT 86.085 157.465 86.265 158.245 ;
        RECT 86.445 157.705 86.780 158.465 ;
        RECT 86.960 157.465 87.130 158.295 ;
        RECT 87.300 157.705 87.630 158.465 ;
        RECT 87.800 157.465 87.970 158.295 ;
        RECT 88.285 157.465 90.875 158.555 ;
        RECT 91.045 158.555 91.565 159.095 ;
        RECT 91.735 158.725 92.255 159.265 ;
        RECT 91.045 157.465 92.255 158.555 ;
        RECT 18.280 157.295 92.340 157.465 ;
        RECT 18.365 156.205 19.575 157.295 ;
        RECT 19.745 156.860 25.090 157.295 ;
        RECT 25.265 156.860 30.610 157.295 ;
        RECT 18.365 155.495 18.885 156.035 ;
        RECT 19.055 155.665 19.575 156.205 ;
        RECT 18.365 154.745 19.575 155.495 ;
        RECT 21.330 155.290 21.670 156.120 ;
        RECT 23.150 155.610 23.500 156.860 ;
        RECT 26.850 155.290 27.190 156.120 ;
        RECT 28.670 155.610 29.020 156.860 ;
        RECT 31.245 156.130 31.535 157.295 ;
        RECT 31.705 156.860 37.050 157.295 ;
        RECT 37.225 156.860 42.570 157.295 ;
        RECT 19.745 154.745 25.090 155.290 ;
        RECT 25.265 154.745 30.610 155.290 ;
        RECT 31.245 154.745 31.535 155.470 ;
        RECT 33.290 155.290 33.630 156.120 ;
        RECT 35.110 155.610 35.460 156.860 ;
        RECT 38.810 155.290 39.150 156.120 ;
        RECT 40.630 155.610 40.980 156.860 ;
        RECT 42.745 156.205 44.415 157.295 ;
        RECT 42.745 155.515 43.495 156.035 ;
        RECT 43.665 155.685 44.415 156.205 ;
        RECT 44.595 156.155 44.925 157.295 ;
        RECT 45.455 156.325 45.785 157.110 ;
        RECT 45.105 156.155 45.785 156.325 ;
        RECT 46.025 156.155 46.235 157.295 ;
        RECT 44.585 155.735 44.935 155.985 ;
        RECT 45.105 155.555 45.275 156.155 ;
        RECT 46.405 156.145 46.735 157.125 ;
        RECT 46.905 156.155 47.135 157.295 ;
        RECT 47.345 156.155 47.730 157.125 ;
        RECT 47.900 156.835 48.225 157.295 ;
        RECT 48.745 156.665 49.025 157.125 ;
        RECT 47.900 156.445 49.025 156.665 ;
        RECT 45.445 155.735 45.795 155.985 ;
        RECT 31.705 154.745 37.050 155.290 ;
        RECT 37.225 154.745 42.570 155.290 ;
        RECT 42.745 154.745 44.415 155.515 ;
        RECT 44.595 154.745 44.865 155.555 ;
        RECT 45.035 154.915 45.365 155.555 ;
        RECT 45.535 154.745 45.775 155.555 ;
        RECT 46.025 154.745 46.235 155.565 ;
        RECT 46.405 155.545 46.655 156.145 ;
        RECT 46.825 155.735 47.155 155.985 ;
        RECT 46.405 154.915 46.735 155.545 ;
        RECT 46.905 154.745 47.135 155.565 ;
        RECT 47.345 155.485 47.625 156.155 ;
        RECT 47.900 155.985 48.350 156.445 ;
        RECT 49.215 156.275 49.615 157.125 ;
        RECT 50.015 156.835 50.285 157.295 ;
        RECT 50.455 156.665 50.740 157.125 ;
        RECT 51.950 156.915 52.285 157.295 ;
        RECT 47.795 155.655 48.350 155.985 ;
        RECT 48.520 155.715 49.615 156.275 ;
        RECT 47.900 155.545 48.350 155.655 ;
        RECT 47.345 154.915 47.730 155.485 ;
        RECT 47.900 155.375 49.025 155.545 ;
        RECT 47.900 154.745 48.225 155.205 ;
        RECT 48.745 154.915 49.025 155.375 ;
        RECT 49.215 154.915 49.615 155.715 ;
        RECT 49.785 156.445 50.740 156.665 ;
        RECT 49.785 155.545 49.995 156.445 ;
        RECT 50.165 155.715 50.855 156.275 ;
        RECT 49.785 155.375 50.740 155.545 ;
        RECT 51.945 155.425 52.185 156.735 ;
        RECT 52.455 156.325 52.705 157.125 ;
        RECT 52.925 156.575 53.255 157.295 ;
        RECT 53.440 156.325 53.690 157.125 ;
        RECT 54.155 156.495 54.485 157.295 ;
        RECT 54.655 156.865 54.995 157.125 ;
        RECT 52.355 156.155 54.545 156.325 ;
        RECT 50.015 154.745 50.285 155.205 ;
        RECT 50.455 154.915 50.740 155.375 ;
        RECT 52.355 155.245 52.525 156.155 ;
        RECT 54.230 155.985 54.545 156.155 ;
        RECT 52.030 154.915 52.525 155.245 ;
        RECT 52.745 155.020 53.095 155.985 ;
        RECT 53.275 155.015 53.575 155.985 ;
        RECT 53.755 155.015 54.035 155.985 ;
        RECT 54.230 155.735 54.560 155.985 ;
        RECT 54.215 154.745 54.485 155.545 ;
        RECT 54.735 155.465 54.995 156.865 ;
        RECT 55.165 156.205 56.835 157.295 ;
        RECT 54.655 154.955 54.995 155.465 ;
        RECT 55.165 155.515 55.915 156.035 ;
        RECT 56.085 155.685 56.835 156.205 ;
        RECT 57.005 156.130 57.295 157.295 ;
        RECT 57.475 156.155 57.805 157.295 ;
        RECT 58.335 156.325 58.665 157.110 ;
        RECT 58.935 156.625 59.105 157.125 ;
        RECT 59.275 156.795 59.605 157.295 ;
        RECT 58.935 156.455 59.600 156.625 ;
        RECT 57.985 156.155 58.665 156.325 ;
        RECT 57.465 155.735 57.815 155.985 ;
        RECT 57.985 155.555 58.155 156.155 ;
        RECT 58.325 155.735 58.675 155.985 ;
        RECT 58.850 155.635 59.200 156.285 ;
        RECT 55.165 154.745 56.835 155.515 ;
        RECT 57.005 154.745 57.295 155.470 ;
        RECT 57.475 154.745 57.745 155.555 ;
        RECT 57.915 154.915 58.245 155.555 ;
        RECT 58.415 154.745 58.655 155.555 ;
        RECT 59.370 155.465 59.600 156.455 ;
        RECT 58.935 155.295 59.600 155.465 ;
        RECT 58.935 155.005 59.105 155.295 ;
        RECT 59.275 154.745 59.605 155.125 ;
        RECT 59.775 155.005 59.960 157.125 ;
        RECT 60.200 156.835 60.465 157.295 ;
        RECT 60.635 156.700 60.885 157.125 ;
        RECT 61.095 156.850 62.200 157.020 ;
        RECT 60.580 156.570 60.885 156.700 ;
        RECT 60.130 155.375 60.410 156.325 ;
        RECT 60.580 155.465 60.750 156.570 ;
        RECT 60.920 155.785 61.160 156.380 ;
        RECT 61.330 156.315 61.860 156.680 ;
        RECT 61.330 155.615 61.500 156.315 ;
        RECT 62.030 156.235 62.200 156.850 ;
        RECT 62.370 156.495 62.540 157.295 ;
        RECT 62.710 156.795 62.960 157.125 ;
        RECT 63.185 156.825 64.070 156.995 ;
        RECT 62.030 156.145 62.540 156.235 ;
        RECT 60.580 155.335 60.805 155.465 ;
        RECT 60.975 155.395 61.500 155.615 ;
        RECT 61.670 155.975 62.540 156.145 ;
        RECT 60.215 154.745 60.465 155.205 ;
        RECT 60.635 155.195 60.805 155.335 ;
        RECT 61.670 155.195 61.840 155.975 ;
        RECT 62.370 155.905 62.540 155.975 ;
        RECT 62.050 155.725 62.250 155.755 ;
        RECT 62.710 155.725 62.880 156.795 ;
        RECT 63.050 155.905 63.240 156.625 ;
        RECT 62.050 155.425 62.880 155.725 ;
        RECT 63.410 155.695 63.730 156.655 ;
        RECT 60.635 155.025 60.970 155.195 ;
        RECT 61.165 155.025 61.840 155.195 ;
        RECT 62.160 154.745 62.530 155.245 ;
        RECT 62.710 155.195 62.880 155.425 ;
        RECT 63.265 155.365 63.730 155.695 ;
        RECT 63.900 155.985 64.070 156.825 ;
        RECT 64.250 156.795 64.565 157.295 ;
        RECT 64.795 156.565 65.135 157.125 ;
        RECT 64.240 156.190 65.135 156.565 ;
        RECT 65.305 156.285 65.475 157.295 ;
        RECT 64.945 155.985 65.135 156.190 ;
        RECT 65.645 156.235 65.975 157.080 ;
        RECT 65.645 156.155 66.035 156.235 ;
        RECT 65.820 156.105 66.035 156.155 ;
        RECT 63.900 155.655 64.775 155.985 ;
        RECT 64.945 155.655 65.695 155.985 ;
        RECT 63.900 155.195 64.070 155.655 ;
        RECT 64.945 155.485 65.145 155.655 ;
        RECT 65.865 155.525 66.035 156.105 ;
        RECT 65.810 155.485 66.035 155.525 ;
        RECT 62.710 155.025 63.115 155.195 ;
        RECT 63.285 155.025 64.070 155.195 ;
        RECT 64.345 154.745 64.555 155.275 ;
        RECT 64.815 154.960 65.145 155.485 ;
        RECT 65.655 155.400 66.035 155.485 ;
        RECT 66.205 156.155 66.590 157.115 ;
        RECT 66.805 156.495 67.095 157.295 ;
        RECT 67.265 156.955 68.630 157.125 ;
        RECT 67.265 156.325 67.435 156.955 ;
        RECT 66.760 156.155 67.435 156.325 ;
        RECT 66.205 156.105 66.435 156.155 ;
        RECT 66.205 155.485 66.380 156.105 ;
        RECT 66.760 155.985 66.930 156.155 ;
        RECT 67.605 155.985 67.930 156.785 ;
        RECT 68.300 156.745 68.630 156.955 ;
        RECT 68.300 156.495 69.255 156.745 ;
        RECT 66.565 155.735 66.930 155.985 ;
        RECT 67.125 155.735 67.375 155.985 ;
        RECT 66.565 155.655 66.755 155.735 ;
        RECT 67.125 155.655 67.295 155.735 ;
        RECT 67.585 155.655 67.930 155.985 ;
        RECT 68.100 155.655 68.375 156.320 ;
        RECT 68.560 155.655 68.915 156.320 ;
        RECT 69.085 155.485 69.255 156.495 ;
        RECT 69.425 156.155 69.715 157.295 ;
        RECT 70.000 156.665 70.285 157.125 ;
        RECT 70.455 156.835 70.725 157.295 ;
        RECT 70.000 156.445 70.955 156.665 ;
        RECT 69.440 155.655 69.715 155.985 ;
        RECT 69.885 155.715 70.575 156.275 ;
        RECT 70.745 155.545 70.955 156.445 ;
        RECT 65.315 154.745 65.485 155.355 ;
        RECT 65.655 154.965 65.985 155.400 ;
        RECT 66.205 154.915 66.715 155.485 ;
        RECT 67.260 155.315 68.660 155.485 ;
        RECT 66.885 154.745 67.055 155.305 ;
        RECT 67.260 154.915 67.590 155.315 ;
        RECT 67.765 154.745 68.095 155.145 ;
        RECT 68.330 155.125 68.660 155.315 ;
        RECT 68.830 155.295 69.255 155.485 ;
        RECT 69.425 155.125 69.715 155.395 ;
        RECT 68.330 154.915 69.715 155.125 ;
        RECT 70.000 155.375 70.955 155.545 ;
        RECT 71.125 156.275 71.525 157.125 ;
        RECT 71.715 156.665 71.995 157.125 ;
        RECT 72.515 156.835 72.840 157.295 ;
        RECT 71.715 156.445 72.840 156.665 ;
        RECT 71.125 155.715 72.220 156.275 ;
        RECT 72.390 155.985 72.840 156.445 ;
        RECT 73.010 156.155 73.395 157.125 ;
        RECT 70.000 154.915 70.285 155.375 ;
        RECT 70.455 154.745 70.725 155.205 ;
        RECT 71.125 154.915 71.525 155.715 ;
        RECT 72.390 155.655 72.945 155.985 ;
        RECT 72.390 155.545 72.840 155.655 ;
        RECT 71.715 155.375 72.840 155.545 ;
        RECT 73.115 155.485 73.395 156.155 ;
        RECT 71.715 154.915 71.995 155.375 ;
        RECT 72.515 154.745 72.840 155.205 ;
        RECT 73.010 154.915 73.395 155.485 ;
        RECT 73.565 156.155 73.950 157.115 ;
        RECT 74.165 156.495 74.455 157.295 ;
        RECT 74.625 156.955 75.990 157.125 ;
        RECT 74.625 156.325 74.795 156.955 ;
        RECT 74.120 156.155 74.795 156.325 ;
        RECT 73.565 155.485 73.740 156.155 ;
        RECT 74.120 155.985 74.290 156.155 ;
        RECT 74.965 155.985 75.290 156.785 ;
        RECT 75.660 156.745 75.990 156.955 ;
        RECT 75.660 156.495 76.615 156.745 ;
        RECT 73.925 155.735 74.290 155.985 ;
        RECT 74.485 155.735 74.735 155.985 ;
        RECT 73.925 155.655 74.115 155.735 ;
        RECT 74.485 155.655 74.655 155.735 ;
        RECT 74.945 155.655 75.290 155.985 ;
        RECT 75.460 155.655 75.735 156.320 ;
        RECT 75.920 155.655 76.275 156.320 ;
        RECT 76.445 155.485 76.615 156.495 ;
        RECT 76.785 156.155 77.075 157.295 ;
        RECT 77.360 156.665 77.645 157.125 ;
        RECT 77.815 156.835 78.085 157.295 ;
        RECT 77.360 156.445 78.315 156.665 ;
        RECT 76.800 155.655 77.075 155.985 ;
        RECT 77.245 155.715 77.935 156.275 ;
        RECT 78.105 155.545 78.315 156.445 ;
        RECT 73.565 154.915 74.075 155.485 ;
        RECT 74.620 155.315 76.020 155.485 ;
        RECT 74.245 154.745 74.415 155.305 ;
        RECT 74.620 154.915 74.950 155.315 ;
        RECT 75.125 154.745 75.455 155.145 ;
        RECT 75.690 155.125 76.020 155.315 ;
        RECT 76.190 155.295 76.615 155.485 ;
        RECT 76.785 155.125 77.075 155.395 ;
        RECT 75.690 154.915 77.075 155.125 ;
        RECT 77.360 155.375 78.315 155.545 ;
        RECT 78.485 156.275 78.885 157.125 ;
        RECT 79.075 156.665 79.355 157.125 ;
        RECT 79.875 156.835 80.200 157.295 ;
        RECT 79.075 156.445 80.200 156.665 ;
        RECT 78.485 155.715 79.580 156.275 ;
        RECT 79.750 155.985 80.200 156.445 ;
        RECT 80.370 156.155 80.755 157.125 ;
        RECT 80.935 156.685 81.265 157.115 ;
        RECT 81.445 156.855 81.640 157.295 ;
        RECT 81.810 156.685 82.140 157.115 ;
        RECT 80.935 156.515 82.140 156.685 ;
        RECT 80.935 156.185 81.830 156.515 ;
        RECT 82.310 156.345 82.585 157.115 ;
        RECT 77.360 154.915 77.645 155.375 ;
        RECT 77.815 154.745 78.085 155.205 ;
        RECT 78.485 154.915 78.885 155.715 ;
        RECT 79.750 155.655 80.305 155.985 ;
        RECT 79.750 155.545 80.200 155.655 ;
        RECT 79.075 155.375 80.200 155.545 ;
        RECT 80.475 155.485 80.755 156.155 ;
        RECT 82.000 156.155 82.585 156.345 ;
        RECT 80.940 155.655 81.235 155.985 ;
        RECT 81.415 155.655 81.830 155.985 ;
        RECT 79.075 154.915 79.355 155.375 ;
        RECT 79.875 154.745 80.200 155.205 ;
        RECT 80.370 154.915 80.755 155.485 ;
        RECT 80.935 154.745 81.235 155.475 ;
        RECT 81.415 155.035 81.645 155.655 ;
        RECT 82.000 155.485 82.175 156.155 ;
        RECT 82.765 156.130 83.055 157.295 ;
        RECT 83.265 156.155 83.495 157.295 ;
        RECT 83.665 156.145 83.995 157.125 ;
        RECT 84.165 156.155 84.375 157.295 ;
        RECT 84.605 156.860 89.950 157.295 ;
        RECT 81.845 155.305 82.175 155.485 ;
        RECT 82.345 155.335 82.585 155.985 ;
        RECT 83.245 155.735 83.575 155.985 ;
        RECT 81.845 154.925 82.070 155.305 ;
        RECT 82.240 154.745 82.570 155.135 ;
        RECT 82.765 154.745 83.055 155.470 ;
        RECT 83.265 154.745 83.495 155.565 ;
        RECT 83.745 155.545 83.995 156.145 ;
        RECT 83.665 154.915 83.995 155.545 ;
        RECT 84.165 154.745 84.375 155.565 ;
        RECT 86.190 155.290 86.530 156.120 ;
        RECT 88.010 155.610 88.360 156.860 ;
        RECT 91.045 156.205 92.255 157.295 ;
        RECT 91.045 155.665 91.565 156.205 ;
        RECT 91.735 155.495 92.255 156.035 ;
        RECT 84.605 154.745 89.950 155.290 ;
        RECT 91.045 154.745 92.255 155.495 ;
        RECT 18.280 154.575 92.340 154.745 ;
        RECT 18.365 153.825 19.575 154.575 ;
        RECT 19.745 154.030 25.090 154.575 ;
        RECT 25.265 154.030 30.610 154.575 ;
        RECT 30.785 154.030 36.130 154.575 ;
        RECT 36.305 154.030 41.650 154.575 ;
        RECT 41.850 154.185 42.180 154.575 ;
        RECT 18.365 153.285 18.885 153.825 ;
        RECT 19.055 153.115 19.575 153.655 ;
        RECT 21.330 153.200 21.670 154.030 ;
        RECT 18.365 152.025 19.575 153.115 ;
        RECT 23.150 152.460 23.500 153.710 ;
        RECT 26.850 153.200 27.190 154.030 ;
        RECT 28.670 152.460 29.020 153.710 ;
        RECT 32.370 153.200 32.710 154.030 ;
        RECT 34.190 152.460 34.540 153.710 ;
        RECT 37.890 153.200 38.230 154.030 ;
        RECT 42.350 154.015 42.575 154.395 ;
        RECT 39.710 152.460 40.060 153.710 ;
        RECT 41.835 153.335 42.075 153.985 ;
        RECT 42.245 153.835 42.575 154.015 ;
        RECT 42.245 153.165 42.420 153.835 ;
        RECT 42.775 153.665 43.005 154.285 ;
        RECT 43.185 153.845 43.485 154.575 ;
        RECT 44.125 153.850 44.415 154.575 ;
        RECT 44.585 153.805 46.255 154.575 ;
        RECT 46.425 153.835 46.935 154.405 ;
        RECT 47.105 154.015 47.275 154.575 ;
        RECT 47.480 154.005 47.810 154.405 ;
        RECT 47.985 154.175 48.315 154.575 ;
        RECT 48.550 154.195 49.935 154.405 ;
        RECT 48.550 154.005 48.880 154.195 ;
        RECT 47.480 153.835 48.880 154.005 ;
        RECT 49.050 153.835 49.475 154.025 ;
        RECT 49.645 153.925 49.935 154.195 ;
        RECT 42.590 153.335 43.005 153.665 ;
        RECT 43.185 153.335 43.480 153.665 ;
        RECT 44.585 153.285 45.335 153.805 ;
        RECT 41.835 152.975 42.420 153.165 ;
        RECT 19.745 152.025 25.090 152.460 ;
        RECT 25.265 152.025 30.610 152.460 ;
        RECT 30.785 152.025 36.130 152.460 ;
        RECT 36.305 152.025 41.650 152.460 ;
        RECT 41.835 152.205 42.110 152.975 ;
        RECT 42.590 152.805 43.485 153.135 ;
        RECT 42.280 152.635 43.485 152.805 ;
        RECT 42.280 152.205 42.610 152.635 ;
        RECT 42.780 152.025 42.975 152.465 ;
        RECT 43.155 152.205 43.485 152.635 ;
        RECT 44.125 152.025 44.415 153.190 ;
        RECT 45.505 153.115 46.255 153.635 ;
        RECT 44.585 152.025 46.255 153.115 ;
        RECT 46.425 153.165 46.600 153.835 ;
        RECT 46.785 153.585 46.975 153.665 ;
        RECT 47.345 153.585 47.515 153.665 ;
        RECT 46.785 153.335 47.150 153.585 ;
        RECT 47.345 153.335 47.595 153.585 ;
        RECT 47.805 153.335 48.150 153.665 ;
        RECT 46.980 153.165 47.150 153.335 ;
        RECT 46.425 152.205 46.810 153.165 ;
        RECT 46.980 152.995 47.655 153.165 ;
        RECT 47.025 152.025 47.315 152.825 ;
        RECT 47.485 152.365 47.655 152.995 ;
        RECT 47.825 152.535 48.150 153.335 ;
        RECT 48.320 153.000 48.595 153.665 ;
        RECT 48.780 153.000 49.135 153.665 ;
        RECT 49.305 152.825 49.475 153.835 ;
        RECT 50.105 153.900 50.380 154.245 ;
        RECT 50.570 154.175 50.945 154.575 ;
        RECT 51.115 154.005 51.285 154.355 ;
        RECT 51.455 154.175 51.785 154.575 ;
        RECT 51.955 154.005 52.215 154.405 ;
        RECT 49.660 153.335 49.935 153.665 ;
        RECT 50.105 153.165 50.275 153.900 ;
        RECT 50.550 153.835 52.215 154.005 ;
        RECT 50.550 153.665 50.720 153.835 ;
        RECT 52.395 153.755 52.725 154.175 ;
        RECT 52.895 153.755 53.155 154.575 ;
        RECT 53.325 153.855 53.665 154.365 ;
        RECT 52.395 153.665 52.645 153.755 ;
        RECT 50.445 153.335 50.720 153.665 ;
        RECT 50.890 153.335 51.715 153.665 ;
        RECT 51.930 153.335 52.645 153.665 ;
        RECT 52.815 153.335 53.150 153.585 ;
        RECT 50.550 153.165 50.720 153.335 ;
        RECT 48.520 152.575 49.475 152.825 ;
        RECT 48.520 152.365 48.850 152.575 ;
        RECT 47.485 152.195 48.850 152.365 ;
        RECT 49.645 152.025 49.935 153.165 ;
        RECT 50.105 152.195 50.380 153.165 ;
        RECT 50.550 152.995 51.210 153.165 ;
        RECT 51.470 153.045 51.715 153.335 ;
        RECT 51.040 152.875 51.210 152.995 ;
        RECT 51.885 152.875 52.215 153.165 ;
        RECT 50.590 152.025 50.870 152.825 ;
        RECT 51.040 152.705 52.215 152.875 ;
        RECT 52.475 152.775 52.645 153.335 ;
        RECT 51.040 152.205 52.655 152.535 ;
        RECT 52.895 152.025 53.155 153.165 ;
        RECT 53.325 152.455 53.585 153.855 ;
        RECT 53.835 153.775 54.105 154.575 ;
        RECT 53.760 153.335 54.090 153.585 ;
        RECT 54.285 153.335 54.565 154.305 ;
        RECT 54.745 153.335 55.045 154.305 ;
        RECT 55.225 153.335 55.575 154.300 ;
        RECT 55.795 154.075 56.290 154.405 ;
        RECT 56.545 154.115 57.105 154.405 ;
        RECT 57.275 154.115 57.525 154.575 ;
        RECT 53.775 153.165 54.090 153.335 ;
        RECT 55.795 153.165 55.965 154.075 ;
        RECT 53.775 152.995 55.965 153.165 ;
        RECT 53.325 152.195 53.665 152.455 ;
        RECT 53.835 152.025 54.165 152.825 ;
        RECT 54.630 152.195 54.880 152.995 ;
        RECT 55.065 152.025 55.395 152.745 ;
        RECT 55.615 152.195 55.865 152.995 ;
        RECT 56.135 152.585 56.375 153.895 ;
        RECT 56.545 152.745 56.795 154.115 ;
        RECT 58.145 153.945 58.475 154.305 ;
        RECT 58.845 154.030 64.190 154.575 ;
        RECT 57.085 153.755 58.475 153.945 ;
        RECT 57.085 153.665 57.255 153.755 ;
        RECT 56.965 153.335 57.255 153.665 ;
        RECT 57.425 153.335 57.765 153.585 ;
        RECT 57.985 153.335 58.660 153.585 ;
        RECT 57.085 153.085 57.255 153.335 ;
        RECT 57.085 152.915 58.025 153.085 ;
        RECT 58.395 152.975 58.660 153.335 ;
        RECT 60.430 153.200 60.770 154.030 ;
        RECT 64.365 153.805 66.035 154.575 ;
        RECT 56.035 152.025 56.370 152.405 ;
        RECT 56.545 152.195 57.005 152.745 ;
        RECT 57.195 152.025 57.525 152.745 ;
        RECT 57.725 152.365 58.025 152.915 ;
        RECT 58.195 152.025 58.475 152.695 ;
        RECT 62.250 152.460 62.600 153.710 ;
        RECT 64.365 153.285 65.115 153.805 ;
        RECT 66.215 153.765 66.485 154.575 ;
        RECT 66.655 153.765 66.985 154.405 ;
        RECT 67.155 153.765 67.395 154.575 ;
        RECT 67.585 153.925 67.845 154.405 ;
        RECT 68.015 154.035 68.265 154.575 ;
        RECT 65.285 153.115 66.035 153.635 ;
        RECT 66.205 153.335 66.555 153.585 ;
        RECT 66.725 153.165 66.895 153.765 ;
        RECT 67.065 153.335 67.415 153.585 ;
        RECT 58.845 152.025 64.190 152.460 ;
        RECT 64.365 152.025 66.035 153.115 ;
        RECT 66.215 152.025 66.545 153.165 ;
        RECT 66.725 152.995 67.405 153.165 ;
        RECT 67.075 152.210 67.405 152.995 ;
        RECT 67.585 152.895 67.755 153.925 ;
        RECT 68.435 153.870 68.655 154.355 ;
        RECT 67.925 153.275 68.155 153.670 ;
        RECT 68.325 153.445 68.655 153.870 ;
        RECT 68.825 154.195 69.715 154.365 ;
        RECT 68.825 153.470 68.995 154.195 ;
        RECT 69.165 153.640 69.715 154.025 ;
        RECT 69.885 153.850 70.175 154.575 ;
        RECT 70.435 154.075 70.930 154.405 ;
        RECT 68.825 153.400 69.715 153.470 ;
        RECT 68.820 153.375 69.715 153.400 ;
        RECT 68.810 153.360 69.715 153.375 ;
        RECT 68.805 153.345 69.715 153.360 ;
        RECT 68.795 153.340 69.715 153.345 ;
        RECT 68.790 153.330 69.715 153.340 ;
        RECT 68.785 153.320 69.715 153.330 ;
        RECT 68.775 153.315 69.715 153.320 ;
        RECT 68.765 153.305 69.715 153.315 ;
        RECT 68.755 153.300 69.715 153.305 ;
        RECT 68.755 153.295 69.090 153.300 ;
        RECT 68.740 153.290 69.090 153.295 ;
        RECT 68.725 153.280 69.090 153.290 ;
        RECT 68.700 153.275 69.090 153.280 ;
        RECT 67.925 153.270 69.090 153.275 ;
        RECT 67.925 153.235 69.060 153.270 ;
        RECT 67.925 153.210 69.025 153.235 ;
        RECT 67.925 153.180 68.995 153.210 ;
        RECT 67.925 153.150 68.975 153.180 ;
        RECT 67.925 153.120 68.955 153.150 ;
        RECT 67.925 153.110 68.885 153.120 ;
        RECT 67.925 153.100 68.860 153.110 ;
        RECT 67.925 153.085 68.840 153.100 ;
        RECT 67.925 153.070 68.820 153.085 ;
        RECT 68.030 153.060 68.815 153.070 ;
        RECT 68.030 153.025 68.800 153.060 ;
        RECT 67.585 152.195 67.860 152.895 ;
        RECT 68.030 152.775 68.785 153.025 ;
        RECT 68.955 152.705 69.285 152.950 ;
        RECT 69.455 152.850 69.715 153.300 ;
        RECT 69.100 152.680 69.285 152.705 ;
        RECT 69.100 152.580 69.715 152.680 ;
        RECT 68.030 152.025 68.285 152.570 ;
        RECT 68.455 152.195 68.935 152.535 ;
        RECT 69.110 152.025 69.715 152.580 ;
        RECT 69.885 152.025 70.175 153.190 ;
        RECT 70.385 152.585 70.590 153.905 ;
        RECT 70.760 153.165 70.930 154.075 ;
        RECT 71.150 153.335 71.505 154.240 ;
        RECT 71.680 153.355 71.980 154.245 ;
        RECT 71.680 153.335 71.850 153.355 ;
        RECT 72.160 153.335 72.420 154.245 ;
        RECT 72.590 153.770 72.825 154.575 ;
        RECT 72.995 154.320 73.325 154.365 ;
        RECT 72.995 153.855 73.330 154.320 ;
        RECT 72.590 153.345 72.985 153.585 ;
        RECT 72.590 153.165 72.815 153.345 ;
        RECT 73.155 153.165 73.330 153.855 ;
        RECT 73.515 153.850 73.845 154.575 ;
        RECT 74.065 153.755 74.295 154.575 ;
        RECT 74.465 153.775 74.795 154.405 ;
        RECT 74.045 153.335 74.375 153.585 ;
        RECT 74.545 153.175 74.795 153.775 ;
        RECT 74.965 153.755 75.175 154.575 ;
        RECT 75.495 154.025 75.665 154.315 ;
        RECT 75.835 154.195 76.165 154.575 ;
        RECT 75.495 153.855 76.160 154.025 ;
        RECT 70.760 152.995 72.815 153.165 ;
        RECT 70.355 152.025 70.685 152.405 ;
        RECT 70.860 152.195 71.110 152.995 ;
        RECT 71.330 152.025 71.660 152.745 ;
        RECT 71.845 152.195 72.095 152.995 ;
        RECT 72.995 152.875 73.330 153.165 ;
        RECT 72.495 152.025 72.825 152.825 ;
        RECT 72.995 152.705 73.335 152.875 ;
        RECT 72.995 152.195 73.330 152.705 ;
        RECT 73.505 152.025 73.835 152.825 ;
        RECT 74.065 152.025 74.295 153.165 ;
        RECT 74.465 152.195 74.795 153.175 ;
        RECT 74.965 152.025 75.175 153.165 ;
        RECT 75.410 153.035 75.760 153.685 ;
        RECT 75.930 152.865 76.160 153.855 ;
        RECT 75.495 152.695 76.160 152.865 ;
        RECT 75.495 152.195 75.665 152.695 ;
        RECT 75.835 152.025 76.165 152.525 ;
        RECT 76.335 152.195 76.520 154.315 ;
        RECT 76.775 154.115 77.025 154.575 ;
        RECT 77.195 154.125 77.530 154.295 ;
        RECT 77.725 154.125 78.400 154.295 ;
        RECT 77.195 153.985 77.365 154.125 ;
        RECT 76.690 152.995 76.970 153.945 ;
        RECT 77.140 153.855 77.365 153.985 ;
        RECT 77.140 152.750 77.310 153.855 ;
        RECT 77.535 153.705 78.060 153.925 ;
        RECT 77.480 152.940 77.720 153.535 ;
        RECT 77.890 153.005 78.060 153.705 ;
        RECT 78.230 153.345 78.400 154.125 ;
        RECT 78.720 154.075 79.090 154.575 ;
        RECT 79.270 154.125 79.675 154.295 ;
        RECT 79.845 154.125 80.630 154.295 ;
        RECT 79.270 153.895 79.440 154.125 ;
        RECT 78.610 153.595 79.440 153.895 ;
        RECT 79.825 153.625 80.290 153.955 ;
        RECT 78.610 153.565 78.810 153.595 ;
        RECT 78.930 153.345 79.100 153.415 ;
        RECT 78.230 153.175 79.100 153.345 ;
        RECT 78.590 153.085 79.100 153.175 ;
        RECT 77.140 152.620 77.445 152.750 ;
        RECT 77.890 152.640 78.420 153.005 ;
        RECT 76.760 152.025 77.025 152.485 ;
        RECT 77.195 152.195 77.445 152.620 ;
        RECT 78.590 152.470 78.760 153.085 ;
        RECT 77.655 152.300 78.760 152.470 ;
        RECT 78.930 152.025 79.100 152.825 ;
        RECT 79.270 152.525 79.440 153.595 ;
        RECT 79.610 152.695 79.800 153.415 ;
        RECT 79.970 152.665 80.290 153.625 ;
        RECT 80.460 153.665 80.630 154.125 ;
        RECT 80.905 154.045 81.115 154.575 ;
        RECT 81.375 153.835 81.705 154.360 ;
        RECT 81.875 153.965 82.045 154.575 ;
        RECT 82.215 153.920 82.545 154.355 ;
        RECT 82.765 154.030 88.110 154.575 ;
        RECT 82.215 153.835 82.595 153.920 ;
        RECT 81.505 153.665 81.705 153.835 ;
        RECT 82.370 153.795 82.595 153.835 ;
        RECT 80.460 153.335 81.335 153.665 ;
        RECT 81.505 153.335 82.255 153.665 ;
        RECT 79.270 152.195 79.520 152.525 ;
        RECT 80.460 152.495 80.630 153.335 ;
        RECT 81.505 153.130 81.695 153.335 ;
        RECT 82.425 153.215 82.595 153.795 ;
        RECT 82.380 153.165 82.595 153.215 ;
        RECT 84.350 153.200 84.690 154.030 ;
        RECT 88.285 153.805 90.875 154.575 ;
        RECT 91.045 153.825 92.255 154.575 ;
        RECT 80.800 152.755 81.695 153.130 ;
        RECT 82.205 153.085 82.595 153.165 ;
        RECT 79.745 152.325 80.630 152.495 ;
        RECT 80.810 152.025 81.125 152.525 ;
        RECT 81.355 152.195 81.695 152.755 ;
        RECT 81.865 152.025 82.035 153.035 ;
        RECT 82.205 152.240 82.535 153.085 ;
        RECT 86.170 152.460 86.520 153.710 ;
        RECT 88.285 153.285 89.495 153.805 ;
        RECT 89.665 153.115 90.875 153.635 ;
        RECT 82.765 152.025 88.110 152.460 ;
        RECT 88.285 152.025 90.875 153.115 ;
        RECT 91.045 153.115 91.565 153.655 ;
        RECT 91.735 153.285 92.255 153.825 ;
        RECT 91.045 152.025 92.255 153.115 ;
        RECT 18.280 151.855 92.340 152.025 ;
        RECT 18.365 150.765 19.575 151.855 ;
        RECT 19.745 151.420 25.090 151.855 ;
        RECT 25.265 151.420 30.610 151.855 ;
        RECT 18.365 150.055 18.885 150.595 ;
        RECT 19.055 150.225 19.575 150.765 ;
        RECT 18.365 149.305 19.575 150.055 ;
        RECT 21.330 149.850 21.670 150.680 ;
        RECT 23.150 150.170 23.500 151.420 ;
        RECT 26.850 149.850 27.190 150.680 ;
        RECT 28.670 150.170 29.020 151.420 ;
        RECT 31.245 150.690 31.535 151.855 ;
        RECT 31.705 150.765 35.215 151.855 ;
        RECT 35.385 150.765 36.595 151.855 ;
        RECT 36.855 151.185 37.025 151.685 ;
        RECT 37.195 151.355 37.525 151.855 ;
        RECT 36.855 151.015 37.520 151.185 ;
        RECT 31.705 150.075 33.355 150.595 ;
        RECT 33.525 150.245 35.215 150.765 ;
        RECT 19.745 149.305 25.090 149.850 ;
        RECT 25.265 149.305 30.610 149.850 ;
        RECT 31.245 149.305 31.535 150.030 ;
        RECT 31.705 149.305 35.215 150.075 ;
        RECT 35.385 150.055 35.905 150.595 ;
        RECT 36.075 150.225 36.595 150.765 ;
        RECT 36.770 150.195 37.120 150.845 ;
        RECT 35.385 149.305 36.595 150.055 ;
        RECT 37.290 150.025 37.520 151.015 ;
        RECT 36.855 149.855 37.520 150.025 ;
        RECT 36.855 149.565 37.025 149.855 ;
        RECT 37.195 149.305 37.525 149.685 ;
        RECT 37.695 149.565 37.880 151.685 ;
        RECT 38.120 151.395 38.385 151.855 ;
        RECT 38.555 151.260 38.805 151.685 ;
        RECT 39.015 151.410 40.120 151.580 ;
        RECT 38.500 151.130 38.805 151.260 ;
        RECT 38.050 149.935 38.330 150.885 ;
        RECT 38.500 150.025 38.670 151.130 ;
        RECT 38.840 150.345 39.080 150.940 ;
        RECT 39.250 150.875 39.780 151.240 ;
        RECT 39.250 150.175 39.420 150.875 ;
        RECT 39.950 150.795 40.120 151.410 ;
        RECT 40.290 151.055 40.460 151.855 ;
        RECT 40.630 151.355 40.880 151.685 ;
        RECT 41.105 151.385 41.990 151.555 ;
        RECT 39.950 150.705 40.460 150.795 ;
        RECT 38.500 149.895 38.725 150.025 ;
        RECT 38.895 149.955 39.420 150.175 ;
        RECT 39.590 150.535 40.460 150.705 ;
        RECT 38.135 149.305 38.385 149.765 ;
        RECT 38.555 149.755 38.725 149.895 ;
        RECT 39.590 149.755 39.760 150.535 ;
        RECT 40.290 150.465 40.460 150.535 ;
        RECT 39.970 150.285 40.170 150.315 ;
        RECT 40.630 150.285 40.800 151.355 ;
        RECT 40.970 150.465 41.160 151.185 ;
        RECT 39.970 149.985 40.800 150.285 ;
        RECT 41.330 150.255 41.650 151.215 ;
        RECT 38.555 149.585 38.890 149.755 ;
        RECT 39.085 149.585 39.760 149.755 ;
        RECT 40.080 149.305 40.450 149.805 ;
        RECT 40.630 149.755 40.800 149.985 ;
        RECT 41.185 149.925 41.650 150.255 ;
        RECT 41.820 150.545 41.990 151.385 ;
        RECT 42.170 151.355 42.485 151.855 ;
        RECT 42.715 151.125 43.055 151.685 ;
        RECT 42.160 150.750 43.055 151.125 ;
        RECT 43.225 150.845 43.395 151.855 ;
        RECT 42.865 150.545 43.055 150.750 ;
        RECT 43.565 150.795 43.895 151.640 ;
        RECT 44.700 151.225 44.985 151.685 ;
        RECT 45.155 151.395 45.425 151.855 ;
        RECT 44.700 151.005 45.655 151.225 ;
        RECT 43.565 150.715 43.955 150.795 ;
        RECT 43.740 150.665 43.955 150.715 ;
        RECT 41.820 150.215 42.695 150.545 ;
        RECT 42.865 150.215 43.615 150.545 ;
        RECT 41.820 149.755 41.990 150.215 ;
        RECT 42.865 150.045 43.065 150.215 ;
        RECT 43.785 150.085 43.955 150.665 ;
        RECT 44.585 150.275 45.275 150.835 ;
        RECT 45.445 150.105 45.655 151.005 ;
        RECT 43.730 150.045 43.955 150.085 ;
        RECT 40.630 149.585 41.035 149.755 ;
        RECT 41.205 149.585 41.990 149.755 ;
        RECT 42.265 149.305 42.475 149.835 ;
        RECT 42.735 149.520 43.065 150.045 ;
        RECT 43.575 149.960 43.955 150.045 ;
        RECT 43.235 149.305 43.405 149.915 ;
        RECT 43.575 149.525 43.905 149.960 ;
        RECT 44.700 149.935 45.655 150.105 ;
        RECT 45.825 150.835 46.225 151.685 ;
        RECT 46.415 151.225 46.695 151.685 ;
        RECT 47.215 151.395 47.540 151.855 ;
        RECT 46.415 151.005 47.540 151.225 ;
        RECT 45.825 150.275 46.920 150.835 ;
        RECT 47.090 150.545 47.540 151.005 ;
        RECT 47.710 150.715 48.095 151.685 ;
        RECT 48.265 150.715 48.545 151.855 ;
        RECT 44.700 149.475 44.985 149.935 ;
        RECT 45.155 149.305 45.425 149.765 ;
        RECT 45.825 149.475 46.225 150.275 ;
        RECT 47.090 150.215 47.645 150.545 ;
        RECT 47.090 150.105 47.540 150.215 ;
        RECT 46.415 149.935 47.540 150.105 ;
        RECT 47.815 150.045 48.095 150.715 ;
        RECT 48.715 150.705 49.045 151.685 ;
        RECT 49.215 150.715 49.475 151.855 ;
        RECT 50.115 150.795 50.445 151.645 ;
        RECT 48.275 150.275 48.610 150.545 ;
        RECT 48.780 150.105 48.950 150.705 ;
        RECT 49.120 150.295 49.455 150.545 ;
        RECT 46.415 149.475 46.695 149.935 ;
        RECT 47.215 149.305 47.540 149.765 ;
        RECT 47.710 149.475 48.095 150.045 ;
        RECT 48.265 149.305 48.575 150.105 ;
        RECT 48.780 149.475 49.475 150.105 ;
        RECT 50.115 150.030 50.305 150.795 ;
        RECT 50.615 150.715 50.865 151.855 ;
        RECT 51.055 151.215 51.305 151.635 ;
        RECT 51.535 151.385 51.865 151.855 ;
        RECT 52.095 151.215 52.345 151.635 ;
        RECT 51.055 151.045 52.345 151.215 ;
        RECT 52.525 151.215 52.855 151.645 ;
        RECT 52.525 151.045 52.980 151.215 ;
        RECT 51.045 150.545 51.260 150.875 ;
        RECT 50.475 150.215 50.785 150.545 ;
        RECT 50.955 150.215 51.260 150.545 ;
        RECT 51.435 150.215 51.720 150.875 ;
        RECT 51.915 150.215 52.180 150.875 ;
        RECT 52.395 150.215 52.640 150.875 ;
        RECT 50.615 150.045 50.785 150.215 ;
        RECT 52.810 150.045 52.980 151.045 ;
        RECT 53.325 150.765 56.835 151.855 ;
        RECT 50.115 149.520 50.445 150.030 ;
        RECT 50.615 149.875 52.980 150.045 ;
        RECT 53.325 150.075 54.975 150.595 ;
        RECT 55.145 150.245 56.835 150.765 ;
        RECT 57.005 150.690 57.295 151.855 ;
        RECT 57.465 150.765 60.055 151.855 ;
        RECT 57.465 150.075 58.675 150.595 ;
        RECT 58.845 150.245 60.055 150.765 ;
        RECT 60.235 150.905 60.510 151.675 ;
        RECT 60.680 151.245 61.010 151.675 ;
        RECT 61.180 151.415 61.375 151.855 ;
        RECT 61.555 151.245 61.885 151.675 ;
        RECT 60.680 151.075 61.885 151.245 ;
        RECT 60.235 150.715 60.820 150.905 ;
        RECT 60.990 150.745 61.885 151.075 ;
        RECT 62.075 150.715 62.405 151.855 ;
        RECT 62.935 150.885 63.265 151.670 ;
        RECT 63.445 151.420 68.790 151.855 ;
        RECT 62.585 150.715 63.265 150.885 ;
        RECT 50.615 149.305 50.945 149.705 ;
        RECT 51.995 149.535 52.325 149.875 ;
        RECT 52.495 149.305 52.825 149.705 ;
        RECT 53.325 149.305 56.835 150.075 ;
        RECT 57.005 149.305 57.295 150.030 ;
        RECT 57.465 149.305 60.055 150.075 ;
        RECT 60.235 149.895 60.475 150.545 ;
        RECT 60.645 150.045 60.820 150.715 ;
        RECT 60.990 150.215 61.405 150.545 ;
        RECT 61.585 150.215 61.880 150.545 ;
        RECT 62.065 150.295 62.415 150.545 ;
        RECT 60.645 149.865 60.975 150.045 ;
        RECT 60.250 149.305 60.580 149.695 ;
        RECT 60.750 149.485 60.975 149.865 ;
        RECT 61.175 149.595 61.405 150.215 ;
        RECT 62.585 150.115 62.755 150.715 ;
        RECT 62.925 150.295 63.275 150.545 ;
        RECT 61.585 149.305 61.885 150.035 ;
        RECT 62.075 149.305 62.345 150.115 ;
        RECT 62.515 149.475 62.845 150.115 ;
        RECT 63.015 149.305 63.255 150.115 ;
        RECT 65.030 149.850 65.370 150.680 ;
        RECT 66.850 150.170 67.200 151.420 ;
        RECT 69.425 151.345 69.725 151.855 ;
        RECT 69.895 151.175 70.225 151.685 ;
        RECT 70.395 151.345 71.025 151.855 ;
        RECT 71.605 151.345 71.985 151.515 ;
        RECT 72.155 151.345 72.455 151.855 ;
        RECT 71.815 151.175 71.985 151.345 ;
        RECT 69.425 151.005 71.645 151.175 ;
        RECT 69.425 150.045 69.595 151.005 ;
        RECT 69.765 150.665 71.305 150.835 ;
        RECT 69.765 150.215 70.010 150.665 ;
        RECT 70.270 150.295 70.965 150.495 ;
        RECT 71.135 150.465 71.305 150.665 ;
        RECT 71.475 150.805 71.645 151.005 ;
        RECT 71.815 150.975 72.475 151.175 ;
        RECT 71.475 150.635 72.135 150.805 ;
        RECT 71.135 150.295 71.735 150.465 ;
        RECT 71.965 150.215 72.135 150.635 ;
        RECT 63.445 149.305 68.790 149.850 ;
        RECT 69.425 149.500 69.890 150.045 ;
        RECT 70.395 149.305 70.565 150.125 ;
        RECT 70.735 150.045 71.645 150.125 ;
        RECT 72.305 150.045 72.475 150.975 ;
        RECT 72.645 150.765 73.855 151.855 ;
        RECT 70.735 149.955 71.985 150.045 ;
        RECT 70.735 149.475 71.065 149.955 ;
        RECT 71.475 149.875 71.985 149.955 ;
        RECT 71.235 149.305 71.585 149.695 ;
        RECT 71.755 149.475 71.985 149.875 ;
        RECT 72.155 149.565 72.475 150.045 ;
        RECT 72.645 150.055 73.165 150.595 ;
        RECT 73.335 150.225 73.855 150.765 ;
        RECT 74.035 150.885 74.365 151.670 ;
        RECT 74.035 150.715 74.715 150.885 ;
        RECT 74.895 150.715 75.225 151.855 ;
        RECT 75.405 151.420 80.750 151.855 ;
        RECT 74.025 150.295 74.375 150.545 ;
        RECT 74.545 150.115 74.715 150.715 ;
        RECT 74.885 150.295 75.235 150.545 ;
        RECT 72.645 149.305 73.855 150.055 ;
        RECT 74.045 149.305 74.285 150.115 ;
        RECT 74.455 149.475 74.785 150.115 ;
        RECT 74.955 149.305 75.225 150.115 ;
        RECT 76.990 149.850 77.330 150.680 ;
        RECT 78.810 150.170 79.160 151.420 ;
        RECT 80.925 150.765 82.595 151.855 ;
        RECT 80.925 150.075 81.675 150.595 ;
        RECT 81.845 150.245 82.595 150.765 ;
        RECT 82.765 150.690 83.055 151.855 ;
        RECT 83.225 151.420 88.570 151.855 ;
        RECT 75.405 149.305 80.750 149.850 ;
        RECT 80.925 149.305 82.595 150.075 ;
        RECT 82.765 149.305 83.055 150.030 ;
        RECT 84.810 149.850 85.150 150.680 ;
        RECT 86.630 150.170 86.980 151.420 ;
        RECT 88.745 150.765 90.415 151.855 ;
        RECT 88.745 150.075 89.495 150.595 ;
        RECT 89.665 150.245 90.415 150.765 ;
        RECT 91.045 150.765 92.255 151.855 ;
        RECT 91.045 150.225 91.565 150.765 ;
        RECT 83.225 149.305 88.570 149.850 ;
        RECT 88.745 149.305 90.415 150.075 ;
        RECT 91.735 150.055 92.255 150.595 ;
        RECT 91.045 149.305 92.255 150.055 ;
        RECT 18.280 149.135 92.340 149.305 ;
        RECT 18.365 148.385 19.575 149.135 ;
        RECT 19.745 148.590 25.090 149.135 ;
        RECT 25.265 148.590 30.610 149.135 ;
        RECT 30.785 148.590 36.130 149.135 ;
        RECT 36.305 148.590 41.650 149.135 ;
        RECT 18.365 147.845 18.885 148.385 ;
        RECT 19.055 147.675 19.575 148.215 ;
        RECT 21.330 147.760 21.670 148.590 ;
        RECT 18.365 146.585 19.575 147.675 ;
        RECT 23.150 147.020 23.500 148.270 ;
        RECT 26.850 147.760 27.190 148.590 ;
        RECT 28.670 147.020 29.020 148.270 ;
        RECT 32.370 147.760 32.710 148.590 ;
        RECT 34.190 147.020 34.540 148.270 ;
        RECT 37.890 147.760 38.230 148.590 ;
        RECT 41.825 148.365 43.495 149.135 ;
        RECT 44.125 148.410 44.415 149.135 ;
        RECT 44.585 148.590 49.930 149.135 ;
        RECT 39.710 147.020 40.060 148.270 ;
        RECT 41.825 147.845 42.575 148.365 ;
        RECT 42.745 147.675 43.495 148.195 ;
        RECT 46.170 147.760 46.510 148.590 ;
        RECT 50.105 148.365 53.615 149.135 ;
        RECT 19.745 146.585 25.090 147.020 ;
        RECT 25.265 146.585 30.610 147.020 ;
        RECT 30.785 146.585 36.130 147.020 ;
        RECT 36.305 146.585 41.650 147.020 ;
        RECT 41.825 146.585 43.495 147.675 ;
        RECT 44.125 146.585 44.415 147.750 ;
        RECT 47.990 147.020 48.340 148.270 ;
        RECT 50.105 147.845 51.755 148.365 ;
        RECT 53.785 148.335 54.095 149.135 ;
        RECT 54.300 148.335 54.995 148.965 ;
        RECT 55.625 148.335 56.320 148.965 ;
        RECT 56.525 148.335 56.835 149.135 ;
        RECT 57.005 148.395 57.390 148.965 ;
        RECT 57.560 148.675 57.885 149.135 ;
        RECT 58.405 148.505 58.685 148.965 ;
        RECT 54.300 148.285 54.475 148.335 ;
        RECT 51.925 147.675 53.615 148.195 ;
        RECT 53.795 147.895 54.130 148.165 ;
        RECT 54.300 147.735 54.470 148.285 ;
        RECT 54.640 147.895 54.975 148.145 ;
        RECT 55.645 147.895 55.980 148.145 ;
        RECT 56.150 147.735 56.320 148.335 ;
        RECT 56.490 147.895 56.825 148.165 ;
        RECT 44.585 146.585 49.930 147.020 ;
        RECT 50.105 146.585 53.615 147.675 ;
        RECT 53.785 146.585 54.065 147.725 ;
        RECT 54.235 146.755 54.565 147.735 ;
        RECT 54.735 146.585 54.995 147.725 ;
        RECT 55.625 146.585 55.885 147.725 ;
        RECT 56.055 146.755 56.385 147.735 ;
        RECT 57.005 147.725 57.285 148.395 ;
        RECT 57.560 148.335 58.685 148.505 ;
        RECT 57.560 148.225 58.010 148.335 ;
        RECT 57.455 147.895 58.010 148.225 ;
        RECT 58.875 148.165 59.275 148.965 ;
        RECT 59.675 148.675 59.945 149.135 ;
        RECT 60.115 148.505 60.400 148.965 ;
        RECT 56.555 146.585 56.835 147.725 ;
        RECT 57.005 146.755 57.390 147.725 ;
        RECT 57.560 147.435 58.010 147.895 ;
        RECT 58.180 147.605 59.275 148.165 ;
        RECT 57.560 147.215 58.685 147.435 ;
        RECT 57.560 146.585 57.885 147.045 ;
        RECT 58.405 146.755 58.685 147.215 ;
        RECT 58.875 146.755 59.275 147.605 ;
        RECT 59.445 148.335 60.400 148.505 ;
        RECT 59.445 147.435 59.655 148.335 ;
        RECT 60.685 148.315 60.945 149.135 ;
        RECT 61.115 148.315 61.445 148.735 ;
        RECT 61.625 148.565 61.885 148.965 ;
        RECT 62.055 148.735 62.385 149.135 ;
        RECT 62.555 148.565 62.725 148.915 ;
        RECT 62.895 148.735 63.270 149.135 ;
        RECT 61.625 148.395 63.290 148.565 ;
        RECT 63.460 148.460 63.735 148.805 ;
        RECT 63.965 148.655 64.245 149.135 ;
        RECT 64.415 148.485 64.675 148.875 ;
        RECT 64.850 148.655 65.105 149.135 ;
        RECT 65.275 148.485 65.570 148.875 ;
        RECT 65.750 148.655 66.025 149.135 ;
        RECT 66.195 148.635 66.495 148.965 ;
        RECT 61.195 148.225 61.445 148.315 ;
        RECT 63.120 148.225 63.290 148.395 ;
        RECT 59.825 147.605 60.515 148.165 ;
        RECT 60.690 147.895 61.025 148.145 ;
        RECT 61.195 147.895 61.910 148.225 ;
        RECT 62.125 147.895 62.950 148.225 ;
        RECT 63.120 147.895 63.395 148.225 ;
        RECT 59.445 147.215 60.400 147.435 ;
        RECT 59.675 146.585 59.945 147.045 ;
        RECT 60.115 146.755 60.400 147.215 ;
        RECT 60.685 146.585 60.945 147.725 ;
        RECT 61.195 147.335 61.365 147.895 ;
        RECT 61.625 147.435 61.955 147.725 ;
        RECT 62.125 147.605 62.370 147.895 ;
        RECT 63.120 147.725 63.290 147.895 ;
        RECT 63.565 147.725 63.735 148.460 ;
        RECT 62.630 147.555 63.290 147.725 ;
        RECT 62.630 147.435 62.800 147.555 ;
        RECT 61.625 147.265 62.800 147.435 ;
        RECT 61.185 146.765 62.800 147.095 ;
        RECT 62.970 146.585 63.250 147.385 ;
        RECT 63.460 146.755 63.735 147.725 ;
        RECT 63.920 148.315 65.570 148.485 ;
        RECT 63.920 147.805 64.325 148.315 ;
        RECT 64.495 147.975 65.635 148.145 ;
        RECT 63.920 147.635 64.675 147.805 ;
        RECT 63.960 146.585 64.245 147.455 ;
        RECT 64.415 147.385 64.675 147.635 ;
        RECT 65.465 147.725 65.635 147.975 ;
        RECT 65.805 147.895 66.155 148.465 ;
        RECT 66.325 147.725 66.495 148.635 ;
        RECT 66.665 148.365 69.255 149.135 ;
        RECT 69.885 148.410 70.175 149.135 ;
        RECT 70.345 148.395 70.685 148.965 ;
        RECT 70.880 148.470 71.050 149.135 ;
        RECT 71.330 148.795 71.550 148.840 ;
        RECT 71.325 148.625 71.550 148.795 ;
        RECT 71.720 148.655 72.165 148.825 ;
        RECT 71.330 148.485 71.550 148.625 ;
        RECT 66.665 147.845 67.875 148.365 ;
        RECT 65.465 147.555 66.495 147.725 ;
        RECT 68.045 147.675 69.255 148.195 ;
        RECT 64.415 147.215 65.535 147.385 ;
        RECT 64.415 146.755 64.675 147.215 ;
        RECT 64.850 146.585 65.105 147.045 ;
        RECT 65.275 146.755 65.535 147.215 ;
        RECT 65.705 146.585 66.015 147.385 ;
        RECT 66.185 146.755 66.495 147.555 ;
        RECT 66.665 146.585 69.255 147.675 ;
        RECT 69.885 146.585 70.175 147.750 ;
        RECT 70.345 147.425 70.520 148.395 ;
        RECT 71.330 148.315 71.825 148.485 ;
        RECT 70.690 147.775 70.860 148.225 ;
        RECT 71.030 147.945 71.480 148.145 ;
        RECT 71.650 148.120 71.825 148.315 ;
        RECT 71.995 147.865 72.165 148.655 ;
        RECT 72.335 148.530 72.585 148.900 ;
        RECT 72.415 148.145 72.585 148.530 ;
        RECT 72.755 148.495 73.005 148.900 ;
        RECT 73.175 148.665 73.345 149.135 ;
        RECT 73.515 148.495 73.855 148.900 ;
        RECT 74.025 148.590 79.370 149.135 ;
        RECT 79.545 148.590 84.890 149.135 ;
        RECT 85.065 148.590 90.410 149.135 ;
        RECT 72.755 148.315 73.855 148.495 ;
        RECT 72.415 147.975 72.610 148.145 ;
        RECT 70.690 147.605 71.085 147.775 ;
        RECT 71.995 147.725 72.270 147.865 ;
        RECT 70.345 146.755 70.605 147.425 ;
        RECT 70.915 147.335 71.085 147.605 ;
        RECT 71.255 147.505 72.270 147.725 ;
        RECT 72.440 147.725 72.610 147.975 ;
        RECT 72.780 147.895 73.340 148.145 ;
        RECT 72.440 147.335 72.995 147.725 ;
        RECT 70.915 147.165 72.995 147.335 ;
        RECT 70.775 146.585 71.105 146.985 ;
        RECT 71.975 146.585 72.375 146.985 ;
        RECT 72.665 146.930 72.995 147.165 ;
        RECT 73.165 146.795 73.340 147.895 ;
        RECT 73.510 147.575 73.855 148.145 ;
        RECT 75.610 147.760 75.950 148.590 ;
        RECT 73.510 146.585 73.855 147.405 ;
        RECT 77.430 147.020 77.780 148.270 ;
        RECT 81.130 147.760 81.470 148.590 ;
        RECT 82.950 147.020 83.300 148.270 ;
        RECT 86.650 147.760 86.990 148.590 ;
        RECT 91.045 148.385 92.255 149.135 ;
        RECT 88.470 147.020 88.820 148.270 ;
        RECT 91.045 147.675 91.565 148.215 ;
        RECT 91.735 147.845 92.255 148.385 ;
        RECT 74.025 146.585 79.370 147.020 ;
        RECT 79.545 146.585 84.890 147.020 ;
        RECT 85.065 146.585 90.410 147.020 ;
        RECT 91.045 146.585 92.255 147.675 ;
        RECT 18.280 146.415 92.340 146.585 ;
        RECT 18.365 145.325 19.575 146.415 ;
        RECT 19.745 145.980 25.090 146.415 ;
        RECT 25.265 145.980 30.610 146.415 ;
        RECT 18.365 144.615 18.885 145.155 ;
        RECT 19.055 144.785 19.575 145.325 ;
        RECT 18.365 143.865 19.575 144.615 ;
        RECT 21.330 144.410 21.670 145.240 ;
        RECT 23.150 144.730 23.500 145.980 ;
        RECT 26.850 144.410 27.190 145.240 ;
        RECT 28.670 144.730 29.020 145.980 ;
        RECT 31.245 145.250 31.535 146.415 ;
        RECT 31.705 145.980 37.050 146.415 ;
        RECT 37.225 145.980 42.570 146.415 ;
        RECT 19.745 143.865 25.090 144.410 ;
        RECT 25.265 143.865 30.610 144.410 ;
        RECT 31.245 143.865 31.535 144.590 ;
        RECT 33.290 144.410 33.630 145.240 ;
        RECT 35.110 144.730 35.460 145.980 ;
        RECT 38.810 144.410 39.150 145.240 ;
        RECT 40.630 144.730 40.980 145.980 ;
        RECT 42.835 145.745 43.005 146.245 ;
        RECT 43.175 145.915 43.505 146.415 ;
        RECT 42.835 145.575 43.500 145.745 ;
        RECT 42.750 144.755 43.100 145.405 ;
        RECT 43.270 144.585 43.500 145.575 ;
        RECT 42.835 144.415 43.500 144.585 ;
        RECT 31.705 143.865 37.050 144.410 ;
        RECT 37.225 143.865 42.570 144.410 ;
        RECT 42.835 144.125 43.005 144.415 ;
        RECT 43.175 143.865 43.505 144.245 ;
        RECT 43.675 144.125 43.860 146.245 ;
        RECT 44.100 145.955 44.365 146.415 ;
        RECT 44.535 145.820 44.785 146.245 ;
        RECT 44.995 145.970 46.100 146.140 ;
        RECT 44.480 145.690 44.785 145.820 ;
        RECT 44.030 144.495 44.310 145.445 ;
        RECT 44.480 144.585 44.650 145.690 ;
        RECT 44.820 144.905 45.060 145.500 ;
        RECT 45.230 145.435 45.760 145.800 ;
        RECT 45.230 144.735 45.400 145.435 ;
        RECT 45.930 145.355 46.100 145.970 ;
        RECT 46.270 145.615 46.440 146.415 ;
        RECT 46.610 145.915 46.860 146.245 ;
        RECT 47.085 145.945 47.970 146.115 ;
        RECT 45.930 145.265 46.440 145.355 ;
        RECT 44.480 144.455 44.705 144.585 ;
        RECT 44.875 144.515 45.400 144.735 ;
        RECT 45.570 145.095 46.440 145.265 ;
        RECT 44.115 143.865 44.365 144.325 ;
        RECT 44.535 144.315 44.705 144.455 ;
        RECT 45.570 144.315 45.740 145.095 ;
        RECT 46.270 145.025 46.440 145.095 ;
        RECT 45.950 144.845 46.150 144.875 ;
        RECT 46.610 144.845 46.780 145.915 ;
        RECT 46.950 145.025 47.140 145.745 ;
        RECT 45.950 144.545 46.780 144.845 ;
        RECT 47.310 144.815 47.630 145.775 ;
        RECT 44.535 144.145 44.870 144.315 ;
        RECT 45.065 144.145 45.740 144.315 ;
        RECT 46.060 143.865 46.430 144.365 ;
        RECT 46.610 144.315 46.780 144.545 ;
        RECT 47.165 144.485 47.630 144.815 ;
        RECT 47.800 145.105 47.970 145.945 ;
        RECT 48.150 145.915 48.465 146.415 ;
        RECT 48.695 145.685 49.035 146.245 ;
        RECT 48.140 145.310 49.035 145.685 ;
        RECT 49.205 145.405 49.375 146.415 ;
        RECT 48.845 145.105 49.035 145.310 ;
        RECT 49.545 145.355 49.875 146.200 ;
        RECT 50.105 145.575 50.365 146.245 ;
        RECT 50.535 146.015 50.865 146.415 ;
        RECT 51.735 146.015 52.135 146.415 ;
        RECT 52.425 145.835 52.755 146.070 ;
        RECT 50.675 145.665 52.755 145.835 ;
        RECT 49.545 145.275 49.935 145.355 ;
        RECT 49.720 145.225 49.935 145.275 ;
        RECT 47.800 144.775 48.675 145.105 ;
        RECT 48.845 144.775 49.595 145.105 ;
        RECT 47.800 144.315 47.970 144.775 ;
        RECT 48.845 144.605 49.045 144.775 ;
        RECT 49.765 144.645 49.935 145.225 ;
        RECT 49.710 144.605 49.935 144.645 ;
        RECT 46.610 144.145 47.015 144.315 ;
        RECT 47.185 144.145 47.970 144.315 ;
        RECT 48.245 143.865 48.455 144.395 ;
        RECT 48.715 144.080 49.045 144.605 ;
        RECT 49.555 144.520 49.935 144.605 ;
        RECT 50.105 144.605 50.280 145.575 ;
        RECT 50.675 145.395 50.845 145.665 ;
        RECT 50.450 145.225 50.845 145.395 ;
        RECT 51.015 145.275 52.030 145.495 ;
        RECT 50.450 144.775 50.620 145.225 ;
        RECT 51.755 145.135 52.030 145.275 ;
        RECT 52.200 145.275 52.755 145.665 ;
        RECT 50.790 144.855 51.240 145.055 ;
        RECT 51.410 144.685 51.585 144.880 ;
        RECT 49.215 143.865 49.385 144.475 ;
        RECT 49.555 144.085 49.885 144.520 ;
        RECT 50.105 144.035 50.445 144.605 ;
        RECT 50.640 143.865 50.810 144.530 ;
        RECT 51.090 144.515 51.585 144.685 ;
        RECT 51.090 144.375 51.310 144.515 ;
        RECT 51.085 144.205 51.310 144.375 ;
        RECT 51.755 144.345 51.925 145.135 ;
        RECT 52.200 145.025 52.370 145.275 ;
        RECT 52.925 145.105 53.100 146.205 ;
        RECT 53.270 145.595 53.615 146.415 ;
        RECT 52.175 144.855 52.370 145.025 ;
        RECT 52.540 144.855 53.100 145.105 ;
        RECT 53.270 144.855 53.615 145.425 ;
        RECT 53.785 145.315 54.105 146.245 ;
        RECT 54.285 145.735 54.685 146.245 ;
        RECT 54.855 145.905 55.025 146.415 ;
        RECT 55.195 145.735 55.525 146.245 ;
        RECT 54.285 145.565 55.525 145.735 ;
        RECT 55.695 145.565 55.865 146.415 ;
        RECT 56.455 145.565 56.835 146.245 ;
        RECT 53.785 145.145 54.415 145.315 ;
        RECT 52.175 144.470 52.345 144.855 ;
        RECT 51.090 144.160 51.310 144.205 ;
        RECT 51.480 144.175 51.925 144.345 ;
        RECT 52.095 144.100 52.345 144.470 ;
        RECT 52.515 144.505 53.615 144.685 ;
        RECT 52.515 144.100 52.765 144.505 ;
        RECT 52.935 143.865 53.105 144.335 ;
        RECT 53.275 144.100 53.615 144.505 ;
        RECT 53.785 143.865 54.075 144.700 ;
        RECT 54.245 144.265 54.415 145.145 ;
        RECT 55.190 145.225 56.495 145.395 ;
        RECT 54.585 144.605 54.815 145.105 ;
        RECT 55.190 145.025 55.360 145.225 ;
        RECT 54.985 144.855 55.360 145.025 ;
        RECT 55.530 144.855 56.080 145.055 ;
        RECT 56.250 144.775 56.495 145.225 ;
        RECT 56.665 144.605 56.835 145.565 ;
        RECT 57.005 145.250 57.295 146.415 ;
        RECT 57.525 145.355 57.855 146.200 ;
        RECT 58.025 145.405 58.195 146.415 ;
        RECT 58.365 145.685 58.705 146.245 ;
        RECT 58.935 145.915 59.250 146.415 ;
        RECT 59.430 145.945 60.315 146.115 ;
        RECT 57.465 145.275 57.855 145.355 ;
        RECT 58.365 145.310 59.260 145.685 ;
        RECT 54.585 144.435 56.835 144.605 ;
        RECT 57.465 145.225 57.680 145.275 ;
        RECT 57.465 144.645 57.635 145.225 ;
        RECT 58.365 145.105 58.555 145.310 ;
        RECT 59.430 145.105 59.600 145.945 ;
        RECT 60.540 145.915 60.790 146.245 ;
        RECT 57.805 144.775 58.555 145.105 ;
        RECT 58.725 144.775 59.600 145.105 ;
        RECT 57.465 144.605 57.690 144.645 ;
        RECT 58.355 144.605 58.555 144.775 ;
        RECT 54.245 144.095 55.200 144.265 ;
        RECT 55.615 143.865 55.945 144.255 ;
        RECT 56.115 144.115 56.285 144.435 ;
        RECT 56.455 143.865 56.785 144.255 ;
        RECT 57.005 143.865 57.295 144.590 ;
        RECT 57.465 144.520 57.845 144.605 ;
        RECT 57.515 144.085 57.845 144.520 ;
        RECT 58.015 143.865 58.185 144.475 ;
        RECT 58.355 144.080 58.685 144.605 ;
        RECT 58.945 143.865 59.155 144.395 ;
        RECT 59.430 144.315 59.600 144.775 ;
        RECT 59.770 144.815 60.090 145.775 ;
        RECT 60.260 145.025 60.450 145.745 ;
        RECT 60.620 144.845 60.790 145.915 ;
        RECT 60.960 145.615 61.130 146.415 ;
        RECT 61.300 145.970 62.405 146.140 ;
        RECT 61.300 145.355 61.470 145.970 ;
        RECT 62.615 145.820 62.865 146.245 ;
        RECT 63.035 145.955 63.300 146.415 ;
        RECT 61.640 145.435 62.170 145.800 ;
        RECT 62.615 145.690 62.920 145.820 ;
        RECT 60.960 145.265 61.470 145.355 ;
        RECT 60.960 145.095 61.830 145.265 ;
        RECT 60.960 145.025 61.130 145.095 ;
        RECT 61.250 144.845 61.450 144.875 ;
        RECT 59.770 144.485 60.235 144.815 ;
        RECT 60.620 144.545 61.450 144.845 ;
        RECT 60.620 144.315 60.790 144.545 ;
        RECT 59.430 144.145 60.215 144.315 ;
        RECT 60.385 144.145 60.790 144.315 ;
        RECT 60.970 143.865 61.340 144.365 ;
        RECT 61.660 144.315 61.830 145.095 ;
        RECT 62.000 144.735 62.170 145.435 ;
        RECT 62.340 144.905 62.580 145.500 ;
        RECT 62.000 144.515 62.525 144.735 ;
        RECT 62.750 144.585 62.920 145.690 ;
        RECT 62.695 144.455 62.920 144.585 ;
        RECT 63.090 144.495 63.370 145.445 ;
        RECT 62.695 144.315 62.865 144.455 ;
        RECT 61.660 144.145 62.335 144.315 ;
        RECT 62.530 144.145 62.865 144.315 ;
        RECT 63.035 143.865 63.285 144.325 ;
        RECT 63.540 144.125 63.725 146.245 ;
        RECT 63.895 145.915 64.225 146.415 ;
        RECT 64.395 145.745 64.565 146.245 ;
        RECT 63.900 145.575 64.565 145.745 ;
        RECT 65.375 145.745 65.545 146.245 ;
        RECT 65.715 145.915 66.045 146.415 ;
        RECT 65.375 145.575 66.040 145.745 ;
        RECT 63.900 144.585 64.130 145.575 ;
        RECT 64.300 144.755 64.650 145.405 ;
        RECT 65.290 144.755 65.640 145.405 ;
        RECT 65.810 144.585 66.040 145.575 ;
        RECT 63.900 144.415 64.565 144.585 ;
        RECT 63.895 143.865 64.225 144.245 ;
        RECT 64.395 144.125 64.565 144.415 ;
        RECT 65.375 144.415 66.040 144.585 ;
        RECT 65.375 144.125 65.545 144.415 ;
        RECT 65.715 143.865 66.045 144.245 ;
        RECT 66.215 144.125 66.400 146.245 ;
        RECT 66.640 145.955 66.905 146.415 ;
        RECT 67.075 145.820 67.325 146.245 ;
        RECT 67.535 145.970 68.640 146.140 ;
        RECT 67.020 145.690 67.325 145.820 ;
        RECT 66.570 144.495 66.850 145.445 ;
        RECT 67.020 144.585 67.190 145.690 ;
        RECT 67.360 144.905 67.600 145.500 ;
        RECT 67.770 145.435 68.300 145.800 ;
        RECT 67.770 144.735 67.940 145.435 ;
        RECT 68.470 145.355 68.640 145.970 ;
        RECT 68.810 145.615 68.980 146.415 ;
        RECT 69.150 145.915 69.400 146.245 ;
        RECT 69.625 145.945 70.510 146.115 ;
        RECT 68.470 145.265 68.980 145.355 ;
        RECT 67.020 144.455 67.245 144.585 ;
        RECT 67.415 144.515 67.940 144.735 ;
        RECT 68.110 145.095 68.980 145.265 ;
        RECT 66.655 143.865 66.905 144.325 ;
        RECT 67.075 144.315 67.245 144.455 ;
        RECT 68.110 144.315 68.280 145.095 ;
        RECT 68.810 145.025 68.980 145.095 ;
        RECT 68.490 144.845 68.690 144.875 ;
        RECT 69.150 144.845 69.320 145.915 ;
        RECT 69.490 145.025 69.680 145.745 ;
        RECT 68.490 144.545 69.320 144.845 ;
        RECT 69.850 144.815 70.170 145.775 ;
        RECT 67.075 144.145 67.410 144.315 ;
        RECT 67.605 144.145 68.280 144.315 ;
        RECT 68.600 143.865 68.970 144.365 ;
        RECT 69.150 144.315 69.320 144.545 ;
        RECT 69.705 144.485 70.170 144.815 ;
        RECT 70.340 145.105 70.510 145.945 ;
        RECT 70.690 145.915 71.005 146.415 ;
        RECT 71.235 145.685 71.575 146.245 ;
        RECT 70.680 145.310 71.575 145.685 ;
        RECT 71.745 145.405 71.915 146.415 ;
        RECT 71.385 145.105 71.575 145.310 ;
        RECT 72.085 145.355 72.415 146.200 ;
        RECT 72.645 145.980 77.990 146.415 ;
        RECT 72.085 145.275 72.475 145.355 ;
        RECT 72.260 145.225 72.475 145.275 ;
        RECT 70.340 144.775 71.215 145.105 ;
        RECT 71.385 144.775 72.135 145.105 ;
        RECT 70.340 144.315 70.510 144.775 ;
        RECT 71.385 144.605 71.585 144.775 ;
        RECT 72.305 144.645 72.475 145.225 ;
        RECT 72.250 144.605 72.475 144.645 ;
        RECT 69.150 144.145 69.555 144.315 ;
        RECT 69.725 144.145 70.510 144.315 ;
        RECT 70.785 143.865 70.995 144.395 ;
        RECT 71.255 144.080 71.585 144.605 ;
        RECT 72.095 144.520 72.475 144.605 ;
        RECT 71.755 143.865 71.925 144.475 ;
        RECT 72.095 144.085 72.425 144.520 ;
        RECT 74.230 144.410 74.570 145.240 ;
        RECT 76.050 144.730 76.400 145.980 ;
        RECT 78.165 145.325 81.675 146.415 ;
        RECT 78.165 144.635 79.815 145.155 ;
        RECT 79.985 144.805 81.675 145.325 ;
        RECT 82.765 145.250 83.055 146.415 ;
        RECT 83.225 145.980 88.570 146.415 ;
        RECT 72.645 143.865 77.990 144.410 ;
        RECT 78.165 143.865 81.675 144.635 ;
        RECT 82.765 143.865 83.055 144.590 ;
        RECT 84.810 144.410 85.150 145.240 ;
        RECT 86.630 144.730 86.980 145.980 ;
        RECT 88.745 145.325 90.415 146.415 ;
        RECT 88.745 144.635 89.495 145.155 ;
        RECT 89.665 144.805 90.415 145.325 ;
        RECT 91.045 145.325 92.255 146.415 ;
        RECT 91.045 144.785 91.565 145.325 ;
        RECT 83.225 143.865 88.570 144.410 ;
        RECT 88.745 143.865 90.415 144.635 ;
        RECT 91.735 144.615 92.255 145.155 ;
        RECT 91.045 143.865 92.255 144.615 ;
        RECT 18.280 143.695 92.340 143.865 ;
        RECT 18.365 142.945 19.575 143.695 ;
        RECT 19.745 143.150 25.090 143.695 ;
        RECT 25.265 143.150 30.610 143.695 ;
        RECT 30.785 143.150 36.130 143.695 ;
        RECT 36.305 143.150 41.650 143.695 ;
        RECT 18.365 142.405 18.885 142.945 ;
        RECT 19.055 142.235 19.575 142.775 ;
        RECT 21.330 142.320 21.670 143.150 ;
        RECT 18.365 141.145 19.575 142.235 ;
        RECT 23.150 141.580 23.500 142.830 ;
        RECT 26.850 142.320 27.190 143.150 ;
        RECT 28.670 141.580 29.020 142.830 ;
        RECT 32.370 142.320 32.710 143.150 ;
        RECT 34.190 141.580 34.540 142.830 ;
        RECT 37.890 142.320 38.230 143.150 ;
        RECT 41.825 142.925 43.495 143.695 ;
        RECT 44.125 142.970 44.415 143.695 ;
        RECT 39.710 141.580 40.060 142.830 ;
        RECT 41.825 142.405 42.575 142.925 ;
        RECT 44.595 142.885 44.865 143.695 ;
        RECT 45.035 142.885 45.365 143.525 ;
        RECT 45.535 142.885 45.775 143.695 ;
        RECT 45.965 143.150 51.310 143.695 ;
        RECT 51.485 143.150 56.830 143.695 ;
        RECT 57.005 143.150 62.350 143.695 ;
        RECT 42.745 142.235 43.495 142.755 ;
        RECT 44.585 142.455 44.935 142.705 ;
        RECT 19.745 141.145 25.090 141.580 ;
        RECT 25.265 141.145 30.610 141.580 ;
        RECT 30.785 141.145 36.130 141.580 ;
        RECT 36.305 141.145 41.650 141.580 ;
        RECT 41.825 141.145 43.495 142.235 ;
        RECT 44.125 141.145 44.415 142.310 ;
        RECT 45.105 142.285 45.275 142.885 ;
        RECT 45.445 142.455 45.795 142.705 ;
        RECT 47.550 142.320 47.890 143.150 ;
        RECT 44.595 141.145 44.925 142.285 ;
        RECT 45.105 142.115 45.785 142.285 ;
        RECT 45.455 141.330 45.785 142.115 ;
        RECT 49.370 141.580 49.720 142.830 ;
        RECT 53.070 142.320 53.410 143.150 ;
        RECT 54.890 141.580 55.240 142.830 ;
        RECT 58.590 142.320 58.930 143.150 ;
        RECT 62.525 142.925 66.035 143.695 ;
        RECT 60.410 141.580 60.760 142.830 ;
        RECT 62.525 142.405 64.175 142.925 ;
        RECT 66.675 142.885 66.945 143.695 ;
        RECT 67.115 142.885 67.445 143.525 ;
        RECT 67.615 142.885 67.855 143.695 ;
        RECT 68.045 142.925 69.715 143.695 ;
        RECT 69.885 142.970 70.175 143.695 ;
        RECT 70.345 143.150 75.690 143.695 ;
        RECT 75.865 143.150 81.210 143.695 ;
        RECT 81.385 143.150 86.730 143.695 ;
        RECT 64.345 142.235 66.035 142.755 ;
        RECT 66.665 142.455 67.015 142.705 ;
        RECT 67.185 142.285 67.355 142.885 ;
        RECT 67.525 142.455 67.875 142.705 ;
        RECT 68.045 142.405 68.795 142.925 ;
        RECT 45.965 141.145 51.310 141.580 ;
        RECT 51.485 141.145 56.830 141.580 ;
        RECT 57.005 141.145 62.350 141.580 ;
        RECT 62.525 141.145 66.035 142.235 ;
        RECT 66.675 141.145 67.005 142.285 ;
        RECT 67.185 142.115 67.865 142.285 ;
        RECT 68.965 142.235 69.715 142.755 ;
        RECT 71.930 142.320 72.270 143.150 ;
        RECT 67.535 141.330 67.865 142.115 ;
        RECT 68.045 141.145 69.715 142.235 ;
        RECT 69.885 141.145 70.175 142.310 ;
        RECT 73.750 141.580 74.100 142.830 ;
        RECT 77.450 142.320 77.790 143.150 ;
        RECT 79.270 141.580 79.620 142.830 ;
        RECT 82.970 142.320 83.310 143.150 ;
        RECT 86.905 142.925 90.415 143.695 ;
        RECT 91.045 142.945 92.255 143.695 ;
        RECT 84.790 141.580 85.140 142.830 ;
        RECT 86.905 142.405 88.555 142.925 ;
        RECT 88.725 142.235 90.415 142.755 ;
        RECT 70.345 141.145 75.690 141.580 ;
        RECT 75.865 141.145 81.210 141.580 ;
        RECT 81.385 141.145 86.730 141.580 ;
        RECT 86.905 141.145 90.415 142.235 ;
        RECT 91.045 142.235 91.565 142.775 ;
        RECT 91.735 142.405 92.255 142.945 ;
        RECT 91.045 141.145 92.255 142.235 ;
        RECT 110.180 141.630 111.830 141.800 ;
        RECT 18.280 140.975 92.340 141.145 ;
        RECT 18.365 139.885 19.575 140.975 ;
        RECT 19.745 140.540 25.090 140.975 ;
        RECT 25.265 140.540 30.610 140.975 ;
        RECT 18.365 139.175 18.885 139.715 ;
        RECT 19.055 139.345 19.575 139.885 ;
        RECT 18.365 138.425 19.575 139.175 ;
        RECT 21.330 138.970 21.670 139.800 ;
        RECT 23.150 139.290 23.500 140.540 ;
        RECT 26.850 138.970 27.190 139.800 ;
        RECT 28.670 139.290 29.020 140.540 ;
        RECT 31.245 139.810 31.535 140.975 ;
        RECT 31.705 140.540 37.050 140.975 ;
        RECT 37.225 140.540 42.570 140.975 ;
        RECT 42.745 140.540 48.090 140.975 ;
        RECT 48.265 140.540 53.610 140.975 ;
        RECT 19.745 138.425 25.090 138.970 ;
        RECT 25.265 138.425 30.610 138.970 ;
        RECT 31.245 138.425 31.535 139.150 ;
        RECT 33.290 138.970 33.630 139.800 ;
        RECT 35.110 139.290 35.460 140.540 ;
        RECT 38.810 138.970 39.150 139.800 ;
        RECT 40.630 139.290 40.980 140.540 ;
        RECT 44.330 138.970 44.670 139.800 ;
        RECT 46.150 139.290 46.500 140.540 ;
        RECT 49.850 138.970 50.190 139.800 ;
        RECT 51.670 139.290 52.020 140.540 ;
        RECT 53.785 139.885 56.375 140.975 ;
        RECT 53.785 139.195 54.995 139.715 ;
        RECT 55.165 139.365 56.375 139.885 ;
        RECT 57.005 139.810 57.295 140.975 ;
        RECT 57.465 140.540 62.810 140.975 ;
        RECT 62.985 140.540 68.330 140.975 ;
        RECT 68.505 140.540 73.850 140.975 ;
        RECT 74.025 140.540 79.370 140.975 ;
        RECT 31.705 138.425 37.050 138.970 ;
        RECT 37.225 138.425 42.570 138.970 ;
        RECT 42.745 138.425 48.090 138.970 ;
        RECT 48.265 138.425 53.610 138.970 ;
        RECT 53.785 138.425 56.375 139.195 ;
        RECT 57.005 138.425 57.295 139.150 ;
        RECT 59.050 138.970 59.390 139.800 ;
        RECT 60.870 139.290 61.220 140.540 ;
        RECT 64.570 138.970 64.910 139.800 ;
        RECT 66.390 139.290 66.740 140.540 ;
        RECT 70.090 138.970 70.430 139.800 ;
        RECT 71.910 139.290 72.260 140.540 ;
        RECT 75.610 138.970 75.950 139.800 ;
        RECT 77.430 139.290 77.780 140.540 ;
        RECT 79.545 139.885 82.135 140.975 ;
        RECT 79.545 139.195 80.755 139.715 ;
        RECT 80.925 139.365 82.135 139.885 ;
        RECT 82.765 139.810 83.055 140.975 ;
        RECT 83.225 140.540 88.570 140.975 ;
        RECT 57.465 138.425 62.810 138.970 ;
        RECT 62.985 138.425 68.330 138.970 ;
        RECT 68.505 138.425 73.850 138.970 ;
        RECT 74.025 138.425 79.370 138.970 ;
        RECT 79.545 138.425 82.135 139.195 ;
        RECT 82.765 138.425 83.055 139.150 ;
        RECT 84.810 138.970 85.150 139.800 ;
        RECT 86.630 139.290 86.980 140.540 ;
        RECT 88.745 139.885 90.415 140.975 ;
        RECT 88.745 139.195 89.495 139.715 ;
        RECT 89.665 139.365 90.415 139.885 ;
        RECT 91.045 139.885 92.255 140.975 ;
        RECT 91.045 139.345 91.565 139.885 ;
        RECT 83.225 138.425 88.570 138.970 ;
        RECT 88.745 138.425 90.415 139.195 ;
        RECT 91.735 139.175 92.255 139.715 ;
        RECT 91.045 138.425 92.255 139.175 ;
        RECT 18.280 138.255 92.340 138.425 ;
        RECT 18.365 137.505 19.575 138.255 ;
        RECT 19.745 137.710 25.090 138.255 ;
        RECT 25.265 137.710 30.610 138.255 ;
        RECT 30.785 137.710 36.130 138.255 ;
        RECT 36.305 137.710 41.650 138.255 ;
        RECT 18.365 136.965 18.885 137.505 ;
        RECT 19.055 136.795 19.575 137.335 ;
        RECT 21.330 136.880 21.670 137.710 ;
        RECT 18.365 135.705 19.575 136.795 ;
        RECT 23.150 136.140 23.500 137.390 ;
        RECT 26.850 136.880 27.190 137.710 ;
        RECT 28.670 136.140 29.020 137.390 ;
        RECT 32.370 136.880 32.710 137.710 ;
        RECT 34.190 136.140 34.540 137.390 ;
        RECT 37.890 136.880 38.230 137.710 ;
        RECT 41.825 137.485 43.495 138.255 ;
        RECT 44.125 137.530 44.415 138.255 ;
        RECT 44.585 137.710 49.930 138.255 ;
        RECT 50.105 137.710 55.450 138.255 ;
        RECT 55.625 137.710 60.970 138.255 ;
        RECT 61.145 137.710 66.490 138.255 ;
        RECT 39.710 136.140 40.060 137.390 ;
        RECT 41.825 136.965 42.575 137.485 ;
        RECT 42.745 136.795 43.495 137.315 ;
        RECT 46.170 136.880 46.510 137.710 ;
        RECT 19.745 135.705 25.090 136.140 ;
        RECT 25.265 135.705 30.610 136.140 ;
        RECT 30.785 135.705 36.130 136.140 ;
        RECT 36.305 135.705 41.650 136.140 ;
        RECT 41.825 135.705 43.495 136.795 ;
        RECT 44.125 135.705 44.415 136.870 ;
        RECT 47.990 136.140 48.340 137.390 ;
        RECT 51.690 136.880 52.030 137.710 ;
        RECT 53.510 136.140 53.860 137.390 ;
        RECT 57.210 136.880 57.550 137.710 ;
        RECT 59.030 136.140 59.380 137.390 ;
        RECT 62.730 136.880 63.070 137.710 ;
        RECT 66.665 137.485 69.255 138.255 ;
        RECT 69.885 137.530 70.175 138.255 ;
        RECT 70.345 137.710 75.690 138.255 ;
        RECT 75.865 137.710 81.210 138.255 ;
        RECT 81.385 137.710 86.730 138.255 ;
        RECT 64.550 136.140 64.900 137.390 ;
        RECT 66.665 136.965 67.875 137.485 ;
        RECT 68.045 136.795 69.255 137.315 ;
        RECT 71.930 136.880 72.270 137.710 ;
        RECT 44.585 135.705 49.930 136.140 ;
        RECT 50.105 135.705 55.450 136.140 ;
        RECT 55.625 135.705 60.970 136.140 ;
        RECT 61.145 135.705 66.490 136.140 ;
        RECT 66.665 135.705 69.255 136.795 ;
        RECT 69.885 135.705 70.175 136.870 ;
        RECT 73.750 136.140 74.100 137.390 ;
        RECT 77.450 136.880 77.790 137.710 ;
        RECT 79.270 136.140 79.620 137.390 ;
        RECT 82.970 136.880 83.310 137.710 ;
        RECT 86.905 137.485 90.415 138.255 ;
        RECT 91.045 137.505 92.255 138.255 ;
        RECT 84.790 136.140 85.140 137.390 ;
        RECT 86.905 136.965 88.555 137.485 ;
        RECT 88.725 136.795 90.415 137.315 ;
        RECT 70.345 135.705 75.690 136.140 ;
        RECT 75.865 135.705 81.210 136.140 ;
        RECT 81.385 135.705 86.730 136.140 ;
        RECT 86.905 135.705 90.415 136.795 ;
        RECT 91.045 136.795 91.565 137.335 ;
        RECT 91.735 136.965 92.255 137.505 ;
        RECT 91.045 135.705 92.255 136.795 ;
        RECT 18.280 135.535 92.340 135.705 ;
        RECT 18.365 134.445 19.575 135.535 ;
        RECT 19.745 135.100 25.090 135.535 ;
        RECT 25.265 135.100 30.610 135.535 ;
        RECT 18.365 133.735 18.885 134.275 ;
        RECT 19.055 133.905 19.575 134.445 ;
        RECT 18.365 132.985 19.575 133.735 ;
        RECT 21.330 133.530 21.670 134.360 ;
        RECT 23.150 133.850 23.500 135.100 ;
        RECT 26.850 133.530 27.190 134.360 ;
        RECT 28.670 133.850 29.020 135.100 ;
        RECT 31.245 134.370 31.535 135.535 ;
        RECT 31.705 135.100 37.050 135.535 ;
        RECT 37.225 135.100 42.570 135.535 ;
        RECT 19.745 132.985 25.090 133.530 ;
        RECT 25.265 132.985 30.610 133.530 ;
        RECT 31.245 132.985 31.535 133.710 ;
        RECT 33.290 133.530 33.630 134.360 ;
        RECT 35.110 133.850 35.460 135.100 ;
        RECT 38.810 133.530 39.150 134.360 ;
        RECT 40.630 133.850 40.980 135.100 ;
        RECT 42.745 134.445 43.955 135.535 ;
        RECT 42.745 133.735 43.265 134.275 ;
        RECT 43.435 133.905 43.955 134.445 ;
        RECT 44.125 134.370 44.415 135.535 ;
        RECT 44.585 135.100 49.930 135.535 ;
        RECT 50.105 135.100 55.450 135.535 ;
        RECT 31.705 132.985 37.050 133.530 ;
        RECT 37.225 132.985 42.570 133.530 ;
        RECT 42.745 132.985 43.955 133.735 ;
        RECT 44.125 132.985 44.415 133.710 ;
        RECT 46.170 133.530 46.510 134.360 ;
        RECT 47.990 133.850 48.340 135.100 ;
        RECT 51.690 133.530 52.030 134.360 ;
        RECT 53.510 133.850 53.860 135.100 ;
        RECT 55.625 134.445 56.835 135.535 ;
        RECT 55.625 133.735 56.145 134.275 ;
        RECT 56.315 133.905 56.835 134.445 ;
        RECT 57.005 134.370 57.295 135.535 ;
        RECT 57.465 135.100 62.810 135.535 ;
        RECT 62.985 135.100 68.330 135.535 ;
        RECT 44.585 132.985 49.930 133.530 ;
        RECT 50.105 132.985 55.450 133.530 ;
        RECT 55.625 132.985 56.835 133.735 ;
        RECT 57.005 132.985 57.295 133.710 ;
        RECT 59.050 133.530 59.390 134.360 ;
        RECT 60.870 133.850 61.220 135.100 ;
        RECT 64.570 133.530 64.910 134.360 ;
        RECT 66.390 133.850 66.740 135.100 ;
        RECT 68.505 134.445 69.715 135.535 ;
        RECT 68.505 133.735 69.025 134.275 ;
        RECT 69.195 133.905 69.715 134.445 ;
        RECT 69.885 134.370 70.175 135.535 ;
        RECT 70.345 135.100 75.690 135.535 ;
        RECT 75.865 135.100 81.210 135.535 ;
        RECT 57.465 132.985 62.810 133.530 ;
        RECT 62.985 132.985 68.330 133.530 ;
        RECT 68.505 132.985 69.715 133.735 ;
        RECT 69.885 132.985 70.175 133.710 ;
        RECT 71.930 133.530 72.270 134.360 ;
        RECT 73.750 133.850 74.100 135.100 ;
        RECT 77.450 133.530 77.790 134.360 ;
        RECT 79.270 133.850 79.620 135.100 ;
        RECT 81.385 134.445 82.595 135.535 ;
        RECT 81.385 133.735 81.905 134.275 ;
        RECT 82.075 133.905 82.595 134.445 ;
        RECT 82.765 134.370 83.055 135.535 ;
        RECT 83.225 135.100 88.570 135.535 ;
        RECT 70.345 132.985 75.690 133.530 ;
        RECT 75.865 132.985 81.210 133.530 ;
        RECT 81.385 132.985 82.595 133.735 ;
        RECT 82.765 132.985 83.055 133.710 ;
        RECT 84.810 133.530 85.150 134.360 ;
        RECT 86.630 133.850 86.980 135.100 ;
        RECT 88.745 134.445 90.415 135.535 ;
        RECT 88.745 133.755 89.495 134.275 ;
        RECT 89.665 133.925 90.415 134.445 ;
        RECT 91.045 134.445 92.255 135.535 ;
        RECT 91.045 133.905 91.565 134.445 ;
        RECT 83.225 132.985 88.570 133.530 ;
        RECT 88.745 132.985 90.415 133.755 ;
        RECT 91.735 133.735 92.255 134.275 ;
        RECT 91.045 132.985 92.255 133.735 ;
        RECT 18.280 132.815 92.340 132.985 ;
        RECT 106.180 114.630 107.830 114.800 ;
        RECT 106.180 69.350 106.350 114.630 ;
        RECT 106.830 111.990 107.180 114.150 ;
        RECT 106.830 69.830 107.180 71.990 ;
        RECT 107.660 69.350 107.830 114.630 ;
        RECT 110.180 96.350 110.350 141.630 ;
        RECT 110.830 138.990 111.180 141.150 ;
        RECT 110.830 96.830 111.180 98.990 ;
        RECT 111.660 96.350 111.830 141.630 ;
        RECT 110.180 96.180 111.830 96.350 ;
        RECT 113.180 141.630 114.830 141.800 ;
        RECT 113.180 96.350 113.350 141.630 ;
        RECT 113.830 138.990 114.180 141.150 ;
        RECT 113.830 96.830 114.180 98.990 ;
        RECT 114.660 96.350 114.830 141.630 ;
        RECT 113.180 96.180 114.830 96.350 ;
        RECT 116.180 141.630 117.830 141.800 ;
        RECT 116.180 96.350 116.350 141.630 ;
        RECT 116.830 138.990 117.180 141.150 ;
        RECT 116.830 96.830 117.180 98.990 ;
        RECT 117.660 96.350 117.830 141.630 ;
        RECT 116.180 96.180 117.830 96.350 ;
        RECT 119.180 141.630 120.830 141.800 ;
        RECT 119.180 96.350 119.350 141.630 ;
        RECT 119.830 138.990 120.180 141.150 ;
        RECT 119.830 96.830 120.180 98.990 ;
        RECT 120.660 96.350 120.830 141.630 ;
        RECT 119.180 96.180 120.830 96.350 ;
        RECT 122.180 141.630 123.830 141.800 ;
        RECT 122.180 96.350 122.350 141.630 ;
        RECT 122.830 138.990 123.180 141.150 ;
        RECT 122.830 96.830 123.180 98.990 ;
        RECT 123.660 96.350 123.830 141.630 ;
        RECT 122.180 96.180 123.830 96.350 ;
        RECT 125.180 141.630 126.830 141.800 ;
        RECT 125.180 96.350 125.350 141.630 ;
        RECT 125.830 138.990 126.180 141.150 ;
        RECT 125.830 96.830 126.180 98.990 ;
        RECT 126.660 96.350 126.830 141.630 ;
        RECT 125.180 96.180 126.830 96.350 ;
        RECT 128.180 141.630 129.830 141.800 ;
        RECT 128.180 96.350 128.350 141.630 ;
        RECT 128.830 138.990 129.180 141.150 ;
        RECT 128.830 96.830 129.180 98.990 ;
        RECT 129.660 96.350 129.830 141.630 ;
        RECT 128.180 96.180 129.830 96.350 ;
        RECT 131.180 141.630 132.830 141.800 ;
        RECT 131.180 96.350 131.350 141.630 ;
        RECT 131.830 138.990 132.180 141.150 ;
        RECT 131.830 96.830 132.180 98.990 ;
        RECT 132.660 96.350 132.830 141.630 ;
        RECT 131.180 96.180 132.830 96.350 ;
        RECT 106.180 69.180 107.830 69.350 ;
        RECT 110.180 94.630 111.830 94.800 ;
        RECT 110.180 69.350 110.350 94.630 ;
        RECT 110.830 91.990 111.180 94.150 ;
        RECT 110.830 69.830 111.180 71.990 ;
        RECT 111.660 69.350 111.830 94.630 ;
        RECT 110.180 69.180 111.830 69.350 ;
        RECT 113.180 94.630 114.830 94.800 ;
        RECT 113.180 69.350 113.350 94.630 ;
        RECT 113.830 91.990 114.180 94.150 ;
        RECT 113.830 69.830 114.180 71.990 ;
        RECT 114.660 69.350 114.830 94.630 ;
        RECT 113.180 69.180 114.830 69.350 ;
        RECT 116.180 94.630 117.830 94.800 ;
        RECT 116.180 69.350 116.350 94.630 ;
        RECT 116.830 91.990 117.180 94.150 ;
        RECT 116.830 69.830 117.180 71.990 ;
        RECT 117.660 69.350 117.830 94.630 ;
        RECT 116.180 69.180 117.830 69.350 ;
        RECT 119.180 94.630 120.830 94.800 ;
        RECT 119.180 69.350 119.350 94.630 ;
        RECT 119.830 91.990 120.180 94.150 ;
        RECT 119.830 69.830 120.180 71.990 ;
        RECT 120.660 69.350 120.830 94.630 ;
        RECT 119.180 69.180 120.830 69.350 ;
        RECT 122.180 94.630 123.830 94.800 ;
        RECT 122.180 69.350 122.350 94.630 ;
        RECT 122.830 91.990 123.180 94.150 ;
        RECT 122.830 69.830 123.180 71.990 ;
        RECT 123.660 69.350 123.830 94.630 ;
        RECT 122.180 69.180 123.830 69.350 ;
        RECT 125.180 94.630 126.830 94.800 ;
        RECT 125.180 69.350 125.350 94.630 ;
        RECT 125.830 91.990 126.180 94.150 ;
        RECT 125.830 69.830 126.180 71.990 ;
        RECT 126.660 69.350 126.830 94.630 ;
        RECT 125.180 69.180 126.830 69.350 ;
        RECT 128.180 94.630 129.830 94.800 ;
        RECT 128.180 69.350 128.350 94.630 ;
        RECT 128.830 91.990 129.180 94.150 ;
        RECT 128.830 69.830 129.180 71.990 ;
        RECT 129.660 69.350 129.830 94.630 ;
        RECT 128.180 69.180 129.830 69.350 ;
      LAYER mcon ;
        RECT 18.425 206.255 18.595 206.425 ;
        RECT 18.885 206.255 19.055 206.425 ;
        RECT 19.345 206.255 19.515 206.425 ;
        RECT 19.805 206.255 19.975 206.425 ;
        RECT 20.265 206.255 20.435 206.425 ;
        RECT 20.725 206.255 20.895 206.425 ;
        RECT 21.185 206.255 21.355 206.425 ;
        RECT 21.645 206.255 21.815 206.425 ;
        RECT 22.105 206.255 22.275 206.425 ;
        RECT 22.565 206.255 22.735 206.425 ;
        RECT 23.025 206.255 23.195 206.425 ;
        RECT 23.485 206.255 23.655 206.425 ;
        RECT 23.945 206.255 24.115 206.425 ;
        RECT 24.405 206.255 24.575 206.425 ;
        RECT 24.865 206.255 25.035 206.425 ;
        RECT 25.325 206.255 25.495 206.425 ;
        RECT 25.785 206.255 25.955 206.425 ;
        RECT 26.245 206.255 26.415 206.425 ;
        RECT 26.705 206.255 26.875 206.425 ;
        RECT 27.165 206.255 27.335 206.425 ;
        RECT 27.625 206.255 27.795 206.425 ;
        RECT 28.085 206.255 28.255 206.425 ;
        RECT 28.545 206.255 28.715 206.425 ;
        RECT 29.005 206.255 29.175 206.425 ;
        RECT 29.465 206.255 29.635 206.425 ;
        RECT 29.925 206.255 30.095 206.425 ;
        RECT 30.385 206.255 30.555 206.425 ;
        RECT 30.845 206.255 31.015 206.425 ;
        RECT 31.305 206.255 31.475 206.425 ;
        RECT 31.765 206.255 31.935 206.425 ;
        RECT 32.225 206.255 32.395 206.425 ;
        RECT 32.685 206.255 32.855 206.425 ;
        RECT 33.145 206.255 33.315 206.425 ;
        RECT 33.605 206.255 33.775 206.425 ;
        RECT 34.065 206.255 34.235 206.425 ;
        RECT 34.525 206.255 34.695 206.425 ;
        RECT 34.985 206.255 35.155 206.425 ;
        RECT 35.445 206.255 35.615 206.425 ;
        RECT 35.905 206.255 36.075 206.425 ;
        RECT 36.365 206.255 36.535 206.425 ;
        RECT 36.825 206.255 36.995 206.425 ;
        RECT 37.285 206.255 37.455 206.425 ;
        RECT 37.745 206.255 37.915 206.425 ;
        RECT 38.205 206.255 38.375 206.425 ;
        RECT 38.665 206.255 38.835 206.425 ;
        RECT 39.125 206.255 39.295 206.425 ;
        RECT 39.585 206.255 39.755 206.425 ;
        RECT 40.045 206.255 40.215 206.425 ;
        RECT 40.505 206.255 40.675 206.425 ;
        RECT 40.965 206.255 41.135 206.425 ;
        RECT 41.425 206.255 41.595 206.425 ;
        RECT 41.885 206.255 42.055 206.425 ;
        RECT 42.345 206.255 42.515 206.425 ;
        RECT 42.805 206.255 42.975 206.425 ;
        RECT 43.265 206.255 43.435 206.425 ;
        RECT 43.725 206.255 43.895 206.425 ;
        RECT 44.185 206.255 44.355 206.425 ;
        RECT 44.645 206.255 44.815 206.425 ;
        RECT 45.105 206.255 45.275 206.425 ;
        RECT 45.565 206.255 45.735 206.425 ;
        RECT 46.025 206.255 46.195 206.425 ;
        RECT 46.485 206.255 46.655 206.425 ;
        RECT 46.945 206.255 47.115 206.425 ;
        RECT 47.405 206.255 47.575 206.425 ;
        RECT 47.865 206.255 48.035 206.425 ;
        RECT 48.325 206.255 48.495 206.425 ;
        RECT 48.785 206.255 48.955 206.425 ;
        RECT 49.245 206.255 49.415 206.425 ;
        RECT 49.705 206.255 49.875 206.425 ;
        RECT 50.165 206.255 50.335 206.425 ;
        RECT 50.625 206.255 50.795 206.425 ;
        RECT 51.085 206.255 51.255 206.425 ;
        RECT 51.545 206.255 51.715 206.425 ;
        RECT 52.005 206.255 52.175 206.425 ;
        RECT 52.465 206.255 52.635 206.425 ;
        RECT 52.925 206.255 53.095 206.425 ;
        RECT 53.385 206.255 53.555 206.425 ;
        RECT 53.845 206.255 54.015 206.425 ;
        RECT 54.305 206.255 54.475 206.425 ;
        RECT 54.765 206.255 54.935 206.425 ;
        RECT 55.225 206.255 55.395 206.425 ;
        RECT 55.685 206.255 55.855 206.425 ;
        RECT 56.145 206.255 56.315 206.425 ;
        RECT 56.605 206.255 56.775 206.425 ;
        RECT 57.065 206.255 57.235 206.425 ;
        RECT 57.525 206.255 57.695 206.425 ;
        RECT 57.985 206.255 58.155 206.425 ;
        RECT 58.445 206.255 58.615 206.425 ;
        RECT 58.905 206.255 59.075 206.425 ;
        RECT 59.365 206.255 59.535 206.425 ;
        RECT 59.825 206.255 59.995 206.425 ;
        RECT 60.285 206.255 60.455 206.425 ;
        RECT 60.745 206.255 60.915 206.425 ;
        RECT 61.205 206.255 61.375 206.425 ;
        RECT 61.665 206.255 61.835 206.425 ;
        RECT 62.125 206.255 62.295 206.425 ;
        RECT 62.585 206.255 62.755 206.425 ;
        RECT 63.045 206.255 63.215 206.425 ;
        RECT 63.505 206.255 63.675 206.425 ;
        RECT 63.965 206.255 64.135 206.425 ;
        RECT 64.425 206.255 64.595 206.425 ;
        RECT 64.885 206.255 65.055 206.425 ;
        RECT 65.345 206.255 65.515 206.425 ;
        RECT 65.805 206.255 65.975 206.425 ;
        RECT 66.265 206.255 66.435 206.425 ;
        RECT 66.725 206.255 66.895 206.425 ;
        RECT 67.185 206.255 67.355 206.425 ;
        RECT 67.645 206.255 67.815 206.425 ;
        RECT 68.105 206.255 68.275 206.425 ;
        RECT 68.565 206.255 68.735 206.425 ;
        RECT 69.025 206.255 69.195 206.425 ;
        RECT 69.485 206.255 69.655 206.425 ;
        RECT 69.945 206.255 70.115 206.425 ;
        RECT 70.405 206.255 70.575 206.425 ;
        RECT 70.865 206.255 71.035 206.425 ;
        RECT 71.325 206.255 71.495 206.425 ;
        RECT 71.785 206.255 71.955 206.425 ;
        RECT 72.245 206.255 72.415 206.425 ;
        RECT 72.705 206.255 72.875 206.425 ;
        RECT 73.165 206.255 73.335 206.425 ;
        RECT 73.625 206.255 73.795 206.425 ;
        RECT 74.085 206.255 74.255 206.425 ;
        RECT 74.545 206.255 74.715 206.425 ;
        RECT 75.005 206.255 75.175 206.425 ;
        RECT 75.465 206.255 75.635 206.425 ;
        RECT 75.925 206.255 76.095 206.425 ;
        RECT 76.385 206.255 76.555 206.425 ;
        RECT 76.845 206.255 77.015 206.425 ;
        RECT 77.305 206.255 77.475 206.425 ;
        RECT 77.765 206.255 77.935 206.425 ;
        RECT 78.225 206.255 78.395 206.425 ;
        RECT 78.685 206.255 78.855 206.425 ;
        RECT 79.145 206.255 79.315 206.425 ;
        RECT 79.605 206.255 79.775 206.425 ;
        RECT 80.065 206.255 80.235 206.425 ;
        RECT 80.525 206.255 80.695 206.425 ;
        RECT 80.985 206.255 81.155 206.425 ;
        RECT 81.445 206.255 81.615 206.425 ;
        RECT 81.905 206.255 82.075 206.425 ;
        RECT 82.365 206.255 82.535 206.425 ;
        RECT 82.825 206.255 82.995 206.425 ;
        RECT 83.285 206.255 83.455 206.425 ;
        RECT 83.745 206.255 83.915 206.425 ;
        RECT 84.205 206.255 84.375 206.425 ;
        RECT 84.665 206.255 84.835 206.425 ;
        RECT 85.125 206.255 85.295 206.425 ;
        RECT 85.585 206.255 85.755 206.425 ;
        RECT 86.045 206.255 86.215 206.425 ;
        RECT 86.505 206.255 86.675 206.425 ;
        RECT 86.965 206.255 87.135 206.425 ;
        RECT 87.425 206.255 87.595 206.425 ;
        RECT 87.885 206.255 88.055 206.425 ;
        RECT 88.345 206.255 88.515 206.425 ;
        RECT 88.805 206.255 88.975 206.425 ;
        RECT 89.265 206.255 89.435 206.425 ;
        RECT 89.725 206.255 89.895 206.425 ;
        RECT 90.185 206.255 90.355 206.425 ;
        RECT 90.645 206.255 90.815 206.425 ;
        RECT 91.105 206.255 91.275 206.425 ;
        RECT 91.565 206.255 91.735 206.425 ;
        RECT 92.025 206.255 92.195 206.425 ;
        RECT 20.725 204.725 20.895 204.895 ;
        RECT 21.645 205.065 21.815 205.235 ;
        RECT 28.085 205.405 28.255 205.575 ;
        RECT 27.165 204.725 27.335 204.895 ;
        RECT 33.145 204.725 33.315 204.895 ;
        RECT 34.065 204.045 34.235 204.215 ;
        RECT 40.045 205.745 40.215 205.915 ;
        RECT 40.045 204.725 40.215 204.895 ;
        RECT 41.425 204.725 41.595 204.895 ;
        RECT 41.885 204.725 42.055 204.895 ;
        RECT 38.665 204.045 38.835 204.215 ;
        RECT 46.025 204.725 46.195 204.895 ;
        RECT 42.805 204.045 42.975 204.215 ;
        RECT 46.945 204.045 47.115 204.215 ;
        RECT 52.465 204.725 52.635 204.895 ;
        RECT 53.385 204.045 53.555 204.215 ;
        RECT 59.825 205.745 59.995 205.915 ;
        RECT 58.905 204.725 59.075 204.895 ;
        RECT 60.285 204.725 60.455 204.895 ;
        RECT 60.745 204.725 60.915 204.895 ;
        RECT 57.525 204.045 57.695 204.215 ;
        RECT 61.665 204.045 61.835 204.215 ;
        RECT 65.345 204.725 65.515 204.895 ;
        RECT 66.265 204.045 66.435 204.215 ;
        RECT 71.785 204.725 71.955 204.895 ;
        RECT 72.705 204.045 72.875 204.215 ;
        RECT 79.145 204.725 79.315 204.895 ;
        RECT 78.225 204.045 78.395 204.215 ;
        RECT 79.605 204.045 79.775 204.215 ;
        RECT 84.665 204.725 84.835 204.895 ;
        RECT 85.585 204.045 85.755 204.215 ;
        RECT 18.425 203.535 18.595 203.705 ;
        RECT 18.885 203.535 19.055 203.705 ;
        RECT 19.345 203.535 19.515 203.705 ;
        RECT 19.805 203.535 19.975 203.705 ;
        RECT 20.265 203.535 20.435 203.705 ;
        RECT 20.725 203.535 20.895 203.705 ;
        RECT 21.185 203.535 21.355 203.705 ;
        RECT 21.645 203.535 21.815 203.705 ;
        RECT 22.105 203.535 22.275 203.705 ;
        RECT 22.565 203.535 22.735 203.705 ;
        RECT 23.025 203.535 23.195 203.705 ;
        RECT 23.485 203.535 23.655 203.705 ;
        RECT 23.945 203.535 24.115 203.705 ;
        RECT 24.405 203.535 24.575 203.705 ;
        RECT 24.865 203.535 25.035 203.705 ;
        RECT 25.325 203.535 25.495 203.705 ;
        RECT 25.785 203.535 25.955 203.705 ;
        RECT 26.245 203.535 26.415 203.705 ;
        RECT 26.705 203.535 26.875 203.705 ;
        RECT 27.165 203.535 27.335 203.705 ;
        RECT 27.625 203.535 27.795 203.705 ;
        RECT 28.085 203.535 28.255 203.705 ;
        RECT 28.545 203.535 28.715 203.705 ;
        RECT 29.005 203.535 29.175 203.705 ;
        RECT 29.465 203.535 29.635 203.705 ;
        RECT 29.925 203.535 30.095 203.705 ;
        RECT 30.385 203.535 30.555 203.705 ;
        RECT 30.845 203.535 31.015 203.705 ;
        RECT 31.305 203.535 31.475 203.705 ;
        RECT 31.765 203.535 31.935 203.705 ;
        RECT 32.225 203.535 32.395 203.705 ;
        RECT 32.685 203.535 32.855 203.705 ;
        RECT 33.145 203.535 33.315 203.705 ;
        RECT 33.605 203.535 33.775 203.705 ;
        RECT 34.065 203.535 34.235 203.705 ;
        RECT 34.525 203.535 34.695 203.705 ;
        RECT 34.985 203.535 35.155 203.705 ;
        RECT 35.445 203.535 35.615 203.705 ;
        RECT 35.905 203.535 36.075 203.705 ;
        RECT 36.365 203.535 36.535 203.705 ;
        RECT 36.825 203.535 36.995 203.705 ;
        RECT 37.285 203.535 37.455 203.705 ;
        RECT 37.745 203.535 37.915 203.705 ;
        RECT 38.205 203.535 38.375 203.705 ;
        RECT 38.665 203.535 38.835 203.705 ;
        RECT 39.125 203.535 39.295 203.705 ;
        RECT 39.585 203.535 39.755 203.705 ;
        RECT 40.045 203.535 40.215 203.705 ;
        RECT 40.505 203.535 40.675 203.705 ;
        RECT 40.965 203.535 41.135 203.705 ;
        RECT 41.425 203.535 41.595 203.705 ;
        RECT 41.885 203.535 42.055 203.705 ;
        RECT 42.345 203.535 42.515 203.705 ;
        RECT 42.805 203.535 42.975 203.705 ;
        RECT 43.265 203.535 43.435 203.705 ;
        RECT 43.725 203.535 43.895 203.705 ;
        RECT 44.185 203.535 44.355 203.705 ;
        RECT 44.645 203.535 44.815 203.705 ;
        RECT 45.105 203.535 45.275 203.705 ;
        RECT 45.565 203.535 45.735 203.705 ;
        RECT 46.025 203.535 46.195 203.705 ;
        RECT 46.485 203.535 46.655 203.705 ;
        RECT 46.945 203.535 47.115 203.705 ;
        RECT 47.405 203.535 47.575 203.705 ;
        RECT 47.865 203.535 48.035 203.705 ;
        RECT 48.325 203.535 48.495 203.705 ;
        RECT 48.785 203.535 48.955 203.705 ;
        RECT 49.245 203.535 49.415 203.705 ;
        RECT 49.705 203.535 49.875 203.705 ;
        RECT 50.165 203.535 50.335 203.705 ;
        RECT 50.625 203.535 50.795 203.705 ;
        RECT 51.085 203.535 51.255 203.705 ;
        RECT 51.545 203.535 51.715 203.705 ;
        RECT 52.005 203.535 52.175 203.705 ;
        RECT 52.465 203.535 52.635 203.705 ;
        RECT 52.925 203.535 53.095 203.705 ;
        RECT 53.385 203.535 53.555 203.705 ;
        RECT 53.845 203.535 54.015 203.705 ;
        RECT 54.305 203.535 54.475 203.705 ;
        RECT 54.765 203.535 54.935 203.705 ;
        RECT 55.225 203.535 55.395 203.705 ;
        RECT 55.685 203.535 55.855 203.705 ;
        RECT 56.145 203.535 56.315 203.705 ;
        RECT 56.605 203.535 56.775 203.705 ;
        RECT 57.065 203.535 57.235 203.705 ;
        RECT 57.525 203.535 57.695 203.705 ;
        RECT 57.985 203.535 58.155 203.705 ;
        RECT 58.445 203.535 58.615 203.705 ;
        RECT 58.905 203.535 59.075 203.705 ;
        RECT 59.365 203.535 59.535 203.705 ;
        RECT 59.825 203.535 59.995 203.705 ;
        RECT 60.285 203.535 60.455 203.705 ;
        RECT 60.745 203.535 60.915 203.705 ;
        RECT 61.205 203.535 61.375 203.705 ;
        RECT 61.665 203.535 61.835 203.705 ;
        RECT 62.125 203.535 62.295 203.705 ;
        RECT 62.585 203.535 62.755 203.705 ;
        RECT 63.045 203.535 63.215 203.705 ;
        RECT 63.505 203.535 63.675 203.705 ;
        RECT 63.965 203.535 64.135 203.705 ;
        RECT 64.425 203.535 64.595 203.705 ;
        RECT 64.885 203.535 65.055 203.705 ;
        RECT 65.345 203.535 65.515 203.705 ;
        RECT 65.805 203.535 65.975 203.705 ;
        RECT 66.265 203.535 66.435 203.705 ;
        RECT 66.725 203.535 66.895 203.705 ;
        RECT 67.185 203.535 67.355 203.705 ;
        RECT 67.645 203.535 67.815 203.705 ;
        RECT 68.105 203.535 68.275 203.705 ;
        RECT 68.565 203.535 68.735 203.705 ;
        RECT 69.025 203.535 69.195 203.705 ;
        RECT 69.485 203.535 69.655 203.705 ;
        RECT 69.945 203.535 70.115 203.705 ;
        RECT 70.405 203.535 70.575 203.705 ;
        RECT 70.865 203.535 71.035 203.705 ;
        RECT 71.325 203.535 71.495 203.705 ;
        RECT 71.785 203.535 71.955 203.705 ;
        RECT 72.245 203.535 72.415 203.705 ;
        RECT 72.705 203.535 72.875 203.705 ;
        RECT 73.165 203.535 73.335 203.705 ;
        RECT 73.625 203.535 73.795 203.705 ;
        RECT 74.085 203.535 74.255 203.705 ;
        RECT 74.545 203.535 74.715 203.705 ;
        RECT 75.005 203.535 75.175 203.705 ;
        RECT 75.465 203.535 75.635 203.705 ;
        RECT 75.925 203.535 76.095 203.705 ;
        RECT 76.385 203.535 76.555 203.705 ;
        RECT 76.845 203.535 77.015 203.705 ;
        RECT 77.305 203.535 77.475 203.705 ;
        RECT 77.765 203.535 77.935 203.705 ;
        RECT 78.225 203.535 78.395 203.705 ;
        RECT 78.685 203.535 78.855 203.705 ;
        RECT 79.145 203.535 79.315 203.705 ;
        RECT 79.605 203.535 79.775 203.705 ;
        RECT 80.065 203.535 80.235 203.705 ;
        RECT 80.525 203.535 80.695 203.705 ;
        RECT 80.985 203.535 81.155 203.705 ;
        RECT 81.445 203.535 81.615 203.705 ;
        RECT 81.905 203.535 82.075 203.705 ;
        RECT 82.365 203.535 82.535 203.705 ;
        RECT 82.825 203.535 82.995 203.705 ;
        RECT 83.285 203.535 83.455 203.705 ;
        RECT 83.745 203.535 83.915 203.705 ;
        RECT 84.205 203.535 84.375 203.705 ;
        RECT 84.665 203.535 84.835 203.705 ;
        RECT 85.125 203.535 85.295 203.705 ;
        RECT 85.585 203.535 85.755 203.705 ;
        RECT 86.045 203.535 86.215 203.705 ;
        RECT 86.505 203.535 86.675 203.705 ;
        RECT 86.965 203.535 87.135 203.705 ;
        RECT 87.425 203.535 87.595 203.705 ;
        RECT 87.885 203.535 88.055 203.705 ;
        RECT 88.345 203.535 88.515 203.705 ;
        RECT 88.805 203.535 88.975 203.705 ;
        RECT 89.265 203.535 89.435 203.705 ;
        RECT 89.725 203.535 89.895 203.705 ;
        RECT 90.185 203.535 90.355 203.705 ;
        RECT 90.645 203.535 90.815 203.705 ;
        RECT 91.105 203.535 91.275 203.705 ;
        RECT 91.565 203.535 91.735 203.705 ;
        RECT 92.025 203.535 92.195 203.705 ;
        RECT 34.065 201.325 34.235 201.495 ;
        RECT 36.375 202.005 36.545 202.175 ;
        RECT 36.810 201.665 36.980 201.835 ;
        RECT 38.895 202.005 39.065 202.175 ;
        RECT 38.380 201.665 38.550 201.835 ;
        RECT 39.685 202.345 39.855 202.515 ;
        RECT 40.085 202.005 40.255 202.175 ;
        RECT 40.965 202.345 41.135 202.515 ;
        RECT 40.480 201.665 40.650 201.835 ;
        RECT 44.645 203.025 44.815 203.195 ;
        RECT 42.805 202.345 42.975 202.515 ;
        RECT 41.885 201.325 42.055 201.495 ;
        RECT 46.955 202.005 47.125 202.175 ;
        RECT 47.390 201.665 47.560 201.835 ;
        RECT 49.475 202.005 49.645 202.175 ;
        RECT 48.960 201.665 49.130 201.835 ;
        RECT 50.210 202.345 50.380 202.515 ;
        RECT 50.665 202.005 50.835 202.175 ;
        RECT 51.545 202.345 51.715 202.515 ;
        RECT 56.145 203.025 56.315 203.195 ;
        RECT 53.385 202.345 53.555 202.515 ;
        RECT 54.765 202.345 54.935 202.515 ;
        RECT 51.060 201.665 51.230 201.835 ;
        RECT 52.005 201.325 52.175 201.495 ;
        RECT 52.925 201.325 53.095 201.495 ;
        RECT 58.455 202.005 58.625 202.175 ;
        RECT 58.890 201.665 59.060 201.835 ;
        RECT 60.975 202.005 61.145 202.175 ;
        RECT 60.460 201.665 60.630 201.835 ;
        RECT 61.710 202.345 61.880 202.515 ;
        RECT 62.165 202.005 62.335 202.175 ;
        RECT 63.045 202.005 63.215 202.175 ;
        RECT 62.560 201.665 62.730 201.835 ;
        RECT 66.265 202.005 66.435 202.175 ;
        RECT 68.105 202.005 68.275 202.175 ;
        RECT 69.485 202.345 69.655 202.515 ;
        RECT 68.565 202.005 68.735 202.175 ;
        RECT 70.405 201.325 70.575 201.495 ;
        RECT 72.715 202.005 72.885 202.175 ;
        RECT 73.150 201.665 73.320 201.835 ;
        RECT 75.235 202.005 75.405 202.175 ;
        RECT 74.720 201.665 74.890 201.835 ;
        RECT 75.970 202.345 76.140 202.515 ;
        RECT 76.425 202.005 76.595 202.175 ;
        RECT 77.305 202.345 77.475 202.515 ;
        RECT 77.765 202.345 77.935 202.515 ;
        RECT 78.230 202.345 78.400 202.515 ;
        RECT 76.820 201.665 76.990 201.835 ;
        RECT 79.145 202.685 79.315 202.855 ;
        RECT 78.635 201.665 78.805 201.835 ;
        RECT 80.065 202.345 80.235 202.515 ;
        RECT 81.425 202.685 81.595 202.855 ;
        RECT 81.785 202.685 81.955 202.855 ;
        RECT 80.525 201.665 80.695 201.835 ;
        RECT 83.645 202.345 83.815 202.515 ;
        RECT 85.025 202.685 85.195 202.855 ;
        RECT 84.725 202.370 84.895 202.540 ;
        RECT 83.645 201.665 83.815 201.835 ;
        RECT 87.425 202.345 87.595 202.515 ;
        RECT 86.505 201.325 86.675 201.495 ;
        RECT 87.885 202.005 88.055 202.175 ;
        RECT 18.425 200.815 18.595 200.985 ;
        RECT 18.885 200.815 19.055 200.985 ;
        RECT 19.345 200.815 19.515 200.985 ;
        RECT 19.805 200.815 19.975 200.985 ;
        RECT 20.265 200.815 20.435 200.985 ;
        RECT 20.725 200.815 20.895 200.985 ;
        RECT 21.185 200.815 21.355 200.985 ;
        RECT 21.645 200.815 21.815 200.985 ;
        RECT 22.105 200.815 22.275 200.985 ;
        RECT 22.565 200.815 22.735 200.985 ;
        RECT 23.025 200.815 23.195 200.985 ;
        RECT 23.485 200.815 23.655 200.985 ;
        RECT 23.945 200.815 24.115 200.985 ;
        RECT 24.405 200.815 24.575 200.985 ;
        RECT 24.865 200.815 25.035 200.985 ;
        RECT 25.325 200.815 25.495 200.985 ;
        RECT 25.785 200.815 25.955 200.985 ;
        RECT 26.245 200.815 26.415 200.985 ;
        RECT 26.705 200.815 26.875 200.985 ;
        RECT 27.165 200.815 27.335 200.985 ;
        RECT 27.625 200.815 27.795 200.985 ;
        RECT 28.085 200.815 28.255 200.985 ;
        RECT 28.545 200.815 28.715 200.985 ;
        RECT 29.005 200.815 29.175 200.985 ;
        RECT 29.465 200.815 29.635 200.985 ;
        RECT 29.925 200.815 30.095 200.985 ;
        RECT 30.385 200.815 30.555 200.985 ;
        RECT 30.845 200.815 31.015 200.985 ;
        RECT 31.305 200.815 31.475 200.985 ;
        RECT 31.765 200.815 31.935 200.985 ;
        RECT 32.225 200.815 32.395 200.985 ;
        RECT 32.685 200.815 32.855 200.985 ;
        RECT 33.145 200.815 33.315 200.985 ;
        RECT 33.605 200.815 33.775 200.985 ;
        RECT 34.065 200.815 34.235 200.985 ;
        RECT 34.525 200.815 34.695 200.985 ;
        RECT 34.985 200.815 35.155 200.985 ;
        RECT 35.445 200.815 35.615 200.985 ;
        RECT 35.905 200.815 36.075 200.985 ;
        RECT 36.365 200.815 36.535 200.985 ;
        RECT 36.825 200.815 36.995 200.985 ;
        RECT 37.285 200.815 37.455 200.985 ;
        RECT 37.745 200.815 37.915 200.985 ;
        RECT 38.205 200.815 38.375 200.985 ;
        RECT 38.665 200.815 38.835 200.985 ;
        RECT 39.125 200.815 39.295 200.985 ;
        RECT 39.585 200.815 39.755 200.985 ;
        RECT 40.045 200.815 40.215 200.985 ;
        RECT 40.505 200.815 40.675 200.985 ;
        RECT 40.965 200.815 41.135 200.985 ;
        RECT 41.425 200.815 41.595 200.985 ;
        RECT 41.885 200.815 42.055 200.985 ;
        RECT 42.345 200.815 42.515 200.985 ;
        RECT 42.805 200.815 42.975 200.985 ;
        RECT 43.265 200.815 43.435 200.985 ;
        RECT 43.725 200.815 43.895 200.985 ;
        RECT 44.185 200.815 44.355 200.985 ;
        RECT 44.645 200.815 44.815 200.985 ;
        RECT 45.105 200.815 45.275 200.985 ;
        RECT 45.565 200.815 45.735 200.985 ;
        RECT 46.025 200.815 46.195 200.985 ;
        RECT 46.485 200.815 46.655 200.985 ;
        RECT 46.945 200.815 47.115 200.985 ;
        RECT 47.405 200.815 47.575 200.985 ;
        RECT 47.865 200.815 48.035 200.985 ;
        RECT 48.325 200.815 48.495 200.985 ;
        RECT 48.785 200.815 48.955 200.985 ;
        RECT 49.245 200.815 49.415 200.985 ;
        RECT 49.705 200.815 49.875 200.985 ;
        RECT 50.165 200.815 50.335 200.985 ;
        RECT 50.625 200.815 50.795 200.985 ;
        RECT 51.085 200.815 51.255 200.985 ;
        RECT 51.545 200.815 51.715 200.985 ;
        RECT 52.005 200.815 52.175 200.985 ;
        RECT 52.465 200.815 52.635 200.985 ;
        RECT 52.925 200.815 53.095 200.985 ;
        RECT 53.385 200.815 53.555 200.985 ;
        RECT 53.845 200.815 54.015 200.985 ;
        RECT 54.305 200.815 54.475 200.985 ;
        RECT 54.765 200.815 54.935 200.985 ;
        RECT 55.225 200.815 55.395 200.985 ;
        RECT 55.685 200.815 55.855 200.985 ;
        RECT 56.145 200.815 56.315 200.985 ;
        RECT 56.605 200.815 56.775 200.985 ;
        RECT 57.065 200.815 57.235 200.985 ;
        RECT 57.525 200.815 57.695 200.985 ;
        RECT 57.985 200.815 58.155 200.985 ;
        RECT 58.445 200.815 58.615 200.985 ;
        RECT 58.905 200.815 59.075 200.985 ;
        RECT 59.365 200.815 59.535 200.985 ;
        RECT 59.825 200.815 59.995 200.985 ;
        RECT 60.285 200.815 60.455 200.985 ;
        RECT 60.745 200.815 60.915 200.985 ;
        RECT 61.205 200.815 61.375 200.985 ;
        RECT 61.665 200.815 61.835 200.985 ;
        RECT 62.125 200.815 62.295 200.985 ;
        RECT 62.585 200.815 62.755 200.985 ;
        RECT 63.045 200.815 63.215 200.985 ;
        RECT 63.505 200.815 63.675 200.985 ;
        RECT 63.965 200.815 64.135 200.985 ;
        RECT 64.425 200.815 64.595 200.985 ;
        RECT 64.885 200.815 65.055 200.985 ;
        RECT 65.345 200.815 65.515 200.985 ;
        RECT 65.805 200.815 65.975 200.985 ;
        RECT 66.265 200.815 66.435 200.985 ;
        RECT 66.725 200.815 66.895 200.985 ;
        RECT 67.185 200.815 67.355 200.985 ;
        RECT 67.645 200.815 67.815 200.985 ;
        RECT 68.105 200.815 68.275 200.985 ;
        RECT 68.565 200.815 68.735 200.985 ;
        RECT 69.025 200.815 69.195 200.985 ;
        RECT 69.485 200.815 69.655 200.985 ;
        RECT 69.945 200.815 70.115 200.985 ;
        RECT 70.405 200.815 70.575 200.985 ;
        RECT 70.865 200.815 71.035 200.985 ;
        RECT 71.325 200.815 71.495 200.985 ;
        RECT 71.785 200.815 71.955 200.985 ;
        RECT 72.245 200.815 72.415 200.985 ;
        RECT 72.705 200.815 72.875 200.985 ;
        RECT 73.165 200.815 73.335 200.985 ;
        RECT 73.625 200.815 73.795 200.985 ;
        RECT 74.085 200.815 74.255 200.985 ;
        RECT 74.545 200.815 74.715 200.985 ;
        RECT 75.005 200.815 75.175 200.985 ;
        RECT 75.465 200.815 75.635 200.985 ;
        RECT 75.925 200.815 76.095 200.985 ;
        RECT 76.385 200.815 76.555 200.985 ;
        RECT 76.845 200.815 77.015 200.985 ;
        RECT 77.305 200.815 77.475 200.985 ;
        RECT 77.765 200.815 77.935 200.985 ;
        RECT 78.225 200.815 78.395 200.985 ;
        RECT 78.685 200.815 78.855 200.985 ;
        RECT 79.145 200.815 79.315 200.985 ;
        RECT 79.605 200.815 79.775 200.985 ;
        RECT 80.065 200.815 80.235 200.985 ;
        RECT 80.525 200.815 80.695 200.985 ;
        RECT 80.985 200.815 81.155 200.985 ;
        RECT 81.445 200.815 81.615 200.985 ;
        RECT 81.905 200.815 82.075 200.985 ;
        RECT 82.365 200.815 82.535 200.985 ;
        RECT 82.825 200.815 82.995 200.985 ;
        RECT 83.285 200.815 83.455 200.985 ;
        RECT 83.745 200.815 83.915 200.985 ;
        RECT 84.205 200.815 84.375 200.985 ;
        RECT 84.665 200.815 84.835 200.985 ;
        RECT 85.125 200.815 85.295 200.985 ;
        RECT 85.585 200.815 85.755 200.985 ;
        RECT 86.045 200.815 86.215 200.985 ;
        RECT 86.505 200.815 86.675 200.985 ;
        RECT 86.965 200.815 87.135 200.985 ;
        RECT 87.425 200.815 87.595 200.985 ;
        RECT 87.885 200.815 88.055 200.985 ;
        RECT 88.345 200.815 88.515 200.985 ;
        RECT 88.805 200.815 88.975 200.985 ;
        RECT 89.265 200.815 89.435 200.985 ;
        RECT 89.725 200.815 89.895 200.985 ;
        RECT 90.185 200.815 90.355 200.985 ;
        RECT 90.645 200.815 90.815 200.985 ;
        RECT 91.105 200.815 91.275 200.985 ;
        RECT 91.565 200.815 91.735 200.985 ;
        RECT 92.025 200.815 92.195 200.985 ;
        RECT 37.285 199.625 37.455 199.795 ;
        RECT 39.125 199.285 39.295 199.455 ;
        RECT 40.505 200.305 40.675 200.475 ;
        RECT 39.585 199.285 39.755 199.455 ;
        RECT 47.405 199.625 47.575 199.795 ;
        RECT 49.245 199.285 49.415 199.455 ;
        RECT 50.625 200.305 50.795 200.475 ;
        RECT 49.705 199.285 49.875 199.455 ;
        RECT 58.445 199.625 58.615 199.795 ;
        RECT 60.285 199.285 60.455 199.455 ;
        RECT 61.665 200.305 61.835 200.475 ;
        RECT 60.745 199.285 60.915 199.455 ;
        RECT 67.645 200.305 67.815 200.475 ;
        RECT 69.945 200.305 70.115 200.475 ;
        RECT 71.785 200.305 71.955 200.475 ;
        RECT 68.565 199.285 68.735 199.455 ;
        RECT 70.375 199.285 70.545 199.455 ;
        RECT 73.165 198.945 73.335 199.115 ;
        RECT 80.065 199.965 80.235 200.135 ;
        RECT 75.005 199.285 75.175 199.455 ;
        RECT 75.925 199.285 76.095 199.455 ;
        RECT 76.385 199.285 76.555 199.455 ;
        RECT 75.465 198.945 75.635 199.115 ;
        RECT 77.305 199.285 77.475 199.455 ;
        RECT 78.685 199.285 78.855 199.455 ;
        RECT 76.845 198.605 77.015 198.775 ;
        RECT 79.145 198.945 79.315 199.115 ;
        RECT 80.065 198.945 80.235 199.115 ;
        RECT 84.665 198.605 84.835 198.775 ;
        RECT 87.885 199.285 88.055 199.455 ;
        RECT 88.345 199.285 88.515 199.455 ;
        RECT 88.805 198.605 88.975 198.775 ;
        RECT 18.425 198.095 18.595 198.265 ;
        RECT 18.885 198.095 19.055 198.265 ;
        RECT 19.345 198.095 19.515 198.265 ;
        RECT 19.805 198.095 19.975 198.265 ;
        RECT 20.265 198.095 20.435 198.265 ;
        RECT 20.725 198.095 20.895 198.265 ;
        RECT 21.185 198.095 21.355 198.265 ;
        RECT 21.645 198.095 21.815 198.265 ;
        RECT 22.105 198.095 22.275 198.265 ;
        RECT 22.565 198.095 22.735 198.265 ;
        RECT 23.025 198.095 23.195 198.265 ;
        RECT 23.485 198.095 23.655 198.265 ;
        RECT 23.945 198.095 24.115 198.265 ;
        RECT 24.405 198.095 24.575 198.265 ;
        RECT 24.865 198.095 25.035 198.265 ;
        RECT 25.325 198.095 25.495 198.265 ;
        RECT 25.785 198.095 25.955 198.265 ;
        RECT 26.245 198.095 26.415 198.265 ;
        RECT 26.705 198.095 26.875 198.265 ;
        RECT 27.165 198.095 27.335 198.265 ;
        RECT 27.625 198.095 27.795 198.265 ;
        RECT 28.085 198.095 28.255 198.265 ;
        RECT 28.545 198.095 28.715 198.265 ;
        RECT 29.005 198.095 29.175 198.265 ;
        RECT 29.465 198.095 29.635 198.265 ;
        RECT 29.925 198.095 30.095 198.265 ;
        RECT 30.385 198.095 30.555 198.265 ;
        RECT 30.845 198.095 31.015 198.265 ;
        RECT 31.305 198.095 31.475 198.265 ;
        RECT 31.765 198.095 31.935 198.265 ;
        RECT 32.225 198.095 32.395 198.265 ;
        RECT 32.685 198.095 32.855 198.265 ;
        RECT 33.145 198.095 33.315 198.265 ;
        RECT 33.605 198.095 33.775 198.265 ;
        RECT 34.065 198.095 34.235 198.265 ;
        RECT 34.525 198.095 34.695 198.265 ;
        RECT 34.985 198.095 35.155 198.265 ;
        RECT 35.445 198.095 35.615 198.265 ;
        RECT 35.905 198.095 36.075 198.265 ;
        RECT 36.365 198.095 36.535 198.265 ;
        RECT 36.825 198.095 36.995 198.265 ;
        RECT 37.285 198.095 37.455 198.265 ;
        RECT 37.745 198.095 37.915 198.265 ;
        RECT 38.205 198.095 38.375 198.265 ;
        RECT 38.665 198.095 38.835 198.265 ;
        RECT 39.125 198.095 39.295 198.265 ;
        RECT 39.585 198.095 39.755 198.265 ;
        RECT 40.045 198.095 40.215 198.265 ;
        RECT 40.505 198.095 40.675 198.265 ;
        RECT 40.965 198.095 41.135 198.265 ;
        RECT 41.425 198.095 41.595 198.265 ;
        RECT 41.885 198.095 42.055 198.265 ;
        RECT 42.345 198.095 42.515 198.265 ;
        RECT 42.805 198.095 42.975 198.265 ;
        RECT 43.265 198.095 43.435 198.265 ;
        RECT 43.725 198.095 43.895 198.265 ;
        RECT 44.185 198.095 44.355 198.265 ;
        RECT 44.645 198.095 44.815 198.265 ;
        RECT 45.105 198.095 45.275 198.265 ;
        RECT 45.565 198.095 45.735 198.265 ;
        RECT 46.025 198.095 46.195 198.265 ;
        RECT 46.485 198.095 46.655 198.265 ;
        RECT 46.945 198.095 47.115 198.265 ;
        RECT 47.405 198.095 47.575 198.265 ;
        RECT 47.865 198.095 48.035 198.265 ;
        RECT 48.325 198.095 48.495 198.265 ;
        RECT 48.785 198.095 48.955 198.265 ;
        RECT 49.245 198.095 49.415 198.265 ;
        RECT 49.705 198.095 49.875 198.265 ;
        RECT 50.165 198.095 50.335 198.265 ;
        RECT 50.625 198.095 50.795 198.265 ;
        RECT 51.085 198.095 51.255 198.265 ;
        RECT 51.545 198.095 51.715 198.265 ;
        RECT 52.005 198.095 52.175 198.265 ;
        RECT 52.465 198.095 52.635 198.265 ;
        RECT 52.925 198.095 53.095 198.265 ;
        RECT 53.385 198.095 53.555 198.265 ;
        RECT 53.845 198.095 54.015 198.265 ;
        RECT 54.305 198.095 54.475 198.265 ;
        RECT 54.765 198.095 54.935 198.265 ;
        RECT 55.225 198.095 55.395 198.265 ;
        RECT 55.685 198.095 55.855 198.265 ;
        RECT 56.145 198.095 56.315 198.265 ;
        RECT 56.605 198.095 56.775 198.265 ;
        RECT 57.065 198.095 57.235 198.265 ;
        RECT 57.525 198.095 57.695 198.265 ;
        RECT 57.985 198.095 58.155 198.265 ;
        RECT 58.445 198.095 58.615 198.265 ;
        RECT 58.905 198.095 59.075 198.265 ;
        RECT 59.365 198.095 59.535 198.265 ;
        RECT 59.825 198.095 59.995 198.265 ;
        RECT 60.285 198.095 60.455 198.265 ;
        RECT 60.745 198.095 60.915 198.265 ;
        RECT 61.205 198.095 61.375 198.265 ;
        RECT 61.665 198.095 61.835 198.265 ;
        RECT 62.125 198.095 62.295 198.265 ;
        RECT 62.585 198.095 62.755 198.265 ;
        RECT 63.045 198.095 63.215 198.265 ;
        RECT 63.505 198.095 63.675 198.265 ;
        RECT 63.965 198.095 64.135 198.265 ;
        RECT 64.425 198.095 64.595 198.265 ;
        RECT 64.885 198.095 65.055 198.265 ;
        RECT 65.345 198.095 65.515 198.265 ;
        RECT 65.805 198.095 65.975 198.265 ;
        RECT 66.265 198.095 66.435 198.265 ;
        RECT 66.725 198.095 66.895 198.265 ;
        RECT 67.185 198.095 67.355 198.265 ;
        RECT 67.645 198.095 67.815 198.265 ;
        RECT 68.105 198.095 68.275 198.265 ;
        RECT 68.565 198.095 68.735 198.265 ;
        RECT 69.025 198.095 69.195 198.265 ;
        RECT 69.485 198.095 69.655 198.265 ;
        RECT 69.945 198.095 70.115 198.265 ;
        RECT 70.405 198.095 70.575 198.265 ;
        RECT 70.865 198.095 71.035 198.265 ;
        RECT 71.325 198.095 71.495 198.265 ;
        RECT 71.785 198.095 71.955 198.265 ;
        RECT 72.245 198.095 72.415 198.265 ;
        RECT 72.705 198.095 72.875 198.265 ;
        RECT 73.165 198.095 73.335 198.265 ;
        RECT 73.625 198.095 73.795 198.265 ;
        RECT 74.085 198.095 74.255 198.265 ;
        RECT 74.545 198.095 74.715 198.265 ;
        RECT 75.005 198.095 75.175 198.265 ;
        RECT 75.465 198.095 75.635 198.265 ;
        RECT 75.925 198.095 76.095 198.265 ;
        RECT 76.385 198.095 76.555 198.265 ;
        RECT 76.845 198.095 77.015 198.265 ;
        RECT 77.305 198.095 77.475 198.265 ;
        RECT 77.765 198.095 77.935 198.265 ;
        RECT 78.225 198.095 78.395 198.265 ;
        RECT 78.685 198.095 78.855 198.265 ;
        RECT 79.145 198.095 79.315 198.265 ;
        RECT 79.605 198.095 79.775 198.265 ;
        RECT 80.065 198.095 80.235 198.265 ;
        RECT 80.525 198.095 80.695 198.265 ;
        RECT 80.985 198.095 81.155 198.265 ;
        RECT 81.445 198.095 81.615 198.265 ;
        RECT 81.905 198.095 82.075 198.265 ;
        RECT 82.365 198.095 82.535 198.265 ;
        RECT 82.825 198.095 82.995 198.265 ;
        RECT 83.285 198.095 83.455 198.265 ;
        RECT 83.745 198.095 83.915 198.265 ;
        RECT 84.205 198.095 84.375 198.265 ;
        RECT 84.665 198.095 84.835 198.265 ;
        RECT 85.125 198.095 85.295 198.265 ;
        RECT 85.585 198.095 85.755 198.265 ;
        RECT 86.045 198.095 86.215 198.265 ;
        RECT 86.505 198.095 86.675 198.265 ;
        RECT 86.965 198.095 87.135 198.265 ;
        RECT 87.425 198.095 87.595 198.265 ;
        RECT 87.885 198.095 88.055 198.265 ;
        RECT 88.345 198.095 88.515 198.265 ;
        RECT 88.805 198.095 88.975 198.265 ;
        RECT 89.265 198.095 89.435 198.265 ;
        RECT 89.725 198.095 89.895 198.265 ;
        RECT 90.185 198.095 90.355 198.265 ;
        RECT 90.645 198.095 90.815 198.265 ;
        RECT 91.105 198.095 91.275 198.265 ;
        RECT 91.565 198.095 91.735 198.265 ;
        RECT 92.025 198.095 92.195 198.265 ;
        RECT 34.985 196.565 35.155 196.735 ;
        RECT 36.825 196.565 36.995 196.735 ;
        RECT 37.285 196.905 37.455 197.075 ;
        RECT 38.205 195.885 38.375 196.055 ;
        RECT 44.645 195.885 44.815 196.055 ;
        RECT 45.565 196.565 45.735 196.735 ;
        RECT 46.025 196.905 46.195 197.075 ;
        RECT 47.865 196.565 48.035 196.735 ;
        RECT 51.545 195.885 51.715 196.055 ;
        RECT 53.855 196.565 54.025 196.735 ;
        RECT 54.290 196.225 54.460 196.395 ;
        RECT 56.375 196.565 56.545 196.735 ;
        RECT 55.860 196.225 56.030 196.395 ;
        RECT 57.165 196.905 57.335 197.075 ;
        RECT 57.565 196.565 57.735 196.735 ;
        RECT 58.445 196.565 58.615 196.735 ;
        RECT 57.960 196.225 58.130 196.395 ;
        RECT 60.745 196.565 60.915 196.735 ;
        RECT 61.230 196.225 61.400 196.395 ;
        RECT 61.625 196.565 61.795 196.735 ;
        RECT 62.080 196.905 62.250 197.075 ;
        RECT 62.815 196.565 62.985 196.735 ;
        RECT 63.330 196.225 63.500 196.395 ;
        RECT 64.900 196.225 65.070 196.395 ;
        RECT 65.335 196.565 65.505 196.735 ;
        RECT 76.385 197.585 76.555 197.755 ;
        RECT 67.645 195.885 67.815 196.055 ;
        RECT 73.855 196.905 74.025 197.075 ;
        RECT 74.545 196.905 74.715 197.075 ;
        RECT 75.005 196.905 75.175 197.075 ;
        RECT 75.465 196.905 75.635 197.075 ;
        RECT 79.145 197.585 79.315 197.755 ;
        RECT 78.225 195.885 78.395 196.055 ;
        RECT 79.145 196.565 79.315 196.735 ;
        RECT 82.365 196.905 82.535 197.075 ;
        RECT 82.830 196.225 83.000 196.395 ;
        RECT 83.290 197.245 83.460 197.415 ;
        RECT 83.745 196.565 83.915 196.735 ;
        RECT 84.690 197.245 84.860 197.415 ;
        RECT 86.530 197.245 86.700 197.415 ;
        RECT 85.150 196.225 85.320 196.395 ;
        RECT 86.530 196.225 86.700 196.395 ;
        RECT 90.185 197.585 90.355 197.755 ;
        RECT 18.425 195.375 18.595 195.545 ;
        RECT 18.885 195.375 19.055 195.545 ;
        RECT 19.345 195.375 19.515 195.545 ;
        RECT 19.805 195.375 19.975 195.545 ;
        RECT 20.265 195.375 20.435 195.545 ;
        RECT 20.725 195.375 20.895 195.545 ;
        RECT 21.185 195.375 21.355 195.545 ;
        RECT 21.645 195.375 21.815 195.545 ;
        RECT 22.105 195.375 22.275 195.545 ;
        RECT 22.565 195.375 22.735 195.545 ;
        RECT 23.025 195.375 23.195 195.545 ;
        RECT 23.485 195.375 23.655 195.545 ;
        RECT 23.945 195.375 24.115 195.545 ;
        RECT 24.405 195.375 24.575 195.545 ;
        RECT 24.865 195.375 25.035 195.545 ;
        RECT 25.325 195.375 25.495 195.545 ;
        RECT 25.785 195.375 25.955 195.545 ;
        RECT 26.245 195.375 26.415 195.545 ;
        RECT 26.705 195.375 26.875 195.545 ;
        RECT 27.165 195.375 27.335 195.545 ;
        RECT 27.625 195.375 27.795 195.545 ;
        RECT 28.085 195.375 28.255 195.545 ;
        RECT 28.545 195.375 28.715 195.545 ;
        RECT 29.005 195.375 29.175 195.545 ;
        RECT 29.465 195.375 29.635 195.545 ;
        RECT 29.925 195.375 30.095 195.545 ;
        RECT 30.385 195.375 30.555 195.545 ;
        RECT 30.845 195.375 31.015 195.545 ;
        RECT 31.305 195.375 31.475 195.545 ;
        RECT 31.765 195.375 31.935 195.545 ;
        RECT 32.225 195.375 32.395 195.545 ;
        RECT 32.685 195.375 32.855 195.545 ;
        RECT 33.145 195.375 33.315 195.545 ;
        RECT 33.605 195.375 33.775 195.545 ;
        RECT 34.065 195.375 34.235 195.545 ;
        RECT 34.525 195.375 34.695 195.545 ;
        RECT 34.985 195.375 35.155 195.545 ;
        RECT 35.445 195.375 35.615 195.545 ;
        RECT 35.905 195.375 36.075 195.545 ;
        RECT 36.365 195.375 36.535 195.545 ;
        RECT 36.825 195.375 36.995 195.545 ;
        RECT 37.285 195.375 37.455 195.545 ;
        RECT 37.745 195.375 37.915 195.545 ;
        RECT 38.205 195.375 38.375 195.545 ;
        RECT 38.665 195.375 38.835 195.545 ;
        RECT 39.125 195.375 39.295 195.545 ;
        RECT 39.585 195.375 39.755 195.545 ;
        RECT 40.045 195.375 40.215 195.545 ;
        RECT 40.505 195.375 40.675 195.545 ;
        RECT 40.965 195.375 41.135 195.545 ;
        RECT 41.425 195.375 41.595 195.545 ;
        RECT 41.885 195.375 42.055 195.545 ;
        RECT 42.345 195.375 42.515 195.545 ;
        RECT 42.805 195.375 42.975 195.545 ;
        RECT 43.265 195.375 43.435 195.545 ;
        RECT 43.725 195.375 43.895 195.545 ;
        RECT 44.185 195.375 44.355 195.545 ;
        RECT 44.645 195.375 44.815 195.545 ;
        RECT 45.105 195.375 45.275 195.545 ;
        RECT 45.565 195.375 45.735 195.545 ;
        RECT 46.025 195.375 46.195 195.545 ;
        RECT 46.485 195.375 46.655 195.545 ;
        RECT 46.945 195.375 47.115 195.545 ;
        RECT 47.405 195.375 47.575 195.545 ;
        RECT 47.865 195.375 48.035 195.545 ;
        RECT 48.325 195.375 48.495 195.545 ;
        RECT 48.785 195.375 48.955 195.545 ;
        RECT 49.245 195.375 49.415 195.545 ;
        RECT 49.705 195.375 49.875 195.545 ;
        RECT 50.165 195.375 50.335 195.545 ;
        RECT 50.625 195.375 50.795 195.545 ;
        RECT 51.085 195.375 51.255 195.545 ;
        RECT 51.545 195.375 51.715 195.545 ;
        RECT 52.005 195.375 52.175 195.545 ;
        RECT 52.465 195.375 52.635 195.545 ;
        RECT 52.925 195.375 53.095 195.545 ;
        RECT 53.385 195.375 53.555 195.545 ;
        RECT 53.845 195.375 54.015 195.545 ;
        RECT 54.305 195.375 54.475 195.545 ;
        RECT 54.765 195.375 54.935 195.545 ;
        RECT 55.225 195.375 55.395 195.545 ;
        RECT 55.685 195.375 55.855 195.545 ;
        RECT 56.145 195.375 56.315 195.545 ;
        RECT 56.605 195.375 56.775 195.545 ;
        RECT 57.065 195.375 57.235 195.545 ;
        RECT 57.525 195.375 57.695 195.545 ;
        RECT 57.985 195.375 58.155 195.545 ;
        RECT 58.445 195.375 58.615 195.545 ;
        RECT 58.905 195.375 59.075 195.545 ;
        RECT 59.365 195.375 59.535 195.545 ;
        RECT 59.825 195.375 59.995 195.545 ;
        RECT 60.285 195.375 60.455 195.545 ;
        RECT 60.745 195.375 60.915 195.545 ;
        RECT 61.205 195.375 61.375 195.545 ;
        RECT 61.665 195.375 61.835 195.545 ;
        RECT 62.125 195.375 62.295 195.545 ;
        RECT 62.585 195.375 62.755 195.545 ;
        RECT 63.045 195.375 63.215 195.545 ;
        RECT 63.505 195.375 63.675 195.545 ;
        RECT 63.965 195.375 64.135 195.545 ;
        RECT 64.425 195.375 64.595 195.545 ;
        RECT 64.885 195.375 65.055 195.545 ;
        RECT 65.345 195.375 65.515 195.545 ;
        RECT 65.805 195.375 65.975 195.545 ;
        RECT 66.265 195.375 66.435 195.545 ;
        RECT 66.725 195.375 66.895 195.545 ;
        RECT 67.185 195.375 67.355 195.545 ;
        RECT 67.645 195.375 67.815 195.545 ;
        RECT 68.105 195.375 68.275 195.545 ;
        RECT 68.565 195.375 68.735 195.545 ;
        RECT 69.025 195.375 69.195 195.545 ;
        RECT 69.485 195.375 69.655 195.545 ;
        RECT 69.945 195.375 70.115 195.545 ;
        RECT 70.405 195.375 70.575 195.545 ;
        RECT 70.865 195.375 71.035 195.545 ;
        RECT 71.325 195.375 71.495 195.545 ;
        RECT 71.785 195.375 71.955 195.545 ;
        RECT 72.245 195.375 72.415 195.545 ;
        RECT 72.705 195.375 72.875 195.545 ;
        RECT 73.165 195.375 73.335 195.545 ;
        RECT 73.625 195.375 73.795 195.545 ;
        RECT 74.085 195.375 74.255 195.545 ;
        RECT 74.545 195.375 74.715 195.545 ;
        RECT 75.005 195.375 75.175 195.545 ;
        RECT 75.465 195.375 75.635 195.545 ;
        RECT 75.925 195.375 76.095 195.545 ;
        RECT 76.385 195.375 76.555 195.545 ;
        RECT 76.845 195.375 77.015 195.545 ;
        RECT 77.305 195.375 77.475 195.545 ;
        RECT 77.765 195.375 77.935 195.545 ;
        RECT 78.225 195.375 78.395 195.545 ;
        RECT 78.685 195.375 78.855 195.545 ;
        RECT 79.145 195.375 79.315 195.545 ;
        RECT 79.605 195.375 79.775 195.545 ;
        RECT 80.065 195.375 80.235 195.545 ;
        RECT 80.525 195.375 80.695 195.545 ;
        RECT 80.985 195.375 81.155 195.545 ;
        RECT 81.445 195.375 81.615 195.545 ;
        RECT 81.905 195.375 82.075 195.545 ;
        RECT 82.365 195.375 82.535 195.545 ;
        RECT 82.825 195.375 82.995 195.545 ;
        RECT 83.285 195.375 83.455 195.545 ;
        RECT 83.745 195.375 83.915 195.545 ;
        RECT 84.205 195.375 84.375 195.545 ;
        RECT 84.665 195.375 84.835 195.545 ;
        RECT 85.125 195.375 85.295 195.545 ;
        RECT 85.585 195.375 85.755 195.545 ;
        RECT 86.045 195.375 86.215 195.545 ;
        RECT 86.505 195.375 86.675 195.545 ;
        RECT 86.965 195.375 87.135 195.545 ;
        RECT 87.425 195.375 87.595 195.545 ;
        RECT 87.885 195.375 88.055 195.545 ;
        RECT 88.345 195.375 88.515 195.545 ;
        RECT 88.805 195.375 88.975 195.545 ;
        RECT 89.265 195.375 89.435 195.545 ;
        RECT 89.725 195.375 89.895 195.545 ;
        RECT 90.185 195.375 90.355 195.545 ;
        RECT 90.645 195.375 90.815 195.545 ;
        RECT 91.105 195.375 91.275 195.545 ;
        RECT 91.565 195.375 91.735 195.545 ;
        RECT 92.025 195.375 92.195 195.545 ;
        RECT 31.765 193.165 31.935 193.335 ;
        RECT 34.075 194.185 34.245 194.355 ;
        RECT 34.510 194.525 34.680 194.695 ;
        RECT 36.080 194.525 36.250 194.695 ;
        RECT 36.595 194.185 36.765 194.355 ;
        RECT 37.385 193.845 37.555 194.015 ;
        RECT 37.785 194.185 37.955 194.355 ;
        RECT 38.180 194.525 38.350 194.695 ;
        RECT 38.665 194.185 38.835 194.355 ;
        RECT 42.370 194.525 42.540 194.695 ;
        RECT 41.885 194.185 42.055 194.355 ;
        RECT 42.765 194.185 42.935 194.355 ;
        RECT 43.220 193.845 43.390 194.015 ;
        RECT 44.470 194.525 44.640 194.695 ;
        RECT 43.955 194.185 44.125 194.355 ;
        RECT 46.040 194.525 46.210 194.695 ;
        RECT 46.475 194.185 46.645 194.355 ;
        RECT 49.245 194.865 49.415 195.035 ;
        RECT 51.085 194.865 51.255 195.035 ;
        RECT 50.625 194.185 50.795 194.355 ;
        RECT 54.305 194.865 54.475 195.035 ;
        RECT 51.055 193.845 51.225 194.015 ;
        RECT 51.545 193.845 51.715 194.015 ;
        RECT 48.785 193.165 48.955 193.335 ;
        RECT 55.225 194.185 55.395 194.355 ;
        RECT 53.845 193.845 54.015 194.015 ;
        RECT 52.005 193.165 52.175 193.335 ;
        RECT 56.605 193.165 56.775 193.335 ;
        RECT 57.525 193.165 57.695 193.335 ;
        RECT 59.365 194.185 59.535 194.355 ;
        RECT 60.745 194.865 60.915 195.035 ;
        RECT 59.825 193.845 59.995 194.015 ;
        RECT 65.345 194.865 65.515 195.035 ;
        RECT 66.265 193.845 66.435 194.015 ;
        RECT 66.725 194.185 66.895 194.355 ;
        RECT 68.565 193.165 68.735 193.335 ;
        RECT 69.945 194.865 70.115 195.035 ;
        RECT 69.945 193.845 70.115 194.015 ;
        RECT 71.785 193.845 71.955 194.015 ;
        RECT 72.245 193.845 72.415 194.015 ;
        RECT 73.165 193.845 73.335 194.015 ;
        RECT 69.025 193.165 69.195 193.335 ;
        RECT 79.145 194.525 79.315 194.695 ;
        RECT 74.545 193.845 74.715 194.015 ;
        RECT 74.085 193.505 74.255 193.675 ;
        RECT 75.465 193.845 75.635 194.015 ;
        RECT 75.925 193.845 76.095 194.015 ;
        RECT 76.385 193.845 76.555 194.015 ;
        RECT 75.005 193.165 75.175 193.335 ;
        RECT 77.765 193.845 77.935 194.015 ;
        RECT 78.225 193.845 78.395 194.015 ;
        RECT 81.445 193.845 81.615 194.015 ;
        RECT 80.525 193.505 80.695 193.675 ;
        RECT 84.665 193.845 84.835 194.015 ;
        RECT 85.125 193.845 85.295 194.015 ;
        RECT 85.585 193.845 85.755 194.015 ;
        RECT 83.285 193.165 83.455 193.335 ;
        RECT 86.505 193.845 86.675 194.015 ;
        RECT 18.425 192.655 18.595 192.825 ;
        RECT 18.885 192.655 19.055 192.825 ;
        RECT 19.345 192.655 19.515 192.825 ;
        RECT 19.805 192.655 19.975 192.825 ;
        RECT 20.265 192.655 20.435 192.825 ;
        RECT 20.725 192.655 20.895 192.825 ;
        RECT 21.185 192.655 21.355 192.825 ;
        RECT 21.645 192.655 21.815 192.825 ;
        RECT 22.105 192.655 22.275 192.825 ;
        RECT 22.565 192.655 22.735 192.825 ;
        RECT 23.025 192.655 23.195 192.825 ;
        RECT 23.485 192.655 23.655 192.825 ;
        RECT 23.945 192.655 24.115 192.825 ;
        RECT 24.405 192.655 24.575 192.825 ;
        RECT 24.865 192.655 25.035 192.825 ;
        RECT 25.325 192.655 25.495 192.825 ;
        RECT 25.785 192.655 25.955 192.825 ;
        RECT 26.245 192.655 26.415 192.825 ;
        RECT 26.705 192.655 26.875 192.825 ;
        RECT 27.165 192.655 27.335 192.825 ;
        RECT 27.625 192.655 27.795 192.825 ;
        RECT 28.085 192.655 28.255 192.825 ;
        RECT 28.545 192.655 28.715 192.825 ;
        RECT 29.005 192.655 29.175 192.825 ;
        RECT 29.465 192.655 29.635 192.825 ;
        RECT 29.925 192.655 30.095 192.825 ;
        RECT 30.385 192.655 30.555 192.825 ;
        RECT 30.845 192.655 31.015 192.825 ;
        RECT 31.305 192.655 31.475 192.825 ;
        RECT 31.765 192.655 31.935 192.825 ;
        RECT 32.225 192.655 32.395 192.825 ;
        RECT 32.685 192.655 32.855 192.825 ;
        RECT 33.145 192.655 33.315 192.825 ;
        RECT 33.605 192.655 33.775 192.825 ;
        RECT 34.065 192.655 34.235 192.825 ;
        RECT 34.525 192.655 34.695 192.825 ;
        RECT 34.985 192.655 35.155 192.825 ;
        RECT 35.445 192.655 35.615 192.825 ;
        RECT 35.905 192.655 36.075 192.825 ;
        RECT 36.365 192.655 36.535 192.825 ;
        RECT 36.825 192.655 36.995 192.825 ;
        RECT 37.285 192.655 37.455 192.825 ;
        RECT 37.745 192.655 37.915 192.825 ;
        RECT 38.205 192.655 38.375 192.825 ;
        RECT 38.665 192.655 38.835 192.825 ;
        RECT 39.125 192.655 39.295 192.825 ;
        RECT 39.585 192.655 39.755 192.825 ;
        RECT 40.045 192.655 40.215 192.825 ;
        RECT 40.505 192.655 40.675 192.825 ;
        RECT 40.965 192.655 41.135 192.825 ;
        RECT 41.425 192.655 41.595 192.825 ;
        RECT 41.885 192.655 42.055 192.825 ;
        RECT 42.345 192.655 42.515 192.825 ;
        RECT 42.805 192.655 42.975 192.825 ;
        RECT 43.265 192.655 43.435 192.825 ;
        RECT 43.725 192.655 43.895 192.825 ;
        RECT 44.185 192.655 44.355 192.825 ;
        RECT 44.645 192.655 44.815 192.825 ;
        RECT 45.105 192.655 45.275 192.825 ;
        RECT 45.565 192.655 45.735 192.825 ;
        RECT 46.025 192.655 46.195 192.825 ;
        RECT 46.485 192.655 46.655 192.825 ;
        RECT 46.945 192.655 47.115 192.825 ;
        RECT 47.405 192.655 47.575 192.825 ;
        RECT 47.865 192.655 48.035 192.825 ;
        RECT 48.325 192.655 48.495 192.825 ;
        RECT 48.785 192.655 48.955 192.825 ;
        RECT 49.245 192.655 49.415 192.825 ;
        RECT 49.705 192.655 49.875 192.825 ;
        RECT 50.165 192.655 50.335 192.825 ;
        RECT 50.625 192.655 50.795 192.825 ;
        RECT 51.085 192.655 51.255 192.825 ;
        RECT 51.545 192.655 51.715 192.825 ;
        RECT 52.005 192.655 52.175 192.825 ;
        RECT 52.465 192.655 52.635 192.825 ;
        RECT 52.925 192.655 53.095 192.825 ;
        RECT 53.385 192.655 53.555 192.825 ;
        RECT 53.845 192.655 54.015 192.825 ;
        RECT 54.305 192.655 54.475 192.825 ;
        RECT 54.765 192.655 54.935 192.825 ;
        RECT 55.225 192.655 55.395 192.825 ;
        RECT 55.685 192.655 55.855 192.825 ;
        RECT 56.145 192.655 56.315 192.825 ;
        RECT 56.605 192.655 56.775 192.825 ;
        RECT 57.065 192.655 57.235 192.825 ;
        RECT 57.525 192.655 57.695 192.825 ;
        RECT 57.985 192.655 58.155 192.825 ;
        RECT 58.445 192.655 58.615 192.825 ;
        RECT 58.905 192.655 59.075 192.825 ;
        RECT 59.365 192.655 59.535 192.825 ;
        RECT 59.825 192.655 59.995 192.825 ;
        RECT 60.285 192.655 60.455 192.825 ;
        RECT 60.745 192.655 60.915 192.825 ;
        RECT 61.205 192.655 61.375 192.825 ;
        RECT 61.665 192.655 61.835 192.825 ;
        RECT 62.125 192.655 62.295 192.825 ;
        RECT 62.585 192.655 62.755 192.825 ;
        RECT 63.045 192.655 63.215 192.825 ;
        RECT 63.505 192.655 63.675 192.825 ;
        RECT 63.965 192.655 64.135 192.825 ;
        RECT 64.425 192.655 64.595 192.825 ;
        RECT 64.885 192.655 65.055 192.825 ;
        RECT 65.345 192.655 65.515 192.825 ;
        RECT 65.805 192.655 65.975 192.825 ;
        RECT 66.265 192.655 66.435 192.825 ;
        RECT 66.725 192.655 66.895 192.825 ;
        RECT 67.185 192.655 67.355 192.825 ;
        RECT 67.645 192.655 67.815 192.825 ;
        RECT 68.105 192.655 68.275 192.825 ;
        RECT 68.565 192.655 68.735 192.825 ;
        RECT 69.025 192.655 69.195 192.825 ;
        RECT 69.485 192.655 69.655 192.825 ;
        RECT 69.945 192.655 70.115 192.825 ;
        RECT 70.405 192.655 70.575 192.825 ;
        RECT 70.865 192.655 71.035 192.825 ;
        RECT 71.325 192.655 71.495 192.825 ;
        RECT 71.785 192.655 71.955 192.825 ;
        RECT 72.245 192.655 72.415 192.825 ;
        RECT 72.705 192.655 72.875 192.825 ;
        RECT 73.165 192.655 73.335 192.825 ;
        RECT 73.625 192.655 73.795 192.825 ;
        RECT 74.085 192.655 74.255 192.825 ;
        RECT 74.545 192.655 74.715 192.825 ;
        RECT 75.005 192.655 75.175 192.825 ;
        RECT 75.465 192.655 75.635 192.825 ;
        RECT 75.925 192.655 76.095 192.825 ;
        RECT 76.385 192.655 76.555 192.825 ;
        RECT 76.845 192.655 77.015 192.825 ;
        RECT 77.305 192.655 77.475 192.825 ;
        RECT 77.765 192.655 77.935 192.825 ;
        RECT 78.225 192.655 78.395 192.825 ;
        RECT 78.685 192.655 78.855 192.825 ;
        RECT 79.145 192.655 79.315 192.825 ;
        RECT 79.605 192.655 79.775 192.825 ;
        RECT 80.065 192.655 80.235 192.825 ;
        RECT 80.525 192.655 80.695 192.825 ;
        RECT 80.985 192.655 81.155 192.825 ;
        RECT 81.445 192.655 81.615 192.825 ;
        RECT 81.905 192.655 82.075 192.825 ;
        RECT 82.365 192.655 82.535 192.825 ;
        RECT 82.825 192.655 82.995 192.825 ;
        RECT 83.285 192.655 83.455 192.825 ;
        RECT 83.745 192.655 83.915 192.825 ;
        RECT 84.205 192.655 84.375 192.825 ;
        RECT 84.665 192.655 84.835 192.825 ;
        RECT 85.125 192.655 85.295 192.825 ;
        RECT 85.585 192.655 85.755 192.825 ;
        RECT 86.045 192.655 86.215 192.825 ;
        RECT 86.505 192.655 86.675 192.825 ;
        RECT 86.965 192.655 87.135 192.825 ;
        RECT 87.425 192.655 87.595 192.825 ;
        RECT 87.885 192.655 88.055 192.825 ;
        RECT 88.345 192.655 88.515 192.825 ;
        RECT 88.805 192.655 88.975 192.825 ;
        RECT 89.265 192.655 89.435 192.825 ;
        RECT 89.725 192.655 89.895 192.825 ;
        RECT 90.185 192.655 90.355 192.825 ;
        RECT 90.645 192.655 90.815 192.825 ;
        RECT 91.105 192.655 91.275 192.825 ;
        RECT 91.565 192.655 91.735 192.825 ;
        RECT 92.025 192.655 92.195 192.825 ;
        RECT 36.825 192.145 36.995 192.315 ;
        RECT 38.205 191.465 38.375 191.635 ;
        RECT 39.585 191.465 39.755 191.635 ;
        RECT 39.125 190.445 39.295 190.615 ;
        RECT 54.765 191.465 54.935 191.635 ;
        RECT 56.145 191.465 56.315 191.635 ;
        RECT 56.605 191.465 56.775 191.635 ;
        RECT 55.225 191.125 55.395 191.295 ;
        RECT 57.525 190.445 57.695 190.615 ;
        RECT 59.365 190.785 59.535 190.955 ;
        RECT 60.285 190.445 60.455 190.615 ;
        RECT 78.685 192.145 78.855 192.315 ;
        RECT 64.885 190.785 65.055 190.955 ;
        RECT 65.345 190.445 65.515 190.615 ;
        RECT 77.765 191.465 77.935 191.635 ;
        RECT 76.845 191.125 77.015 191.295 ;
        RECT 82.365 191.465 82.535 191.635 ;
        RECT 82.830 190.785 83.000 190.955 ;
        RECT 83.290 191.805 83.460 191.975 ;
        RECT 83.745 191.465 83.915 191.635 ;
        RECT 84.690 191.805 84.860 191.975 ;
        RECT 86.530 191.805 86.700 191.975 ;
        RECT 85.150 190.785 85.320 190.955 ;
        RECT 86.530 190.785 86.700 190.955 ;
        RECT 90.645 191.805 90.815 191.975 ;
        RECT 18.425 189.935 18.595 190.105 ;
        RECT 18.885 189.935 19.055 190.105 ;
        RECT 19.345 189.935 19.515 190.105 ;
        RECT 19.805 189.935 19.975 190.105 ;
        RECT 20.265 189.935 20.435 190.105 ;
        RECT 20.725 189.935 20.895 190.105 ;
        RECT 21.185 189.935 21.355 190.105 ;
        RECT 21.645 189.935 21.815 190.105 ;
        RECT 22.105 189.935 22.275 190.105 ;
        RECT 22.565 189.935 22.735 190.105 ;
        RECT 23.025 189.935 23.195 190.105 ;
        RECT 23.485 189.935 23.655 190.105 ;
        RECT 23.945 189.935 24.115 190.105 ;
        RECT 24.405 189.935 24.575 190.105 ;
        RECT 24.865 189.935 25.035 190.105 ;
        RECT 25.325 189.935 25.495 190.105 ;
        RECT 25.785 189.935 25.955 190.105 ;
        RECT 26.245 189.935 26.415 190.105 ;
        RECT 26.705 189.935 26.875 190.105 ;
        RECT 27.165 189.935 27.335 190.105 ;
        RECT 27.625 189.935 27.795 190.105 ;
        RECT 28.085 189.935 28.255 190.105 ;
        RECT 28.545 189.935 28.715 190.105 ;
        RECT 29.005 189.935 29.175 190.105 ;
        RECT 29.465 189.935 29.635 190.105 ;
        RECT 29.925 189.935 30.095 190.105 ;
        RECT 30.385 189.935 30.555 190.105 ;
        RECT 30.845 189.935 31.015 190.105 ;
        RECT 31.305 189.935 31.475 190.105 ;
        RECT 31.765 189.935 31.935 190.105 ;
        RECT 32.225 189.935 32.395 190.105 ;
        RECT 32.685 189.935 32.855 190.105 ;
        RECT 33.145 189.935 33.315 190.105 ;
        RECT 33.605 189.935 33.775 190.105 ;
        RECT 34.065 189.935 34.235 190.105 ;
        RECT 34.525 189.935 34.695 190.105 ;
        RECT 34.985 189.935 35.155 190.105 ;
        RECT 35.445 189.935 35.615 190.105 ;
        RECT 35.905 189.935 36.075 190.105 ;
        RECT 36.365 189.935 36.535 190.105 ;
        RECT 36.825 189.935 36.995 190.105 ;
        RECT 37.285 189.935 37.455 190.105 ;
        RECT 37.745 189.935 37.915 190.105 ;
        RECT 38.205 189.935 38.375 190.105 ;
        RECT 38.665 189.935 38.835 190.105 ;
        RECT 39.125 189.935 39.295 190.105 ;
        RECT 39.585 189.935 39.755 190.105 ;
        RECT 40.045 189.935 40.215 190.105 ;
        RECT 40.505 189.935 40.675 190.105 ;
        RECT 40.965 189.935 41.135 190.105 ;
        RECT 41.425 189.935 41.595 190.105 ;
        RECT 41.885 189.935 42.055 190.105 ;
        RECT 42.345 189.935 42.515 190.105 ;
        RECT 42.805 189.935 42.975 190.105 ;
        RECT 43.265 189.935 43.435 190.105 ;
        RECT 43.725 189.935 43.895 190.105 ;
        RECT 44.185 189.935 44.355 190.105 ;
        RECT 44.645 189.935 44.815 190.105 ;
        RECT 45.105 189.935 45.275 190.105 ;
        RECT 45.565 189.935 45.735 190.105 ;
        RECT 46.025 189.935 46.195 190.105 ;
        RECT 46.485 189.935 46.655 190.105 ;
        RECT 46.945 189.935 47.115 190.105 ;
        RECT 47.405 189.935 47.575 190.105 ;
        RECT 47.865 189.935 48.035 190.105 ;
        RECT 48.325 189.935 48.495 190.105 ;
        RECT 48.785 189.935 48.955 190.105 ;
        RECT 49.245 189.935 49.415 190.105 ;
        RECT 49.705 189.935 49.875 190.105 ;
        RECT 50.165 189.935 50.335 190.105 ;
        RECT 50.625 189.935 50.795 190.105 ;
        RECT 51.085 189.935 51.255 190.105 ;
        RECT 51.545 189.935 51.715 190.105 ;
        RECT 52.005 189.935 52.175 190.105 ;
        RECT 52.465 189.935 52.635 190.105 ;
        RECT 52.925 189.935 53.095 190.105 ;
        RECT 53.385 189.935 53.555 190.105 ;
        RECT 53.845 189.935 54.015 190.105 ;
        RECT 54.305 189.935 54.475 190.105 ;
        RECT 54.765 189.935 54.935 190.105 ;
        RECT 55.225 189.935 55.395 190.105 ;
        RECT 55.685 189.935 55.855 190.105 ;
        RECT 56.145 189.935 56.315 190.105 ;
        RECT 56.605 189.935 56.775 190.105 ;
        RECT 57.065 189.935 57.235 190.105 ;
        RECT 57.525 189.935 57.695 190.105 ;
        RECT 57.985 189.935 58.155 190.105 ;
        RECT 58.445 189.935 58.615 190.105 ;
        RECT 58.905 189.935 59.075 190.105 ;
        RECT 59.365 189.935 59.535 190.105 ;
        RECT 59.825 189.935 59.995 190.105 ;
        RECT 60.285 189.935 60.455 190.105 ;
        RECT 60.745 189.935 60.915 190.105 ;
        RECT 61.205 189.935 61.375 190.105 ;
        RECT 61.665 189.935 61.835 190.105 ;
        RECT 62.125 189.935 62.295 190.105 ;
        RECT 62.585 189.935 62.755 190.105 ;
        RECT 63.045 189.935 63.215 190.105 ;
        RECT 63.505 189.935 63.675 190.105 ;
        RECT 63.965 189.935 64.135 190.105 ;
        RECT 64.425 189.935 64.595 190.105 ;
        RECT 64.885 189.935 65.055 190.105 ;
        RECT 65.345 189.935 65.515 190.105 ;
        RECT 65.805 189.935 65.975 190.105 ;
        RECT 66.265 189.935 66.435 190.105 ;
        RECT 66.725 189.935 66.895 190.105 ;
        RECT 67.185 189.935 67.355 190.105 ;
        RECT 67.645 189.935 67.815 190.105 ;
        RECT 68.105 189.935 68.275 190.105 ;
        RECT 68.565 189.935 68.735 190.105 ;
        RECT 69.025 189.935 69.195 190.105 ;
        RECT 69.485 189.935 69.655 190.105 ;
        RECT 69.945 189.935 70.115 190.105 ;
        RECT 70.405 189.935 70.575 190.105 ;
        RECT 70.865 189.935 71.035 190.105 ;
        RECT 71.325 189.935 71.495 190.105 ;
        RECT 71.785 189.935 71.955 190.105 ;
        RECT 72.245 189.935 72.415 190.105 ;
        RECT 72.705 189.935 72.875 190.105 ;
        RECT 73.165 189.935 73.335 190.105 ;
        RECT 73.625 189.935 73.795 190.105 ;
        RECT 74.085 189.935 74.255 190.105 ;
        RECT 74.545 189.935 74.715 190.105 ;
        RECT 75.005 189.935 75.175 190.105 ;
        RECT 75.465 189.935 75.635 190.105 ;
        RECT 75.925 189.935 76.095 190.105 ;
        RECT 76.385 189.935 76.555 190.105 ;
        RECT 76.845 189.935 77.015 190.105 ;
        RECT 77.305 189.935 77.475 190.105 ;
        RECT 77.765 189.935 77.935 190.105 ;
        RECT 78.225 189.935 78.395 190.105 ;
        RECT 78.685 189.935 78.855 190.105 ;
        RECT 79.145 189.935 79.315 190.105 ;
        RECT 79.605 189.935 79.775 190.105 ;
        RECT 80.065 189.935 80.235 190.105 ;
        RECT 80.525 189.935 80.695 190.105 ;
        RECT 80.985 189.935 81.155 190.105 ;
        RECT 81.445 189.935 81.615 190.105 ;
        RECT 81.905 189.935 82.075 190.105 ;
        RECT 82.365 189.935 82.535 190.105 ;
        RECT 82.825 189.935 82.995 190.105 ;
        RECT 83.285 189.935 83.455 190.105 ;
        RECT 83.745 189.935 83.915 190.105 ;
        RECT 84.205 189.935 84.375 190.105 ;
        RECT 84.665 189.935 84.835 190.105 ;
        RECT 85.125 189.935 85.295 190.105 ;
        RECT 85.585 189.935 85.755 190.105 ;
        RECT 86.045 189.935 86.215 190.105 ;
        RECT 86.505 189.935 86.675 190.105 ;
        RECT 86.965 189.935 87.135 190.105 ;
        RECT 87.425 189.935 87.595 190.105 ;
        RECT 87.885 189.935 88.055 190.105 ;
        RECT 88.345 189.935 88.515 190.105 ;
        RECT 88.805 189.935 88.975 190.105 ;
        RECT 89.265 189.935 89.435 190.105 ;
        RECT 89.725 189.935 89.895 190.105 ;
        RECT 90.185 189.935 90.355 190.105 ;
        RECT 90.645 189.935 90.815 190.105 ;
        RECT 91.105 189.935 91.275 190.105 ;
        RECT 91.565 189.935 91.735 190.105 ;
        RECT 92.025 189.935 92.195 190.105 ;
        RECT 34.985 188.745 35.155 188.915 ;
        RECT 35.445 188.405 35.615 188.575 ;
        RECT 37.285 188.745 37.455 188.915 ;
        RECT 40.965 188.405 41.135 188.575 ;
        RECT 41.885 188.405 42.055 188.575 ;
        RECT 42.345 188.405 42.515 188.575 ;
        RECT 42.805 188.405 42.975 188.575 ;
        RECT 44.185 187.725 44.355 187.895 ;
        RECT 48.785 189.085 48.955 189.255 ;
        RECT 49.705 188.405 49.875 188.575 ;
        RECT 50.445 188.405 50.615 188.575 ;
        RECT 51.085 188.405 51.255 188.575 ;
        RECT 49.245 187.725 49.415 187.895 ;
        RECT 52.235 188.405 52.405 188.575 ;
        RECT 51.545 188.065 51.715 188.235 ;
        RECT 52.925 187.725 53.095 187.895 ;
        RECT 54.305 188.405 54.475 188.575 ;
        RECT 54.765 188.405 54.935 188.575 ;
        RECT 53.385 187.725 53.555 187.895 ;
        RECT 56.145 188.745 56.315 188.915 ;
        RECT 56.605 188.065 56.775 188.235 ;
        RECT 64.450 189.085 64.620 189.255 ;
        RECT 59.135 188.405 59.305 188.575 ;
        RECT 58.445 187.725 58.615 187.895 ;
        RECT 59.825 188.065 59.995 188.235 ;
        RECT 61.200 188.405 61.370 188.575 ;
        RECT 61.665 188.405 61.835 188.575 ;
        RECT 60.285 188.065 60.455 188.235 ;
        RECT 63.965 188.745 64.135 188.915 ;
        RECT 64.845 188.745 65.015 188.915 ;
        RECT 65.190 188.065 65.360 188.235 ;
        RECT 66.550 189.085 66.720 189.255 ;
        RECT 66.035 188.745 66.205 188.915 ;
        RECT 68.120 189.085 68.290 189.255 ;
        RECT 68.555 188.745 68.725 188.915 ;
        RECT 70.865 187.725 71.035 187.895 ;
        RECT 71.325 187.725 71.495 187.895 ;
        RECT 74.085 188.745 74.255 188.915 ;
        RECT 75.925 188.405 76.095 188.575 ;
        RECT 76.845 188.405 77.015 188.575 ;
        RECT 76.385 187.725 76.555 187.895 ;
        RECT 79.145 189.425 79.315 189.595 ;
        RECT 80.065 189.425 80.235 189.595 ;
        RECT 79.985 187.725 80.155 187.895 ;
        RECT 80.985 188.065 81.155 188.235 ;
        RECT 84.665 188.405 84.835 188.575 ;
        RECT 85.125 188.405 85.295 188.575 ;
        RECT 85.585 188.405 85.755 188.575 ;
        RECT 83.285 187.725 83.455 187.895 ;
        RECT 86.505 188.405 86.675 188.575 ;
        RECT 18.425 187.215 18.595 187.385 ;
        RECT 18.885 187.215 19.055 187.385 ;
        RECT 19.345 187.215 19.515 187.385 ;
        RECT 19.805 187.215 19.975 187.385 ;
        RECT 20.265 187.215 20.435 187.385 ;
        RECT 20.725 187.215 20.895 187.385 ;
        RECT 21.185 187.215 21.355 187.385 ;
        RECT 21.645 187.215 21.815 187.385 ;
        RECT 22.105 187.215 22.275 187.385 ;
        RECT 22.565 187.215 22.735 187.385 ;
        RECT 23.025 187.215 23.195 187.385 ;
        RECT 23.485 187.215 23.655 187.385 ;
        RECT 23.945 187.215 24.115 187.385 ;
        RECT 24.405 187.215 24.575 187.385 ;
        RECT 24.865 187.215 25.035 187.385 ;
        RECT 25.325 187.215 25.495 187.385 ;
        RECT 25.785 187.215 25.955 187.385 ;
        RECT 26.245 187.215 26.415 187.385 ;
        RECT 26.705 187.215 26.875 187.385 ;
        RECT 27.165 187.215 27.335 187.385 ;
        RECT 27.625 187.215 27.795 187.385 ;
        RECT 28.085 187.215 28.255 187.385 ;
        RECT 28.545 187.215 28.715 187.385 ;
        RECT 29.005 187.215 29.175 187.385 ;
        RECT 29.465 187.215 29.635 187.385 ;
        RECT 29.925 187.215 30.095 187.385 ;
        RECT 30.385 187.215 30.555 187.385 ;
        RECT 30.845 187.215 31.015 187.385 ;
        RECT 31.305 187.215 31.475 187.385 ;
        RECT 31.765 187.215 31.935 187.385 ;
        RECT 32.225 187.215 32.395 187.385 ;
        RECT 32.685 187.215 32.855 187.385 ;
        RECT 33.145 187.215 33.315 187.385 ;
        RECT 33.605 187.215 33.775 187.385 ;
        RECT 34.065 187.215 34.235 187.385 ;
        RECT 34.525 187.215 34.695 187.385 ;
        RECT 34.985 187.215 35.155 187.385 ;
        RECT 35.445 187.215 35.615 187.385 ;
        RECT 35.905 187.215 36.075 187.385 ;
        RECT 36.365 187.215 36.535 187.385 ;
        RECT 36.825 187.215 36.995 187.385 ;
        RECT 37.285 187.215 37.455 187.385 ;
        RECT 37.745 187.215 37.915 187.385 ;
        RECT 38.205 187.215 38.375 187.385 ;
        RECT 38.665 187.215 38.835 187.385 ;
        RECT 39.125 187.215 39.295 187.385 ;
        RECT 39.585 187.215 39.755 187.385 ;
        RECT 40.045 187.215 40.215 187.385 ;
        RECT 40.505 187.215 40.675 187.385 ;
        RECT 40.965 187.215 41.135 187.385 ;
        RECT 41.425 187.215 41.595 187.385 ;
        RECT 41.885 187.215 42.055 187.385 ;
        RECT 42.345 187.215 42.515 187.385 ;
        RECT 42.805 187.215 42.975 187.385 ;
        RECT 43.265 187.215 43.435 187.385 ;
        RECT 43.725 187.215 43.895 187.385 ;
        RECT 44.185 187.215 44.355 187.385 ;
        RECT 44.645 187.215 44.815 187.385 ;
        RECT 45.105 187.215 45.275 187.385 ;
        RECT 45.565 187.215 45.735 187.385 ;
        RECT 46.025 187.215 46.195 187.385 ;
        RECT 46.485 187.215 46.655 187.385 ;
        RECT 46.945 187.215 47.115 187.385 ;
        RECT 47.405 187.215 47.575 187.385 ;
        RECT 47.865 187.215 48.035 187.385 ;
        RECT 48.325 187.215 48.495 187.385 ;
        RECT 48.785 187.215 48.955 187.385 ;
        RECT 49.245 187.215 49.415 187.385 ;
        RECT 49.705 187.215 49.875 187.385 ;
        RECT 50.165 187.215 50.335 187.385 ;
        RECT 50.625 187.215 50.795 187.385 ;
        RECT 51.085 187.215 51.255 187.385 ;
        RECT 51.545 187.215 51.715 187.385 ;
        RECT 52.005 187.215 52.175 187.385 ;
        RECT 52.465 187.215 52.635 187.385 ;
        RECT 52.925 187.215 53.095 187.385 ;
        RECT 53.385 187.215 53.555 187.385 ;
        RECT 53.845 187.215 54.015 187.385 ;
        RECT 54.305 187.215 54.475 187.385 ;
        RECT 54.765 187.215 54.935 187.385 ;
        RECT 55.225 187.215 55.395 187.385 ;
        RECT 55.685 187.215 55.855 187.385 ;
        RECT 56.145 187.215 56.315 187.385 ;
        RECT 56.605 187.215 56.775 187.385 ;
        RECT 57.065 187.215 57.235 187.385 ;
        RECT 57.525 187.215 57.695 187.385 ;
        RECT 57.985 187.215 58.155 187.385 ;
        RECT 58.445 187.215 58.615 187.385 ;
        RECT 58.905 187.215 59.075 187.385 ;
        RECT 59.365 187.215 59.535 187.385 ;
        RECT 59.825 187.215 59.995 187.385 ;
        RECT 60.285 187.215 60.455 187.385 ;
        RECT 60.745 187.215 60.915 187.385 ;
        RECT 61.205 187.215 61.375 187.385 ;
        RECT 61.665 187.215 61.835 187.385 ;
        RECT 62.125 187.215 62.295 187.385 ;
        RECT 62.585 187.215 62.755 187.385 ;
        RECT 63.045 187.215 63.215 187.385 ;
        RECT 63.505 187.215 63.675 187.385 ;
        RECT 63.965 187.215 64.135 187.385 ;
        RECT 64.425 187.215 64.595 187.385 ;
        RECT 64.885 187.215 65.055 187.385 ;
        RECT 65.345 187.215 65.515 187.385 ;
        RECT 65.805 187.215 65.975 187.385 ;
        RECT 66.265 187.215 66.435 187.385 ;
        RECT 66.725 187.215 66.895 187.385 ;
        RECT 67.185 187.215 67.355 187.385 ;
        RECT 67.645 187.215 67.815 187.385 ;
        RECT 68.105 187.215 68.275 187.385 ;
        RECT 68.565 187.215 68.735 187.385 ;
        RECT 69.025 187.215 69.195 187.385 ;
        RECT 69.485 187.215 69.655 187.385 ;
        RECT 69.945 187.215 70.115 187.385 ;
        RECT 70.405 187.215 70.575 187.385 ;
        RECT 70.865 187.215 71.035 187.385 ;
        RECT 71.325 187.215 71.495 187.385 ;
        RECT 71.785 187.215 71.955 187.385 ;
        RECT 72.245 187.215 72.415 187.385 ;
        RECT 72.705 187.215 72.875 187.385 ;
        RECT 73.165 187.215 73.335 187.385 ;
        RECT 73.625 187.215 73.795 187.385 ;
        RECT 74.085 187.215 74.255 187.385 ;
        RECT 74.545 187.215 74.715 187.385 ;
        RECT 75.005 187.215 75.175 187.385 ;
        RECT 75.465 187.215 75.635 187.385 ;
        RECT 75.925 187.215 76.095 187.385 ;
        RECT 76.385 187.215 76.555 187.385 ;
        RECT 76.845 187.215 77.015 187.385 ;
        RECT 77.305 187.215 77.475 187.385 ;
        RECT 77.765 187.215 77.935 187.385 ;
        RECT 78.225 187.215 78.395 187.385 ;
        RECT 78.685 187.215 78.855 187.385 ;
        RECT 79.145 187.215 79.315 187.385 ;
        RECT 79.605 187.215 79.775 187.385 ;
        RECT 80.065 187.215 80.235 187.385 ;
        RECT 80.525 187.215 80.695 187.385 ;
        RECT 80.985 187.215 81.155 187.385 ;
        RECT 81.445 187.215 81.615 187.385 ;
        RECT 81.905 187.215 82.075 187.385 ;
        RECT 82.365 187.215 82.535 187.385 ;
        RECT 82.825 187.215 82.995 187.385 ;
        RECT 83.285 187.215 83.455 187.385 ;
        RECT 83.745 187.215 83.915 187.385 ;
        RECT 84.205 187.215 84.375 187.385 ;
        RECT 84.665 187.215 84.835 187.385 ;
        RECT 85.125 187.215 85.295 187.385 ;
        RECT 85.585 187.215 85.755 187.385 ;
        RECT 86.045 187.215 86.215 187.385 ;
        RECT 86.505 187.215 86.675 187.385 ;
        RECT 86.965 187.215 87.135 187.385 ;
        RECT 87.425 187.215 87.595 187.385 ;
        RECT 87.885 187.215 88.055 187.385 ;
        RECT 88.345 187.215 88.515 187.385 ;
        RECT 88.805 187.215 88.975 187.385 ;
        RECT 89.265 187.215 89.435 187.385 ;
        RECT 89.725 187.215 89.895 187.385 ;
        RECT 90.185 187.215 90.355 187.385 ;
        RECT 90.645 187.215 90.815 187.385 ;
        RECT 91.105 187.215 91.275 187.385 ;
        RECT 91.565 187.215 91.735 187.385 ;
        RECT 92.025 187.215 92.195 187.385 ;
        RECT 36.825 186.705 36.995 186.875 ;
        RECT 34.525 186.025 34.695 186.195 ;
        RECT 39.585 186.705 39.755 186.875 ;
        RECT 37.285 186.025 37.455 186.195 ;
        RECT 34.985 185.005 35.155 185.175 ;
        RECT 40.045 186.025 40.215 186.195 ;
        RECT 38.665 185.005 38.835 185.175 ;
        RECT 40.505 185.005 40.675 185.175 ;
        RECT 42.805 185.345 42.975 185.515 ;
        RECT 45.105 186.025 45.275 186.195 ;
        RECT 45.565 186.025 45.735 186.195 ;
        RECT 46.485 186.025 46.655 186.195 ;
        RECT 46.025 185.345 46.195 185.515 ;
        RECT 47.405 185.005 47.575 185.175 ;
        RECT 48.785 186.025 48.955 186.195 ;
        RECT 50.625 186.025 50.795 186.195 ;
        RECT 47.865 185.345 48.035 185.515 ;
        RECT 50.165 185.345 50.335 185.515 ;
        RECT 54.305 186.705 54.475 186.875 ;
        RECT 52.465 186.025 52.635 186.195 ;
        RECT 51.085 185.005 51.255 185.175 ;
        RECT 52.925 185.345 53.095 185.515 ;
        RECT 60.285 186.705 60.455 186.875 ;
        RECT 54.765 186.025 54.935 186.195 ;
        RECT 53.385 185.005 53.555 185.175 ;
        RECT 57.985 186.025 58.155 186.195 ;
        RECT 63.965 186.705 64.135 186.875 ;
        RECT 59.365 185.005 59.535 185.175 ;
        RECT 64.885 186.025 65.055 186.195 ;
        RECT 65.345 185.345 65.515 185.515 ;
        RECT 66.265 186.025 66.435 186.195 ;
        RECT 68.105 186.365 68.275 186.535 ;
        RECT 67.185 186.025 67.355 186.195 ;
        RECT 68.565 186.025 68.735 186.195 ;
        RECT 65.805 185.345 65.975 185.515 ;
        RECT 73.625 185.685 73.795 185.855 ;
        RECT 75.005 186.705 75.175 186.875 ;
        RECT 74.545 185.685 74.715 185.855 ;
        RECT 77.305 186.025 77.475 186.195 ;
        RECT 78.685 186.025 78.855 186.195 ;
        RECT 79.145 186.025 79.315 186.195 ;
        RECT 76.845 185.005 77.015 185.175 ;
        RECT 82.365 186.025 82.535 186.195 ;
        RECT 82.830 185.345 83.000 185.515 ;
        RECT 83.290 186.365 83.460 186.535 ;
        RECT 83.745 186.025 83.915 186.195 ;
        RECT 84.690 186.365 84.860 186.535 ;
        RECT 86.530 186.365 86.700 186.535 ;
        RECT 85.150 185.345 85.320 185.515 ;
        RECT 86.530 185.345 86.700 185.515 ;
        RECT 90.185 185.005 90.355 185.175 ;
        RECT 18.425 184.495 18.595 184.665 ;
        RECT 18.885 184.495 19.055 184.665 ;
        RECT 19.345 184.495 19.515 184.665 ;
        RECT 19.805 184.495 19.975 184.665 ;
        RECT 20.265 184.495 20.435 184.665 ;
        RECT 20.725 184.495 20.895 184.665 ;
        RECT 21.185 184.495 21.355 184.665 ;
        RECT 21.645 184.495 21.815 184.665 ;
        RECT 22.105 184.495 22.275 184.665 ;
        RECT 22.565 184.495 22.735 184.665 ;
        RECT 23.025 184.495 23.195 184.665 ;
        RECT 23.485 184.495 23.655 184.665 ;
        RECT 23.945 184.495 24.115 184.665 ;
        RECT 24.405 184.495 24.575 184.665 ;
        RECT 24.865 184.495 25.035 184.665 ;
        RECT 25.325 184.495 25.495 184.665 ;
        RECT 25.785 184.495 25.955 184.665 ;
        RECT 26.245 184.495 26.415 184.665 ;
        RECT 26.705 184.495 26.875 184.665 ;
        RECT 27.165 184.495 27.335 184.665 ;
        RECT 27.625 184.495 27.795 184.665 ;
        RECT 28.085 184.495 28.255 184.665 ;
        RECT 28.545 184.495 28.715 184.665 ;
        RECT 29.005 184.495 29.175 184.665 ;
        RECT 29.465 184.495 29.635 184.665 ;
        RECT 29.925 184.495 30.095 184.665 ;
        RECT 30.385 184.495 30.555 184.665 ;
        RECT 30.845 184.495 31.015 184.665 ;
        RECT 31.305 184.495 31.475 184.665 ;
        RECT 31.765 184.495 31.935 184.665 ;
        RECT 32.225 184.495 32.395 184.665 ;
        RECT 32.685 184.495 32.855 184.665 ;
        RECT 33.145 184.495 33.315 184.665 ;
        RECT 33.605 184.495 33.775 184.665 ;
        RECT 34.065 184.495 34.235 184.665 ;
        RECT 34.525 184.495 34.695 184.665 ;
        RECT 34.985 184.495 35.155 184.665 ;
        RECT 35.445 184.495 35.615 184.665 ;
        RECT 35.905 184.495 36.075 184.665 ;
        RECT 36.365 184.495 36.535 184.665 ;
        RECT 36.825 184.495 36.995 184.665 ;
        RECT 37.285 184.495 37.455 184.665 ;
        RECT 37.745 184.495 37.915 184.665 ;
        RECT 38.205 184.495 38.375 184.665 ;
        RECT 38.665 184.495 38.835 184.665 ;
        RECT 39.125 184.495 39.295 184.665 ;
        RECT 39.585 184.495 39.755 184.665 ;
        RECT 40.045 184.495 40.215 184.665 ;
        RECT 40.505 184.495 40.675 184.665 ;
        RECT 40.965 184.495 41.135 184.665 ;
        RECT 41.425 184.495 41.595 184.665 ;
        RECT 41.885 184.495 42.055 184.665 ;
        RECT 42.345 184.495 42.515 184.665 ;
        RECT 42.805 184.495 42.975 184.665 ;
        RECT 43.265 184.495 43.435 184.665 ;
        RECT 43.725 184.495 43.895 184.665 ;
        RECT 44.185 184.495 44.355 184.665 ;
        RECT 44.645 184.495 44.815 184.665 ;
        RECT 45.105 184.495 45.275 184.665 ;
        RECT 45.565 184.495 45.735 184.665 ;
        RECT 46.025 184.495 46.195 184.665 ;
        RECT 46.485 184.495 46.655 184.665 ;
        RECT 46.945 184.495 47.115 184.665 ;
        RECT 47.405 184.495 47.575 184.665 ;
        RECT 47.865 184.495 48.035 184.665 ;
        RECT 48.325 184.495 48.495 184.665 ;
        RECT 48.785 184.495 48.955 184.665 ;
        RECT 49.245 184.495 49.415 184.665 ;
        RECT 49.705 184.495 49.875 184.665 ;
        RECT 50.165 184.495 50.335 184.665 ;
        RECT 50.625 184.495 50.795 184.665 ;
        RECT 51.085 184.495 51.255 184.665 ;
        RECT 51.545 184.495 51.715 184.665 ;
        RECT 52.005 184.495 52.175 184.665 ;
        RECT 52.465 184.495 52.635 184.665 ;
        RECT 52.925 184.495 53.095 184.665 ;
        RECT 53.385 184.495 53.555 184.665 ;
        RECT 53.845 184.495 54.015 184.665 ;
        RECT 54.305 184.495 54.475 184.665 ;
        RECT 54.765 184.495 54.935 184.665 ;
        RECT 55.225 184.495 55.395 184.665 ;
        RECT 55.685 184.495 55.855 184.665 ;
        RECT 56.145 184.495 56.315 184.665 ;
        RECT 56.605 184.495 56.775 184.665 ;
        RECT 57.065 184.495 57.235 184.665 ;
        RECT 57.525 184.495 57.695 184.665 ;
        RECT 57.985 184.495 58.155 184.665 ;
        RECT 58.445 184.495 58.615 184.665 ;
        RECT 58.905 184.495 59.075 184.665 ;
        RECT 59.365 184.495 59.535 184.665 ;
        RECT 59.825 184.495 59.995 184.665 ;
        RECT 60.285 184.495 60.455 184.665 ;
        RECT 60.745 184.495 60.915 184.665 ;
        RECT 61.205 184.495 61.375 184.665 ;
        RECT 61.665 184.495 61.835 184.665 ;
        RECT 62.125 184.495 62.295 184.665 ;
        RECT 62.585 184.495 62.755 184.665 ;
        RECT 63.045 184.495 63.215 184.665 ;
        RECT 63.505 184.495 63.675 184.665 ;
        RECT 63.965 184.495 64.135 184.665 ;
        RECT 64.425 184.495 64.595 184.665 ;
        RECT 64.885 184.495 65.055 184.665 ;
        RECT 65.345 184.495 65.515 184.665 ;
        RECT 65.805 184.495 65.975 184.665 ;
        RECT 66.265 184.495 66.435 184.665 ;
        RECT 66.725 184.495 66.895 184.665 ;
        RECT 67.185 184.495 67.355 184.665 ;
        RECT 67.645 184.495 67.815 184.665 ;
        RECT 68.105 184.495 68.275 184.665 ;
        RECT 68.565 184.495 68.735 184.665 ;
        RECT 69.025 184.495 69.195 184.665 ;
        RECT 69.485 184.495 69.655 184.665 ;
        RECT 69.945 184.495 70.115 184.665 ;
        RECT 70.405 184.495 70.575 184.665 ;
        RECT 70.865 184.495 71.035 184.665 ;
        RECT 71.325 184.495 71.495 184.665 ;
        RECT 71.785 184.495 71.955 184.665 ;
        RECT 72.245 184.495 72.415 184.665 ;
        RECT 72.705 184.495 72.875 184.665 ;
        RECT 73.165 184.495 73.335 184.665 ;
        RECT 73.625 184.495 73.795 184.665 ;
        RECT 74.085 184.495 74.255 184.665 ;
        RECT 74.545 184.495 74.715 184.665 ;
        RECT 75.005 184.495 75.175 184.665 ;
        RECT 75.465 184.495 75.635 184.665 ;
        RECT 75.925 184.495 76.095 184.665 ;
        RECT 76.385 184.495 76.555 184.665 ;
        RECT 76.845 184.495 77.015 184.665 ;
        RECT 77.305 184.495 77.475 184.665 ;
        RECT 77.765 184.495 77.935 184.665 ;
        RECT 78.225 184.495 78.395 184.665 ;
        RECT 78.685 184.495 78.855 184.665 ;
        RECT 79.145 184.495 79.315 184.665 ;
        RECT 79.605 184.495 79.775 184.665 ;
        RECT 80.065 184.495 80.235 184.665 ;
        RECT 80.525 184.495 80.695 184.665 ;
        RECT 80.985 184.495 81.155 184.665 ;
        RECT 81.445 184.495 81.615 184.665 ;
        RECT 81.905 184.495 82.075 184.665 ;
        RECT 82.365 184.495 82.535 184.665 ;
        RECT 82.825 184.495 82.995 184.665 ;
        RECT 83.285 184.495 83.455 184.665 ;
        RECT 83.745 184.495 83.915 184.665 ;
        RECT 84.205 184.495 84.375 184.665 ;
        RECT 84.665 184.495 84.835 184.665 ;
        RECT 85.125 184.495 85.295 184.665 ;
        RECT 85.585 184.495 85.755 184.665 ;
        RECT 86.045 184.495 86.215 184.665 ;
        RECT 86.505 184.495 86.675 184.665 ;
        RECT 86.965 184.495 87.135 184.665 ;
        RECT 87.425 184.495 87.595 184.665 ;
        RECT 87.885 184.495 88.055 184.665 ;
        RECT 88.345 184.495 88.515 184.665 ;
        RECT 88.805 184.495 88.975 184.665 ;
        RECT 89.265 184.495 89.435 184.665 ;
        RECT 89.725 184.495 89.895 184.665 ;
        RECT 90.185 184.495 90.355 184.665 ;
        RECT 90.645 184.495 90.815 184.665 ;
        RECT 91.105 184.495 91.275 184.665 ;
        RECT 91.565 184.495 91.735 184.665 ;
        RECT 92.025 184.495 92.195 184.665 ;
        RECT 38.205 183.305 38.375 183.475 ;
        RECT 40.505 183.985 40.675 184.155 ;
        RECT 39.585 183.645 39.755 183.815 ;
        RECT 43.265 183.985 43.435 184.155 ;
        RECT 50.625 182.625 50.795 182.795 ;
        RECT 64.885 182.965 65.055 183.135 ;
        RECT 65.345 183.305 65.515 183.475 ;
        RECT 65.805 183.305 65.975 183.475 ;
        RECT 67.185 183.985 67.355 184.155 ;
        RECT 66.265 182.965 66.435 183.135 ;
        RECT 67.645 182.625 67.815 182.795 ;
        RECT 76.385 182.625 76.555 182.795 ;
        RECT 78.685 183.985 78.855 184.155 ;
        RECT 81.905 183.985 82.075 184.155 ;
        RECT 79.605 182.965 79.775 183.135 ;
        RECT 80.985 182.965 81.155 183.135 ;
        RECT 81.445 182.965 81.615 183.135 ;
        RECT 82.365 182.965 82.535 183.135 ;
        RECT 80.525 182.285 80.695 182.455 ;
        RECT 18.425 181.775 18.595 181.945 ;
        RECT 18.885 181.775 19.055 181.945 ;
        RECT 19.345 181.775 19.515 181.945 ;
        RECT 19.805 181.775 19.975 181.945 ;
        RECT 20.265 181.775 20.435 181.945 ;
        RECT 20.725 181.775 20.895 181.945 ;
        RECT 21.185 181.775 21.355 181.945 ;
        RECT 21.645 181.775 21.815 181.945 ;
        RECT 22.105 181.775 22.275 181.945 ;
        RECT 22.565 181.775 22.735 181.945 ;
        RECT 23.025 181.775 23.195 181.945 ;
        RECT 23.485 181.775 23.655 181.945 ;
        RECT 23.945 181.775 24.115 181.945 ;
        RECT 24.405 181.775 24.575 181.945 ;
        RECT 24.865 181.775 25.035 181.945 ;
        RECT 25.325 181.775 25.495 181.945 ;
        RECT 25.785 181.775 25.955 181.945 ;
        RECT 26.245 181.775 26.415 181.945 ;
        RECT 26.705 181.775 26.875 181.945 ;
        RECT 27.165 181.775 27.335 181.945 ;
        RECT 27.625 181.775 27.795 181.945 ;
        RECT 28.085 181.775 28.255 181.945 ;
        RECT 28.545 181.775 28.715 181.945 ;
        RECT 29.005 181.775 29.175 181.945 ;
        RECT 29.465 181.775 29.635 181.945 ;
        RECT 29.925 181.775 30.095 181.945 ;
        RECT 30.385 181.775 30.555 181.945 ;
        RECT 30.845 181.775 31.015 181.945 ;
        RECT 31.305 181.775 31.475 181.945 ;
        RECT 31.765 181.775 31.935 181.945 ;
        RECT 32.225 181.775 32.395 181.945 ;
        RECT 32.685 181.775 32.855 181.945 ;
        RECT 33.145 181.775 33.315 181.945 ;
        RECT 33.605 181.775 33.775 181.945 ;
        RECT 34.065 181.775 34.235 181.945 ;
        RECT 34.525 181.775 34.695 181.945 ;
        RECT 34.985 181.775 35.155 181.945 ;
        RECT 35.445 181.775 35.615 181.945 ;
        RECT 35.905 181.775 36.075 181.945 ;
        RECT 36.365 181.775 36.535 181.945 ;
        RECT 36.825 181.775 36.995 181.945 ;
        RECT 37.285 181.775 37.455 181.945 ;
        RECT 37.745 181.775 37.915 181.945 ;
        RECT 38.205 181.775 38.375 181.945 ;
        RECT 38.665 181.775 38.835 181.945 ;
        RECT 39.125 181.775 39.295 181.945 ;
        RECT 39.585 181.775 39.755 181.945 ;
        RECT 40.045 181.775 40.215 181.945 ;
        RECT 40.505 181.775 40.675 181.945 ;
        RECT 40.965 181.775 41.135 181.945 ;
        RECT 41.425 181.775 41.595 181.945 ;
        RECT 41.885 181.775 42.055 181.945 ;
        RECT 42.345 181.775 42.515 181.945 ;
        RECT 42.805 181.775 42.975 181.945 ;
        RECT 43.265 181.775 43.435 181.945 ;
        RECT 43.725 181.775 43.895 181.945 ;
        RECT 44.185 181.775 44.355 181.945 ;
        RECT 44.645 181.775 44.815 181.945 ;
        RECT 45.105 181.775 45.275 181.945 ;
        RECT 45.565 181.775 45.735 181.945 ;
        RECT 46.025 181.775 46.195 181.945 ;
        RECT 46.485 181.775 46.655 181.945 ;
        RECT 46.945 181.775 47.115 181.945 ;
        RECT 47.405 181.775 47.575 181.945 ;
        RECT 47.865 181.775 48.035 181.945 ;
        RECT 48.325 181.775 48.495 181.945 ;
        RECT 48.785 181.775 48.955 181.945 ;
        RECT 49.245 181.775 49.415 181.945 ;
        RECT 49.705 181.775 49.875 181.945 ;
        RECT 50.165 181.775 50.335 181.945 ;
        RECT 50.625 181.775 50.795 181.945 ;
        RECT 51.085 181.775 51.255 181.945 ;
        RECT 51.545 181.775 51.715 181.945 ;
        RECT 52.005 181.775 52.175 181.945 ;
        RECT 52.465 181.775 52.635 181.945 ;
        RECT 52.925 181.775 53.095 181.945 ;
        RECT 53.385 181.775 53.555 181.945 ;
        RECT 53.845 181.775 54.015 181.945 ;
        RECT 54.305 181.775 54.475 181.945 ;
        RECT 54.765 181.775 54.935 181.945 ;
        RECT 55.225 181.775 55.395 181.945 ;
        RECT 55.685 181.775 55.855 181.945 ;
        RECT 56.145 181.775 56.315 181.945 ;
        RECT 56.605 181.775 56.775 181.945 ;
        RECT 57.065 181.775 57.235 181.945 ;
        RECT 57.525 181.775 57.695 181.945 ;
        RECT 57.985 181.775 58.155 181.945 ;
        RECT 58.445 181.775 58.615 181.945 ;
        RECT 58.905 181.775 59.075 181.945 ;
        RECT 59.365 181.775 59.535 181.945 ;
        RECT 59.825 181.775 59.995 181.945 ;
        RECT 60.285 181.775 60.455 181.945 ;
        RECT 60.745 181.775 60.915 181.945 ;
        RECT 61.205 181.775 61.375 181.945 ;
        RECT 61.665 181.775 61.835 181.945 ;
        RECT 62.125 181.775 62.295 181.945 ;
        RECT 62.585 181.775 62.755 181.945 ;
        RECT 63.045 181.775 63.215 181.945 ;
        RECT 63.505 181.775 63.675 181.945 ;
        RECT 63.965 181.775 64.135 181.945 ;
        RECT 64.425 181.775 64.595 181.945 ;
        RECT 64.885 181.775 65.055 181.945 ;
        RECT 65.345 181.775 65.515 181.945 ;
        RECT 65.805 181.775 65.975 181.945 ;
        RECT 66.265 181.775 66.435 181.945 ;
        RECT 66.725 181.775 66.895 181.945 ;
        RECT 67.185 181.775 67.355 181.945 ;
        RECT 67.645 181.775 67.815 181.945 ;
        RECT 68.105 181.775 68.275 181.945 ;
        RECT 68.565 181.775 68.735 181.945 ;
        RECT 69.025 181.775 69.195 181.945 ;
        RECT 69.485 181.775 69.655 181.945 ;
        RECT 69.945 181.775 70.115 181.945 ;
        RECT 70.405 181.775 70.575 181.945 ;
        RECT 70.865 181.775 71.035 181.945 ;
        RECT 71.325 181.775 71.495 181.945 ;
        RECT 71.785 181.775 71.955 181.945 ;
        RECT 72.245 181.775 72.415 181.945 ;
        RECT 72.705 181.775 72.875 181.945 ;
        RECT 73.165 181.775 73.335 181.945 ;
        RECT 73.625 181.775 73.795 181.945 ;
        RECT 74.085 181.775 74.255 181.945 ;
        RECT 74.545 181.775 74.715 181.945 ;
        RECT 75.005 181.775 75.175 181.945 ;
        RECT 75.465 181.775 75.635 181.945 ;
        RECT 75.925 181.775 76.095 181.945 ;
        RECT 76.385 181.775 76.555 181.945 ;
        RECT 76.845 181.775 77.015 181.945 ;
        RECT 77.305 181.775 77.475 181.945 ;
        RECT 77.765 181.775 77.935 181.945 ;
        RECT 78.225 181.775 78.395 181.945 ;
        RECT 78.685 181.775 78.855 181.945 ;
        RECT 79.145 181.775 79.315 181.945 ;
        RECT 79.605 181.775 79.775 181.945 ;
        RECT 80.065 181.775 80.235 181.945 ;
        RECT 80.525 181.775 80.695 181.945 ;
        RECT 80.985 181.775 81.155 181.945 ;
        RECT 81.445 181.775 81.615 181.945 ;
        RECT 81.905 181.775 82.075 181.945 ;
        RECT 82.365 181.775 82.535 181.945 ;
        RECT 82.825 181.775 82.995 181.945 ;
        RECT 83.285 181.775 83.455 181.945 ;
        RECT 83.745 181.775 83.915 181.945 ;
        RECT 84.205 181.775 84.375 181.945 ;
        RECT 84.665 181.775 84.835 181.945 ;
        RECT 85.125 181.775 85.295 181.945 ;
        RECT 85.585 181.775 85.755 181.945 ;
        RECT 86.045 181.775 86.215 181.945 ;
        RECT 86.505 181.775 86.675 181.945 ;
        RECT 86.965 181.775 87.135 181.945 ;
        RECT 87.425 181.775 87.595 181.945 ;
        RECT 87.885 181.775 88.055 181.945 ;
        RECT 88.345 181.775 88.515 181.945 ;
        RECT 88.805 181.775 88.975 181.945 ;
        RECT 89.265 181.775 89.435 181.945 ;
        RECT 89.725 181.775 89.895 181.945 ;
        RECT 90.185 181.775 90.355 181.945 ;
        RECT 90.645 181.775 90.815 181.945 ;
        RECT 91.105 181.775 91.275 181.945 ;
        RECT 91.565 181.775 91.735 181.945 ;
        RECT 92.025 181.775 92.195 181.945 ;
        RECT 41.425 180.585 41.595 180.755 ;
        RECT 42.345 180.585 42.515 180.755 ;
        RECT 42.345 179.565 42.515 179.735 ;
        RECT 45.105 180.925 45.275 181.095 ;
        RECT 47.865 180.925 48.035 181.095 ;
        RECT 48.325 180.585 48.495 180.755 ;
        RECT 52.465 181.265 52.635 181.435 ;
        RECT 46.485 179.565 46.655 179.735 ;
        RECT 53.845 181.265 54.015 181.435 ;
        RECT 52.925 180.585 53.095 180.755 ;
        RECT 58.445 181.265 58.615 181.435 ;
        RECT 54.305 180.585 54.475 180.755 ;
        RECT 57.985 180.585 58.155 180.755 ;
        RECT 59.365 180.585 59.535 180.755 ;
        RECT 60.745 180.585 60.915 180.755 ;
        RECT 60.285 180.245 60.455 180.415 ;
        RECT 64.885 181.265 65.055 181.435 ;
        RECT 61.665 180.585 61.835 180.755 ;
        RECT 62.125 180.585 62.295 180.755 ;
        RECT 62.585 180.585 62.755 180.755 ;
        RECT 64.425 180.585 64.595 180.755 ;
        RECT 65.805 180.585 65.975 180.755 ;
        RECT 63.965 179.905 64.135 180.075 ;
        RECT 65.805 179.565 65.975 179.735 ;
        RECT 72.705 181.265 72.875 181.435 ;
        RECT 72.245 180.925 72.415 181.095 ;
        RECT 76.845 180.585 77.015 180.755 ;
        RECT 77.765 180.585 77.935 180.755 ;
        RECT 79.605 180.585 79.775 180.755 ;
        RECT 78.225 180.245 78.395 180.415 ;
        RECT 80.925 180.585 81.095 180.755 ;
        RECT 81.445 180.585 81.615 180.755 ;
        RECT 81.905 180.585 82.075 180.755 ;
        RECT 80.525 179.905 80.695 180.075 ;
        RECT 82.365 180.245 82.535 180.415 ;
        RECT 82.830 179.905 83.000 180.075 ;
        RECT 83.290 180.925 83.460 181.095 ;
        RECT 83.745 180.245 83.915 180.415 ;
        RECT 84.690 180.925 84.860 181.095 ;
        RECT 86.530 180.925 86.700 181.095 ;
        RECT 85.150 179.905 85.320 180.075 ;
        RECT 86.530 179.905 86.700 180.075 ;
        RECT 90.185 179.565 90.355 179.735 ;
        RECT 18.425 179.055 18.595 179.225 ;
        RECT 18.885 179.055 19.055 179.225 ;
        RECT 19.345 179.055 19.515 179.225 ;
        RECT 19.805 179.055 19.975 179.225 ;
        RECT 20.265 179.055 20.435 179.225 ;
        RECT 20.725 179.055 20.895 179.225 ;
        RECT 21.185 179.055 21.355 179.225 ;
        RECT 21.645 179.055 21.815 179.225 ;
        RECT 22.105 179.055 22.275 179.225 ;
        RECT 22.565 179.055 22.735 179.225 ;
        RECT 23.025 179.055 23.195 179.225 ;
        RECT 23.485 179.055 23.655 179.225 ;
        RECT 23.945 179.055 24.115 179.225 ;
        RECT 24.405 179.055 24.575 179.225 ;
        RECT 24.865 179.055 25.035 179.225 ;
        RECT 25.325 179.055 25.495 179.225 ;
        RECT 25.785 179.055 25.955 179.225 ;
        RECT 26.245 179.055 26.415 179.225 ;
        RECT 26.705 179.055 26.875 179.225 ;
        RECT 27.165 179.055 27.335 179.225 ;
        RECT 27.625 179.055 27.795 179.225 ;
        RECT 28.085 179.055 28.255 179.225 ;
        RECT 28.545 179.055 28.715 179.225 ;
        RECT 29.005 179.055 29.175 179.225 ;
        RECT 29.465 179.055 29.635 179.225 ;
        RECT 29.925 179.055 30.095 179.225 ;
        RECT 30.385 179.055 30.555 179.225 ;
        RECT 30.845 179.055 31.015 179.225 ;
        RECT 31.305 179.055 31.475 179.225 ;
        RECT 31.765 179.055 31.935 179.225 ;
        RECT 32.225 179.055 32.395 179.225 ;
        RECT 32.685 179.055 32.855 179.225 ;
        RECT 33.145 179.055 33.315 179.225 ;
        RECT 33.605 179.055 33.775 179.225 ;
        RECT 34.065 179.055 34.235 179.225 ;
        RECT 34.525 179.055 34.695 179.225 ;
        RECT 34.985 179.055 35.155 179.225 ;
        RECT 35.445 179.055 35.615 179.225 ;
        RECT 35.905 179.055 36.075 179.225 ;
        RECT 36.365 179.055 36.535 179.225 ;
        RECT 36.825 179.055 36.995 179.225 ;
        RECT 37.285 179.055 37.455 179.225 ;
        RECT 37.745 179.055 37.915 179.225 ;
        RECT 38.205 179.055 38.375 179.225 ;
        RECT 38.665 179.055 38.835 179.225 ;
        RECT 39.125 179.055 39.295 179.225 ;
        RECT 39.585 179.055 39.755 179.225 ;
        RECT 40.045 179.055 40.215 179.225 ;
        RECT 40.505 179.055 40.675 179.225 ;
        RECT 40.965 179.055 41.135 179.225 ;
        RECT 41.425 179.055 41.595 179.225 ;
        RECT 41.885 179.055 42.055 179.225 ;
        RECT 42.345 179.055 42.515 179.225 ;
        RECT 42.805 179.055 42.975 179.225 ;
        RECT 43.265 179.055 43.435 179.225 ;
        RECT 43.725 179.055 43.895 179.225 ;
        RECT 44.185 179.055 44.355 179.225 ;
        RECT 44.645 179.055 44.815 179.225 ;
        RECT 45.105 179.055 45.275 179.225 ;
        RECT 45.565 179.055 45.735 179.225 ;
        RECT 46.025 179.055 46.195 179.225 ;
        RECT 46.485 179.055 46.655 179.225 ;
        RECT 46.945 179.055 47.115 179.225 ;
        RECT 47.405 179.055 47.575 179.225 ;
        RECT 47.865 179.055 48.035 179.225 ;
        RECT 48.325 179.055 48.495 179.225 ;
        RECT 48.785 179.055 48.955 179.225 ;
        RECT 49.245 179.055 49.415 179.225 ;
        RECT 49.705 179.055 49.875 179.225 ;
        RECT 50.165 179.055 50.335 179.225 ;
        RECT 50.625 179.055 50.795 179.225 ;
        RECT 51.085 179.055 51.255 179.225 ;
        RECT 51.545 179.055 51.715 179.225 ;
        RECT 52.005 179.055 52.175 179.225 ;
        RECT 52.465 179.055 52.635 179.225 ;
        RECT 52.925 179.055 53.095 179.225 ;
        RECT 53.385 179.055 53.555 179.225 ;
        RECT 53.845 179.055 54.015 179.225 ;
        RECT 54.305 179.055 54.475 179.225 ;
        RECT 54.765 179.055 54.935 179.225 ;
        RECT 55.225 179.055 55.395 179.225 ;
        RECT 55.685 179.055 55.855 179.225 ;
        RECT 56.145 179.055 56.315 179.225 ;
        RECT 56.605 179.055 56.775 179.225 ;
        RECT 57.065 179.055 57.235 179.225 ;
        RECT 57.525 179.055 57.695 179.225 ;
        RECT 57.985 179.055 58.155 179.225 ;
        RECT 58.445 179.055 58.615 179.225 ;
        RECT 58.905 179.055 59.075 179.225 ;
        RECT 59.365 179.055 59.535 179.225 ;
        RECT 59.825 179.055 59.995 179.225 ;
        RECT 60.285 179.055 60.455 179.225 ;
        RECT 60.745 179.055 60.915 179.225 ;
        RECT 61.205 179.055 61.375 179.225 ;
        RECT 61.665 179.055 61.835 179.225 ;
        RECT 62.125 179.055 62.295 179.225 ;
        RECT 62.585 179.055 62.755 179.225 ;
        RECT 63.045 179.055 63.215 179.225 ;
        RECT 63.505 179.055 63.675 179.225 ;
        RECT 63.965 179.055 64.135 179.225 ;
        RECT 64.425 179.055 64.595 179.225 ;
        RECT 64.885 179.055 65.055 179.225 ;
        RECT 65.345 179.055 65.515 179.225 ;
        RECT 65.805 179.055 65.975 179.225 ;
        RECT 66.265 179.055 66.435 179.225 ;
        RECT 66.725 179.055 66.895 179.225 ;
        RECT 67.185 179.055 67.355 179.225 ;
        RECT 67.645 179.055 67.815 179.225 ;
        RECT 68.105 179.055 68.275 179.225 ;
        RECT 68.565 179.055 68.735 179.225 ;
        RECT 69.025 179.055 69.195 179.225 ;
        RECT 69.485 179.055 69.655 179.225 ;
        RECT 69.945 179.055 70.115 179.225 ;
        RECT 70.405 179.055 70.575 179.225 ;
        RECT 70.865 179.055 71.035 179.225 ;
        RECT 71.325 179.055 71.495 179.225 ;
        RECT 71.785 179.055 71.955 179.225 ;
        RECT 72.245 179.055 72.415 179.225 ;
        RECT 72.705 179.055 72.875 179.225 ;
        RECT 73.165 179.055 73.335 179.225 ;
        RECT 73.625 179.055 73.795 179.225 ;
        RECT 74.085 179.055 74.255 179.225 ;
        RECT 74.545 179.055 74.715 179.225 ;
        RECT 75.005 179.055 75.175 179.225 ;
        RECT 75.465 179.055 75.635 179.225 ;
        RECT 75.925 179.055 76.095 179.225 ;
        RECT 76.385 179.055 76.555 179.225 ;
        RECT 76.845 179.055 77.015 179.225 ;
        RECT 77.305 179.055 77.475 179.225 ;
        RECT 77.765 179.055 77.935 179.225 ;
        RECT 78.225 179.055 78.395 179.225 ;
        RECT 78.685 179.055 78.855 179.225 ;
        RECT 79.145 179.055 79.315 179.225 ;
        RECT 79.605 179.055 79.775 179.225 ;
        RECT 80.065 179.055 80.235 179.225 ;
        RECT 80.525 179.055 80.695 179.225 ;
        RECT 80.985 179.055 81.155 179.225 ;
        RECT 81.445 179.055 81.615 179.225 ;
        RECT 81.905 179.055 82.075 179.225 ;
        RECT 82.365 179.055 82.535 179.225 ;
        RECT 82.825 179.055 82.995 179.225 ;
        RECT 83.285 179.055 83.455 179.225 ;
        RECT 83.745 179.055 83.915 179.225 ;
        RECT 84.205 179.055 84.375 179.225 ;
        RECT 84.665 179.055 84.835 179.225 ;
        RECT 85.125 179.055 85.295 179.225 ;
        RECT 85.585 179.055 85.755 179.225 ;
        RECT 86.045 179.055 86.215 179.225 ;
        RECT 86.505 179.055 86.675 179.225 ;
        RECT 86.965 179.055 87.135 179.225 ;
        RECT 87.425 179.055 87.595 179.225 ;
        RECT 87.885 179.055 88.055 179.225 ;
        RECT 88.345 179.055 88.515 179.225 ;
        RECT 88.805 179.055 88.975 179.225 ;
        RECT 89.265 179.055 89.435 179.225 ;
        RECT 89.725 179.055 89.895 179.225 ;
        RECT 90.185 179.055 90.355 179.225 ;
        RECT 90.645 179.055 90.815 179.225 ;
        RECT 91.105 179.055 91.275 179.225 ;
        RECT 91.565 179.055 91.735 179.225 ;
        RECT 92.025 179.055 92.195 179.225 ;
        RECT 40.530 178.205 40.700 178.375 ;
        RECT 40.045 177.865 40.215 178.035 ;
        RECT 40.925 177.865 41.095 178.035 ;
        RECT 41.380 177.525 41.550 177.695 ;
        RECT 42.630 178.205 42.800 178.375 ;
        RECT 42.115 177.865 42.285 178.035 ;
        RECT 44.200 178.205 44.370 178.375 ;
        RECT 44.635 177.865 44.805 178.035 ;
        RECT 46.945 178.205 47.115 178.375 ;
        RECT 49.245 178.545 49.415 178.715 ;
        RECT 50.165 177.525 50.335 177.695 ;
        RECT 50.625 177.525 50.795 177.695 ;
        RECT 51.085 177.865 51.255 178.035 ;
        RECT 51.545 177.525 51.715 177.695 ;
        RECT 53.385 178.545 53.555 178.715 ;
        RECT 54.305 178.545 54.475 178.715 ;
        RECT 52.465 177.525 52.635 177.695 ;
        RECT 54.175 176.845 54.345 177.015 ;
        RECT 55.225 177.185 55.395 177.355 ;
        RECT 58.445 178.545 58.615 178.715 ;
        RECT 59.365 178.205 59.535 178.375 ;
        RECT 57.525 177.185 57.695 177.355 ;
        RECT 62.125 178.545 62.295 178.715 ;
        RECT 58.575 176.845 58.745 177.015 ;
        RECT 64.435 177.865 64.605 178.035 ;
        RECT 64.870 178.205 65.040 178.375 ;
        RECT 66.440 178.205 66.610 178.375 ;
        RECT 66.955 177.865 67.125 178.035 ;
        RECT 67.690 177.525 67.860 177.695 ;
        RECT 68.145 177.865 68.315 178.035 ;
        RECT 68.540 178.205 68.710 178.375 ;
        RECT 69.025 177.865 69.195 178.035 ;
        RECT 72.245 178.545 72.415 178.715 ;
        RECT 69.485 177.525 69.655 177.695 ;
        RECT 70.405 177.525 70.575 177.695 ;
        RECT 71.325 177.525 71.495 177.695 ;
        RECT 70.405 176.845 70.575 177.015 ;
        RECT 77.765 177.525 77.935 177.695 ;
        RECT 78.505 177.525 78.675 177.695 ;
        RECT 79.145 177.525 79.315 177.695 ;
        RECT 79.605 177.525 79.775 177.695 ;
        RECT 80.090 177.525 80.260 177.695 ;
        RECT 82.365 178.545 82.535 178.715 ;
        RECT 81.445 177.525 81.615 177.695 ;
        RECT 82.365 177.525 82.535 177.695 ;
        RECT 84.665 177.525 84.835 177.695 ;
        RECT 85.125 177.525 85.295 177.695 ;
        RECT 85.585 177.525 85.755 177.695 ;
        RECT 83.285 176.845 83.455 177.015 ;
        RECT 86.505 177.525 86.675 177.695 ;
        RECT 18.425 176.335 18.595 176.505 ;
        RECT 18.885 176.335 19.055 176.505 ;
        RECT 19.345 176.335 19.515 176.505 ;
        RECT 19.805 176.335 19.975 176.505 ;
        RECT 20.265 176.335 20.435 176.505 ;
        RECT 20.725 176.335 20.895 176.505 ;
        RECT 21.185 176.335 21.355 176.505 ;
        RECT 21.645 176.335 21.815 176.505 ;
        RECT 22.105 176.335 22.275 176.505 ;
        RECT 22.565 176.335 22.735 176.505 ;
        RECT 23.025 176.335 23.195 176.505 ;
        RECT 23.485 176.335 23.655 176.505 ;
        RECT 23.945 176.335 24.115 176.505 ;
        RECT 24.405 176.335 24.575 176.505 ;
        RECT 24.865 176.335 25.035 176.505 ;
        RECT 25.325 176.335 25.495 176.505 ;
        RECT 25.785 176.335 25.955 176.505 ;
        RECT 26.245 176.335 26.415 176.505 ;
        RECT 26.705 176.335 26.875 176.505 ;
        RECT 27.165 176.335 27.335 176.505 ;
        RECT 27.625 176.335 27.795 176.505 ;
        RECT 28.085 176.335 28.255 176.505 ;
        RECT 28.545 176.335 28.715 176.505 ;
        RECT 29.005 176.335 29.175 176.505 ;
        RECT 29.465 176.335 29.635 176.505 ;
        RECT 29.925 176.335 30.095 176.505 ;
        RECT 30.385 176.335 30.555 176.505 ;
        RECT 30.845 176.335 31.015 176.505 ;
        RECT 31.305 176.335 31.475 176.505 ;
        RECT 31.765 176.335 31.935 176.505 ;
        RECT 32.225 176.335 32.395 176.505 ;
        RECT 32.685 176.335 32.855 176.505 ;
        RECT 33.145 176.335 33.315 176.505 ;
        RECT 33.605 176.335 33.775 176.505 ;
        RECT 34.065 176.335 34.235 176.505 ;
        RECT 34.525 176.335 34.695 176.505 ;
        RECT 34.985 176.335 35.155 176.505 ;
        RECT 35.445 176.335 35.615 176.505 ;
        RECT 35.905 176.335 36.075 176.505 ;
        RECT 36.365 176.335 36.535 176.505 ;
        RECT 36.825 176.335 36.995 176.505 ;
        RECT 37.285 176.335 37.455 176.505 ;
        RECT 37.745 176.335 37.915 176.505 ;
        RECT 38.205 176.335 38.375 176.505 ;
        RECT 38.665 176.335 38.835 176.505 ;
        RECT 39.125 176.335 39.295 176.505 ;
        RECT 39.585 176.335 39.755 176.505 ;
        RECT 40.045 176.335 40.215 176.505 ;
        RECT 40.505 176.335 40.675 176.505 ;
        RECT 40.965 176.335 41.135 176.505 ;
        RECT 41.425 176.335 41.595 176.505 ;
        RECT 41.885 176.335 42.055 176.505 ;
        RECT 42.345 176.335 42.515 176.505 ;
        RECT 42.805 176.335 42.975 176.505 ;
        RECT 43.265 176.335 43.435 176.505 ;
        RECT 43.725 176.335 43.895 176.505 ;
        RECT 44.185 176.335 44.355 176.505 ;
        RECT 44.645 176.335 44.815 176.505 ;
        RECT 45.105 176.335 45.275 176.505 ;
        RECT 45.565 176.335 45.735 176.505 ;
        RECT 46.025 176.335 46.195 176.505 ;
        RECT 46.485 176.335 46.655 176.505 ;
        RECT 46.945 176.335 47.115 176.505 ;
        RECT 47.405 176.335 47.575 176.505 ;
        RECT 47.865 176.335 48.035 176.505 ;
        RECT 48.325 176.335 48.495 176.505 ;
        RECT 48.785 176.335 48.955 176.505 ;
        RECT 49.245 176.335 49.415 176.505 ;
        RECT 49.705 176.335 49.875 176.505 ;
        RECT 50.165 176.335 50.335 176.505 ;
        RECT 50.625 176.335 50.795 176.505 ;
        RECT 51.085 176.335 51.255 176.505 ;
        RECT 51.545 176.335 51.715 176.505 ;
        RECT 52.005 176.335 52.175 176.505 ;
        RECT 52.465 176.335 52.635 176.505 ;
        RECT 52.925 176.335 53.095 176.505 ;
        RECT 53.385 176.335 53.555 176.505 ;
        RECT 53.845 176.335 54.015 176.505 ;
        RECT 54.305 176.335 54.475 176.505 ;
        RECT 54.765 176.335 54.935 176.505 ;
        RECT 55.225 176.335 55.395 176.505 ;
        RECT 55.685 176.335 55.855 176.505 ;
        RECT 56.145 176.335 56.315 176.505 ;
        RECT 56.605 176.335 56.775 176.505 ;
        RECT 57.065 176.335 57.235 176.505 ;
        RECT 57.525 176.335 57.695 176.505 ;
        RECT 57.985 176.335 58.155 176.505 ;
        RECT 58.445 176.335 58.615 176.505 ;
        RECT 58.905 176.335 59.075 176.505 ;
        RECT 59.365 176.335 59.535 176.505 ;
        RECT 59.825 176.335 59.995 176.505 ;
        RECT 60.285 176.335 60.455 176.505 ;
        RECT 60.745 176.335 60.915 176.505 ;
        RECT 61.205 176.335 61.375 176.505 ;
        RECT 61.665 176.335 61.835 176.505 ;
        RECT 62.125 176.335 62.295 176.505 ;
        RECT 62.585 176.335 62.755 176.505 ;
        RECT 63.045 176.335 63.215 176.505 ;
        RECT 63.505 176.335 63.675 176.505 ;
        RECT 63.965 176.335 64.135 176.505 ;
        RECT 64.425 176.335 64.595 176.505 ;
        RECT 64.885 176.335 65.055 176.505 ;
        RECT 65.345 176.335 65.515 176.505 ;
        RECT 65.805 176.335 65.975 176.505 ;
        RECT 66.265 176.335 66.435 176.505 ;
        RECT 66.725 176.335 66.895 176.505 ;
        RECT 67.185 176.335 67.355 176.505 ;
        RECT 67.645 176.335 67.815 176.505 ;
        RECT 68.105 176.335 68.275 176.505 ;
        RECT 68.565 176.335 68.735 176.505 ;
        RECT 69.025 176.335 69.195 176.505 ;
        RECT 69.485 176.335 69.655 176.505 ;
        RECT 69.945 176.335 70.115 176.505 ;
        RECT 70.405 176.335 70.575 176.505 ;
        RECT 70.865 176.335 71.035 176.505 ;
        RECT 71.325 176.335 71.495 176.505 ;
        RECT 71.785 176.335 71.955 176.505 ;
        RECT 72.245 176.335 72.415 176.505 ;
        RECT 72.705 176.335 72.875 176.505 ;
        RECT 73.165 176.335 73.335 176.505 ;
        RECT 73.625 176.335 73.795 176.505 ;
        RECT 74.085 176.335 74.255 176.505 ;
        RECT 74.545 176.335 74.715 176.505 ;
        RECT 75.005 176.335 75.175 176.505 ;
        RECT 75.465 176.335 75.635 176.505 ;
        RECT 75.925 176.335 76.095 176.505 ;
        RECT 76.385 176.335 76.555 176.505 ;
        RECT 76.845 176.335 77.015 176.505 ;
        RECT 77.305 176.335 77.475 176.505 ;
        RECT 77.765 176.335 77.935 176.505 ;
        RECT 78.225 176.335 78.395 176.505 ;
        RECT 78.685 176.335 78.855 176.505 ;
        RECT 79.145 176.335 79.315 176.505 ;
        RECT 79.605 176.335 79.775 176.505 ;
        RECT 80.065 176.335 80.235 176.505 ;
        RECT 80.525 176.335 80.695 176.505 ;
        RECT 80.985 176.335 81.155 176.505 ;
        RECT 81.445 176.335 81.615 176.505 ;
        RECT 81.905 176.335 82.075 176.505 ;
        RECT 82.365 176.335 82.535 176.505 ;
        RECT 82.825 176.335 82.995 176.505 ;
        RECT 83.285 176.335 83.455 176.505 ;
        RECT 83.745 176.335 83.915 176.505 ;
        RECT 84.205 176.335 84.375 176.505 ;
        RECT 84.665 176.335 84.835 176.505 ;
        RECT 85.125 176.335 85.295 176.505 ;
        RECT 85.585 176.335 85.755 176.505 ;
        RECT 86.045 176.335 86.215 176.505 ;
        RECT 86.505 176.335 86.675 176.505 ;
        RECT 86.965 176.335 87.135 176.505 ;
        RECT 87.425 176.335 87.595 176.505 ;
        RECT 87.885 176.335 88.055 176.505 ;
        RECT 88.345 176.335 88.515 176.505 ;
        RECT 88.805 176.335 88.975 176.505 ;
        RECT 89.265 176.335 89.435 176.505 ;
        RECT 89.725 176.335 89.895 176.505 ;
        RECT 90.185 176.335 90.355 176.505 ;
        RECT 90.645 176.335 90.815 176.505 ;
        RECT 91.105 176.335 91.275 176.505 ;
        RECT 91.565 176.335 91.735 176.505 ;
        RECT 92.025 176.335 92.195 176.505 ;
        RECT 34.525 174.125 34.695 174.295 ;
        RECT 36.835 174.805 37.005 174.975 ;
        RECT 37.270 174.465 37.440 174.635 ;
        RECT 39.355 174.805 39.525 174.975 ;
        RECT 38.840 174.465 39.010 174.635 ;
        RECT 40.145 175.145 40.315 175.315 ;
        RECT 40.545 174.805 40.715 174.975 ;
        RECT 41.425 175.145 41.595 175.315 ;
        RECT 41.885 175.145 42.055 175.315 ;
        RECT 42.805 175.145 42.975 175.315 ;
        RECT 40.940 174.465 41.110 174.635 ;
        RECT 42.345 174.805 42.515 174.975 ;
        RECT 46.485 175.145 46.655 175.315 ;
        RECT 45.565 174.805 45.735 174.975 ;
        RECT 47.405 175.145 47.575 175.315 ;
        RECT 47.865 174.805 48.035 174.975 ;
        RECT 46.945 174.465 47.115 174.635 ;
        RECT 49.705 175.825 49.875 175.995 ;
        RECT 48.785 175.145 48.955 175.315 ;
        RECT 49.245 175.145 49.415 175.315 ;
        RECT 51.085 175.145 51.255 175.315 ;
        RECT 52.005 175.485 52.175 175.655 ;
        RECT 53.845 175.825 54.015 175.995 ;
        RECT 52.465 175.145 52.635 175.315 ;
        RECT 53.385 175.145 53.555 175.315 ;
        RECT 51.085 174.465 51.255 174.635 ;
        RECT 66.725 175.485 66.895 175.655 ;
        RECT 60.285 174.125 60.455 174.295 ;
        RECT 70.865 174.805 71.035 174.975 ;
        RECT 71.325 174.805 71.495 174.975 ;
        RECT 71.780 175.145 71.950 175.315 ;
        RECT 72.245 175.145 72.415 175.315 ;
        RECT 73.165 174.125 73.335 174.295 ;
        RECT 73.625 175.825 73.795 175.995 ;
        RECT 75.005 175.145 75.175 175.315 ;
        RECT 75.465 175.145 75.635 175.315 ;
        RECT 77.305 175.145 77.475 175.315 ;
        RECT 79.145 175.485 79.315 175.655 ;
        RECT 78.225 175.145 78.395 175.315 ;
        RECT 74.545 174.125 74.715 174.295 ;
        RECT 82.365 175.145 82.535 175.315 ;
        RECT 82.830 174.465 83.000 174.635 ;
        RECT 83.290 175.485 83.460 175.655 ;
        RECT 83.745 175.145 83.915 175.315 ;
        RECT 84.690 175.485 84.860 175.655 ;
        RECT 86.530 175.485 86.700 175.655 ;
        RECT 85.150 174.465 85.320 174.635 ;
        RECT 86.530 174.465 86.700 174.635 ;
        RECT 90.185 174.125 90.355 174.295 ;
        RECT 18.425 173.615 18.595 173.785 ;
        RECT 18.885 173.615 19.055 173.785 ;
        RECT 19.345 173.615 19.515 173.785 ;
        RECT 19.805 173.615 19.975 173.785 ;
        RECT 20.265 173.615 20.435 173.785 ;
        RECT 20.725 173.615 20.895 173.785 ;
        RECT 21.185 173.615 21.355 173.785 ;
        RECT 21.645 173.615 21.815 173.785 ;
        RECT 22.105 173.615 22.275 173.785 ;
        RECT 22.565 173.615 22.735 173.785 ;
        RECT 23.025 173.615 23.195 173.785 ;
        RECT 23.485 173.615 23.655 173.785 ;
        RECT 23.945 173.615 24.115 173.785 ;
        RECT 24.405 173.615 24.575 173.785 ;
        RECT 24.865 173.615 25.035 173.785 ;
        RECT 25.325 173.615 25.495 173.785 ;
        RECT 25.785 173.615 25.955 173.785 ;
        RECT 26.245 173.615 26.415 173.785 ;
        RECT 26.705 173.615 26.875 173.785 ;
        RECT 27.165 173.615 27.335 173.785 ;
        RECT 27.625 173.615 27.795 173.785 ;
        RECT 28.085 173.615 28.255 173.785 ;
        RECT 28.545 173.615 28.715 173.785 ;
        RECT 29.005 173.615 29.175 173.785 ;
        RECT 29.465 173.615 29.635 173.785 ;
        RECT 29.925 173.615 30.095 173.785 ;
        RECT 30.385 173.615 30.555 173.785 ;
        RECT 30.845 173.615 31.015 173.785 ;
        RECT 31.305 173.615 31.475 173.785 ;
        RECT 31.765 173.615 31.935 173.785 ;
        RECT 32.225 173.615 32.395 173.785 ;
        RECT 32.685 173.615 32.855 173.785 ;
        RECT 33.145 173.615 33.315 173.785 ;
        RECT 33.605 173.615 33.775 173.785 ;
        RECT 34.065 173.615 34.235 173.785 ;
        RECT 34.525 173.615 34.695 173.785 ;
        RECT 34.985 173.615 35.155 173.785 ;
        RECT 35.445 173.615 35.615 173.785 ;
        RECT 35.905 173.615 36.075 173.785 ;
        RECT 36.365 173.615 36.535 173.785 ;
        RECT 36.825 173.615 36.995 173.785 ;
        RECT 37.285 173.615 37.455 173.785 ;
        RECT 37.745 173.615 37.915 173.785 ;
        RECT 38.205 173.615 38.375 173.785 ;
        RECT 38.665 173.615 38.835 173.785 ;
        RECT 39.125 173.615 39.295 173.785 ;
        RECT 39.585 173.615 39.755 173.785 ;
        RECT 40.045 173.615 40.215 173.785 ;
        RECT 40.505 173.615 40.675 173.785 ;
        RECT 40.965 173.615 41.135 173.785 ;
        RECT 41.425 173.615 41.595 173.785 ;
        RECT 41.885 173.615 42.055 173.785 ;
        RECT 42.345 173.615 42.515 173.785 ;
        RECT 42.805 173.615 42.975 173.785 ;
        RECT 43.265 173.615 43.435 173.785 ;
        RECT 43.725 173.615 43.895 173.785 ;
        RECT 44.185 173.615 44.355 173.785 ;
        RECT 44.645 173.615 44.815 173.785 ;
        RECT 45.105 173.615 45.275 173.785 ;
        RECT 45.565 173.615 45.735 173.785 ;
        RECT 46.025 173.615 46.195 173.785 ;
        RECT 46.485 173.615 46.655 173.785 ;
        RECT 46.945 173.615 47.115 173.785 ;
        RECT 47.405 173.615 47.575 173.785 ;
        RECT 47.865 173.615 48.035 173.785 ;
        RECT 48.325 173.615 48.495 173.785 ;
        RECT 48.785 173.615 48.955 173.785 ;
        RECT 49.245 173.615 49.415 173.785 ;
        RECT 49.705 173.615 49.875 173.785 ;
        RECT 50.165 173.615 50.335 173.785 ;
        RECT 50.625 173.615 50.795 173.785 ;
        RECT 51.085 173.615 51.255 173.785 ;
        RECT 51.545 173.615 51.715 173.785 ;
        RECT 52.005 173.615 52.175 173.785 ;
        RECT 52.465 173.615 52.635 173.785 ;
        RECT 52.925 173.615 53.095 173.785 ;
        RECT 53.385 173.615 53.555 173.785 ;
        RECT 53.845 173.615 54.015 173.785 ;
        RECT 54.305 173.615 54.475 173.785 ;
        RECT 54.765 173.615 54.935 173.785 ;
        RECT 55.225 173.615 55.395 173.785 ;
        RECT 55.685 173.615 55.855 173.785 ;
        RECT 56.145 173.615 56.315 173.785 ;
        RECT 56.605 173.615 56.775 173.785 ;
        RECT 57.065 173.615 57.235 173.785 ;
        RECT 57.525 173.615 57.695 173.785 ;
        RECT 57.985 173.615 58.155 173.785 ;
        RECT 58.445 173.615 58.615 173.785 ;
        RECT 58.905 173.615 59.075 173.785 ;
        RECT 59.365 173.615 59.535 173.785 ;
        RECT 59.825 173.615 59.995 173.785 ;
        RECT 60.285 173.615 60.455 173.785 ;
        RECT 60.745 173.615 60.915 173.785 ;
        RECT 61.205 173.615 61.375 173.785 ;
        RECT 61.665 173.615 61.835 173.785 ;
        RECT 62.125 173.615 62.295 173.785 ;
        RECT 62.585 173.615 62.755 173.785 ;
        RECT 63.045 173.615 63.215 173.785 ;
        RECT 63.505 173.615 63.675 173.785 ;
        RECT 63.965 173.615 64.135 173.785 ;
        RECT 64.425 173.615 64.595 173.785 ;
        RECT 64.885 173.615 65.055 173.785 ;
        RECT 65.345 173.615 65.515 173.785 ;
        RECT 65.805 173.615 65.975 173.785 ;
        RECT 66.265 173.615 66.435 173.785 ;
        RECT 66.725 173.615 66.895 173.785 ;
        RECT 67.185 173.615 67.355 173.785 ;
        RECT 67.645 173.615 67.815 173.785 ;
        RECT 68.105 173.615 68.275 173.785 ;
        RECT 68.565 173.615 68.735 173.785 ;
        RECT 69.025 173.615 69.195 173.785 ;
        RECT 69.485 173.615 69.655 173.785 ;
        RECT 69.945 173.615 70.115 173.785 ;
        RECT 70.405 173.615 70.575 173.785 ;
        RECT 70.865 173.615 71.035 173.785 ;
        RECT 71.325 173.615 71.495 173.785 ;
        RECT 71.785 173.615 71.955 173.785 ;
        RECT 72.245 173.615 72.415 173.785 ;
        RECT 72.705 173.615 72.875 173.785 ;
        RECT 73.165 173.615 73.335 173.785 ;
        RECT 73.625 173.615 73.795 173.785 ;
        RECT 74.085 173.615 74.255 173.785 ;
        RECT 74.545 173.615 74.715 173.785 ;
        RECT 75.005 173.615 75.175 173.785 ;
        RECT 75.465 173.615 75.635 173.785 ;
        RECT 75.925 173.615 76.095 173.785 ;
        RECT 76.385 173.615 76.555 173.785 ;
        RECT 76.845 173.615 77.015 173.785 ;
        RECT 77.305 173.615 77.475 173.785 ;
        RECT 77.765 173.615 77.935 173.785 ;
        RECT 78.225 173.615 78.395 173.785 ;
        RECT 78.685 173.615 78.855 173.785 ;
        RECT 79.145 173.615 79.315 173.785 ;
        RECT 79.605 173.615 79.775 173.785 ;
        RECT 80.065 173.615 80.235 173.785 ;
        RECT 80.525 173.615 80.695 173.785 ;
        RECT 80.985 173.615 81.155 173.785 ;
        RECT 81.445 173.615 81.615 173.785 ;
        RECT 81.905 173.615 82.075 173.785 ;
        RECT 82.365 173.615 82.535 173.785 ;
        RECT 82.825 173.615 82.995 173.785 ;
        RECT 83.285 173.615 83.455 173.785 ;
        RECT 83.745 173.615 83.915 173.785 ;
        RECT 84.205 173.615 84.375 173.785 ;
        RECT 84.665 173.615 84.835 173.785 ;
        RECT 85.125 173.615 85.295 173.785 ;
        RECT 85.585 173.615 85.755 173.785 ;
        RECT 86.045 173.615 86.215 173.785 ;
        RECT 86.505 173.615 86.675 173.785 ;
        RECT 86.965 173.615 87.135 173.785 ;
        RECT 87.425 173.615 87.595 173.785 ;
        RECT 87.885 173.615 88.055 173.785 ;
        RECT 88.345 173.615 88.515 173.785 ;
        RECT 88.805 173.615 88.975 173.785 ;
        RECT 89.265 173.615 89.435 173.785 ;
        RECT 89.725 173.615 89.895 173.785 ;
        RECT 90.185 173.615 90.355 173.785 ;
        RECT 90.645 173.615 90.815 173.785 ;
        RECT 91.105 173.615 91.275 173.785 ;
        RECT 91.565 173.615 91.735 173.785 ;
        RECT 92.025 173.615 92.195 173.785 ;
        RECT 38.205 172.085 38.375 172.255 ;
        RECT 41.425 171.405 41.595 171.575 ;
        RECT 46.485 173.105 46.655 173.275 ;
        RECT 45.105 172.085 45.275 172.255 ;
        RECT 45.565 171.405 45.735 171.575 ;
        RECT 46.485 172.085 46.655 172.255 ;
        RECT 51.085 172.085 51.255 172.255 ;
        RECT 54.305 172.425 54.475 172.595 ;
        RECT 52.005 172.085 52.175 172.255 ;
        RECT 52.465 172.085 52.635 172.255 ;
        RECT 53.385 172.085 53.555 172.255 ;
        RECT 52.005 171.405 52.175 171.575 ;
        RECT 55.685 171.745 55.855 171.915 ;
        RECT 58.315 172.085 58.485 172.255 ;
        RECT 56.605 171.405 56.775 171.575 ;
        RECT 59.825 172.085 59.995 172.255 ;
        RECT 58.905 171.745 59.075 171.915 ;
        RECT 59.365 171.745 59.535 171.915 ;
        RECT 62.585 172.765 62.755 172.935 ;
        RECT 61.205 172.085 61.375 172.255 ;
        RECT 62.125 172.085 62.295 172.255 ;
        RECT 60.745 171.405 60.915 171.575 ;
        RECT 61.665 171.745 61.835 171.915 ;
        RECT 64.895 172.425 65.065 172.595 ;
        RECT 65.330 172.765 65.500 172.935 ;
        RECT 66.900 172.765 67.070 172.935 ;
        RECT 67.415 172.425 67.585 172.595 ;
        RECT 68.150 171.745 68.320 171.915 ;
        RECT 68.605 172.425 68.775 172.595 ;
        RECT 69.000 172.765 69.170 172.935 ;
        RECT 69.485 172.085 69.655 172.255 ;
        RECT 74.545 173.105 74.715 173.275 ;
        RECT 75.465 173.105 75.635 173.275 ;
        RECT 76.385 173.105 76.555 173.275 ;
        RECT 73.165 172.085 73.335 172.255 ;
        RECT 73.625 172.085 73.795 172.255 ;
        RECT 74.545 171.745 74.715 171.915 ;
        RECT 76.305 171.405 76.475 171.575 ;
        RECT 77.305 171.745 77.475 171.915 ;
        RECT 81.905 173.105 82.075 173.275 ;
        RECT 79.145 172.425 79.315 172.595 ;
        RECT 80.065 171.745 80.235 171.915 ;
        RECT 80.525 171.405 80.695 171.575 ;
        RECT 80.985 171.405 81.155 171.575 ;
        RECT 84.205 172.085 84.375 172.255 ;
        RECT 85.585 172.085 85.755 172.255 ;
        RECT 86.505 172.085 86.675 172.255 ;
        RECT 87.425 172.085 87.595 172.255 ;
        RECT 90.185 172.085 90.355 172.255 ;
        RECT 18.425 170.895 18.595 171.065 ;
        RECT 18.885 170.895 19.055 171.065 ;
        RECT 19.345 170.895 19.515 171.065 ;
        RECT 19.805 170.895 19.975 171.065 ;
        RECT 20.265 170.895 20.435 171.065 ;
        RECT 20.725 170.895 20.895 171.065 ;
        RECT 21.185 170.895 21.355 171.065 ;
        RECT 21.645 170.895 21.815 171.065 ;
        RECT 22.105 170.895 22.275 171.065 ;
        RECT 22.565 170.895 22.735 171.065 ;
        RECT 23.025 170.895 23.195 171.065 ;
        RECT 23.485 170.895 23.655 171.065 ;
        RECT 23.945 170.895 24.115 171.065 ;
        RECT 24.405 170.895 24.575 171.065 ;
        RECT 24.865 170.895 25.035 171.065 ;
        RECT 25.325 170.895 25.495 171.065 ;
        RECT 25.785 170.895 25.955 171.065 ;
        RECT 26.245 170.895 26.415 171.065 ;
        RECT 26.705 170.895 26.875 171.065 ;
        RECT 27.165 170.895 27.335 171.065 ;
        RECT 27.625 170.895 27.795 171.065 ;
        RECT 28.085 170.895 28.255 171.065 ;
        RECT 28.545 170.895 28.715 171.065 ;
        RECT 29.005 170.895 29.175 171.065 ;
        RECT 29.465 170.895 29.635 171.065 ;
        RECT 29.925 170.895 30.095 171.065 ;
        RECT 30.385 170.895 30.555 171.065 ;
        RECT 30.845 170.895 31.015 171.065 ;
        RECT 31.305 170.895 31.475 171.065 ;
        RECT 31.765 170.895 31.935 171.065 ;
        RECT 32.225 170.895 32.395 171.065 ;
        RECT 32.685 170.895 32.855 171.065 ;
        RECT 33.145 170.895 33.315 171.065 ;
        RECT 33.605 170.895 33.775 171.065 ;
        RECT 34.065 170.895 34.235 171.065 ;
        RECT 34.525 170.895 34.695 171.065 ;
        RECT 34.985 170.895 35.155 171.065 ;
        RECT 35.445 170.895 35.615 171.065 ;
        RECT 35.905 170.895 36.075 171.065 ;
        RECT 36.365 170.895 36.535 171.065 ;
        RECT 36.825 170.895 36.995 171.065 ;
        RECT 37.285 170.895 37.455 171.065 ;
        RECT 37.745 170.895 37.915 171.065 ;
        RECT 38.205 170.895 38.375 171.065 ;
        RECT 38.665 170.895 38.835 171.065 ;
        RECT 39.125 170.895 39.295 171.065 ;
        RECT 39.585 170.895 39.755 171.065 ;
        RECT 40.045 170.895 40.215 171.065 ;
        RECT 40.505 170.895 40.675 171.065 ;
        RECT 40.965 170.895 41.135 171.065 ;
        RECT 41.425 170.895 41.595 171.065 ;
        RECT 41.885 170.895 42.055 171.065 ;
        RECT 42.345 170.895 42.515 171.065 ;
        RECT 42.805 170.895 42.975 171.065 ;
        RECT 43.265 170.895 43.435 171.065 ;
        RECT 43.725 170.895 43.895 171.065 ;
        RECT 44.185 170.895 44.355 171.065 ;
        RECT 44.645 170.895 44.815 171.065 ;
        RECT 45.105 170.895 45.275 171.065 ;
        RECT 45.565 170.895 45.735 171.065 ;
        RECT 46.025 170.895 46.195 171.065 ;
        RECT 46.485 170.895 46.655 171.065 ;
        RECT 46.945 170.895 47.115 171.065 ;
        RECT 47.405 170.895 47.575 171.065 ;
        RECT 47.865 170.895 48.035 171.065 ;
        RECT 48.325 170.895 48.495 171.065 ;
        RECT 48.785 170.895 48.955 171.065 ;
        RECT 49.245 170.895 49.415 171.065 ;
        RECT 49.705 170.895 49.875 171.065 ;
        RECT 50.165 170.895 50.335 171.065 ;
        RECT 50.625 170.895 50.795 171.065 ;
        RECT 51.085 170.895 51.255 171.065 ;
        RECT 51.545 170.895 51.715 171.065 ;
        RECT 52.005 170.895 52.175 171.065 ;
        RECT 52.465 170.895 52.635 171.065 ;
        RECT 52.925 170.895 53.095 171.065 ;
        RECT 53.385 170.895 53.555 171.065 ;
        RECT 53.845 170.895 54.015 171.065 ;
        RECT 54.305 170.895 54.475 171.065 ;
        RECT 54.765 170.895 54.935 171.065 ;
        RECT 55.225 170.895 55.395 171.065 ;
        RECT 55.685 170.895 55.855 171.065 ;
        RECT 56.145 170.895 56.315 171.065 ;
        RECT 56.605 170.895 56.775 171.065 ;
        RECT 57.065 170.895 57.235 171.065 ;
        RECT 57.525 170.895 57.695 171.065 ;
        RECT 57.985 170.895 58.155 171.065 ;
        RECT 58.445 170.895 58.615 171.065 ;
        RECT 58.905 170.895 59.075 171.065 ;
        RECT 59.365 170.895 59.535 171.065 ;
        RECT 59.825 170.895 59.995 171.065 ;
        RECT 60.285 170.895 60.455 171.065 ;
        RECT 60.745 170.895 60.915 171.065 ;
        RECT 61.205 170.895 61.375 171.065 ;
        RECT 61.665 170.895 61.835 171.065 ;
        RECT 62.125 170.895 62.295 171.065 ;
        RECT 62.585 170.895 62.755 171.065 ;
        RECT 63.045 170.895 63.215 171.065 ;
        RECT 63.505 170.895 63.675 171.065 ;
        RECT 63.965 170.895 64.135 171.065 ;
        RECT 64.425 170.895 64.595 171.065 ;
        RECT 64.885 170.895 65.055 171.065 ;
        RECT 65.345 170.895 65.515 171.065 ;
        RECT 65.805 170.895 65.975 171.065 ;
        RECT 66.265 170.895 66.435 171.065 ;
        RECT 66.725 170.895 66.895 171.065 ;
        RECT 67.185 170.895 67.355 171.065 ;
        RECT 67.645 170.895 67.815 171.065 ;
        RECT 68.105 170.895 68.275 171.065 ;
        RECT 68.565 170.895 68.735 171.065 ;
        RECT 69.025 170.895 69.195 171.065 ;
        RECT 69.485 170.895 69.655 171.065 ;
        RECT 69.945 170.895 70.115 171.065 ;
        RECT 70.405 170.895 70.575 171.065 ;
        RECT 70.865 170.895 71.035 171.065 ;
        RECT 71.325 170.895 71.495 171.065 ;
        RECT 71.785 170.895 71.955 171.065 ;
        RECT 72.245 170.895 72.415 171.065 ;
        RECT 72.705 170.895 72.875 171.065 ;
        RECT 73.165 170.895 73.335 171.065 ;
        RECT 73.625 170.895 73.795 171.065 ;
        RECT 74.085 170.895 74.255 171.065 ;
        RECT 74.545 170.895 74.715 171.065 ;
        RECT 75.005 170.895 75.175 171.065 ;
        RECT 75.465 170.895 75.635 171.065 ;
        RECT 75.925 170.895 76.095 171.065 ;
        RECT 76.385 170.895 76.555 171.065 ;
        RECT 76.845 170.895 77.015 171.065 ;
        RECT 77.305 170.895 77.475 171.065 ;
        RECT 77.765 170.895 77.935 171.065 ;
        RECT 78.225 170.895 78.395 171.065 ;
        RECT 78.685 170.895 78.855 171.065 ;
        RECT 79.145 170.895 79.315 171.065 ;
        RECT 79.605 170.895 79.775 171.065 ;
        RECT 80.065 170.895 80.235 171.065 ;
        RECT 80.525 170.895 80.695 171.065 ;
        RECT 80.985 170.895 81.155 171.065 ;
        RECT 81.445 170.895 81.615 171.065 ;
        RECT 81.905 170.895 82.075 171.065 ;
        RECT 82.365 170.895 82.535 171.065 ;
        RECT 82.825 170.895 82.995 171.065 ;
        RECT 83.285 170.895 83.455 171.065 ;
        RECT 83.745 170.895 83.915 171.065 ;
        RECT 84.205 170.895 84.375 171.065 ;
        RECT 84.665 170.895 84.835 171.065 ;
        RECT 85.125 170.895 85.295 171.065 ;
        RECT 85.585 170.895 85.755 171.065 ;
        RECT 86.045 170.895 86.215 171.065 ;
        RECT 86.505 170.895 86.675 171.065 ;
        RECT 86.965 170.895 87.135 171.065 ;
        RECT 87.425 170.895 87.595 171.065 ;
        RECT 87.885 170.895 88.055 171.065 ;
        RECT 88.345 170.895 88.515 171.065 ;
        RECT 88.805 170.895 88.975 171.065 ;
        RECT 89.265 170.895 89.435 171.065 ;
        RECT 89.725 170.895 89.895 171.065 ;
        RECT 90.185 170.895 90.355 171.065 ;
        RECT 90.645 170.895 90.815 171.065 ;
        RECT 91.105 170.895 91.275 171.065 ;
        RECT 91.565 170.895 91.735 171.065 ;
        RECT 92.025 170.895 92.195 171.065 ;
        RECT 33.145 170.385 33.315 170.555 ;
        RECT 35.455 169.365 35.625 169.535 ;
        RECT 35.890 169.025 36.060 169.195 ;
        RECT 37.975 169.365 38.145 169.535 ;
        RECT 37.460 169.025 37.630 169.195 ;
        RECT 38.820 170.045 38.990 170.215 ;
        RECT 39.165 169.365 39.335 169.535 ;
        RECT 40.505 169.705 40.675 169.875 ;
        RECT 40.045 169.365 40.215 169.535 ;
        RECT 41.425 170.045 41.595 170.215 ;
        RECT 42.805 170.045 42.975 170.215 ;
        RECT 41.885 169.705 42.055 169.875 ;
        RECT 42.345 169.705 42.515 169.875 ;
        RECT 43.265 169.705 43.435 169.875 ;
        RECT 39.560 169.025 39.730 169.195 ;
        RECT 40.505 169.025 40.675 169.195 ;
        RECT 44.645 169.365 44.815 169.535 ;
        RECT 45.565 169.705 45.735 169.875 ;
        RECT 46.025 169.705 46.195 169.875 ;
        RECT 46.945 169.705 47.115 169.875 ;
        RECT 47.405 169.705 47.575 169.875 ;
        RECT 47.865 169.705 48.035 169.875 ;
        RECT 49.245 170.045 49.415 170.215 ;
        RECT 48.785 169.705 48.955 169.875 ;
        RECT 48.325 169.365 48.495 169.535 ;
        RECT 50.165 170.385 50.335 170.555 ;
        RECT 50.625 170.045 50.795 170.215 ;
        RECT 51.085 169.705 51.255 169.875 ;
        RECT 52.005 168.685 52.175 168.855 ;
        RECT 61.665 169.705 61.835 169.875 ;
        RECT 63.965 170.385 64.135 170.555 ;
        RECT 62.585 169.705 62.755 169.875 ;
        RECT 60.745 169.365 60.915 169.535 ;
        RECT 63.045 169.705 63.215 169.875 ;
        RECT 73.625 170.045 73.795 170.215 ;
        RECT 72.705 169.705 72.875 169.875 ;
        RECT 74.085 169.705 74.255 169.875 ;
        RECT 74.545 169.705 74.715 169.875 ;
        RECT 76.385 170.045 76.555 170.215 ;
        RECT 75.925 169.705 76.095 169.875 ;
        RECT 76.845 169.705 77.015 169.875 ;
        RECT 75.465 168.685 75.635 168.855 ;
        RECT 82.365 169.365 82.535 169.535 ;
        RECT 82.830 169.025 83.000 169.195 ;
        RECT 83.290 170.045 83.460 170.215 ;
        RECT 83.745 169.705 83.915 169.875 ;
        RECT 84.690 170.045 84.860 170.215 ;
        RECT 86.530 170.045 86.700 170.215 ;
        RECT 85.150 169.025 85.320 169.195 ;
        RECT 86.530 169.025 86.700 169.195 ;
        RECT 90.185 168.685 90.355 168.855 ;
        RECT 18.425 168.175 18.595 168.345 ;
        RECT 18.885 168.175 19.055 168.345 ;
        RECT 19.345 168.175 19.515 168.345 ;
        RECT 19.805 168.175 19.975 168.345 ;
        RECT 20.265 168.175 20.435 168.345 ;
        RECT 20.725 168.175 20.895 168.345 ;
        RECT 21.185 168.175 21.355 168.345 ;
        RECT 21.645 168.175 21.815 168.345 ;
        RECT 22.105 168.175 22.275 168.345 ;
        RECT 22.565 168.175 22.735 168.345 ;
        RECT 23.025 168.175 23.195 168.345 ;
        RECT 23.485 168.175 23.655 168.345 ;
        RECT 23.945 168.175 24.115 168.345 ;
        RECT 24.405 168.175 24.575 168.345 ;
        RECT 24.865 168.175 25.035 168.345 ;
        RECT 25.325 168.175 25.495 168.345 ;
        RECT 25.785 168.175 25.955 168.345 ;
        RECT 26.245 168.175 26.415 168.345 ;
        RECT 26.705 168.175 26.875 168.345 ;
        RECT 27.165 168.175 27.335 168.345 ;
        RECT 27.625 168.175 27.795 168.345 ;
        RECT 28.085 168.175 28.255 168.345 ;
        RECT 28.545 168.175 28.715 168.345 ;
        RECT 29.005 168.175 29.175 168.345 ;
        RECT 29.465 168.175 29.635 168.345 ;
        RECT 29.925 168.175 30.095 168.345 ;
        RECT 30.385 168.175 30.555 168.345 ;
        RECT 30.845 168.175 31.015 168.345 ;
        RECT 31.305 168.175 31.475 168.345 ;
        RECT 31.765 168.175 31.935 168.345 ;
        RECT 32.225 168.175 32.395 168.345 ;
        RECT 32.685 168.175 32.855 168.345 ;
        RECT 33.145 168.175 33.315 168.345 ;
        RECT 33.605 168.175 33.775 168.345 ;
        RECT 34.065 168.175 34.235 168.345 ;
        RECT 34.525 168.175 34.695 168.345 ;
        RECT 34.985 168.175 35.155 168.345 ;
        RECT 35.445 168.175 35.615 168.345 ;
        RECT 35.905 168.175 36.075 168.345 ;
        RECT 36.365 168.175 36.535 168.345 ;
        RECT 36.825 168.175 36.995 168.345 ;
        RECT 37.285 168.175 37.455 168.345 ;
        RECT 37.745 168.175 37.915 168.345 ;
        RECT 38.205 168.175 38.375 168.345 ;
        RECT 38.665 168.175 38.835 168.345 ;
        RECT 39.125 168.175 39.295 168.345 ;
        RECT 39.585 168.175 39.755 168.345 ;
        RECT 40.045 168.175 40.215 168.345 ;
        RECT 40.505 168.175 40.675 168.345 ;
        RECT 40.965 168.175 41.135 168.345 ;
        RECT 41.425 168.175 41.595 168.345 ;
        RECT 41.885 168.175 42.055 168.345 ;
        RECT 42.345 168.175 42.515 168.345 ;
        RECT 42.805 168.175 42.975 168.345 ;
        RECT 43.265 168.175 43.435 168.345 ;
        RECT 43.725 168.175 43.895 168.345 ;
        RECT 44.185 168.175 44.355 168.345 ;
        RECT 44.645 168.175 44.815 168.345 ;
        RECT 45.105 168.175 45.275 168.345 ;
        RECT 45.565 168.175 45.735 168.345 ;
        RECT 46.025 168.175 46.195 168.345 ;
        RECT 46.485 168.175 46.655 168.345 ;
        RECT 46.945 168.175 47.115 168.345 ;
        RECT 47.405 168.175 47.575 168.345 ;
        RECT 47.865 168.175 48.035 168.345 ;
        RECT 48.325 168.175 48.495 168.345 ;
        RECT 48.785 168.175 48.955 168.345 ;
        RECT 49.245 168.175 49.415 168.345 ;
        RECT 49.705 168.175 49.875 168.345 ;
        RECT 50.165 168.175 50.335 168.345 ;
        RECT 50.625 168.175 50.795 168.345 ;
        RECT 51.085 168.175 51.255 168.345 ;
        RECT 51.545 168.175 51.715 168.345 ;
        RECT 52.005 168.175 52.175 168.345 ;
        RECT 52.465 168.175 52.635 168.345 ;
        RECT 52.925 168.175 53.095 168.345 ;
        RECT 53.385 168.175 53.555 168.345 ;
        RECT 53.845 168.175 54.015 168.345 ;
        RECT 54.305 168.175 54.475 168.345 ;
        RECT 54.765 168.175 54.935 168.345 ;
        RECT 55.225 168.175 55.395 168.345 ;
        RECT 55.685 168.175 55.855 168.345 ;
        RECT 56.145 168.175 56.315 168.345 ;
        RECT 56.605 168.175 56.775 168.345 ;
        RECT 57.065 168.175 57.235 168.345 ;
        RECT 57.525 168.175 57.695 168.345 ;
        RECT 57.985 168.175 58.155 168.345 ;
        RECT 58.445 168.175 58.615 168.345 ;
        RECT 58.905 168.175 59.075 168.345 ;
        RECT 59.365 168.175 59.535 168.345 ;
        RECT 59.825 168.175 59.995 168.345 ;
        RECT 60.285 168.175 60.455 168.345 ;
        RECT 60.745 168.175 60.915 168.345 ;
        RECT 61.205 168.175 61.375 168.345 ;
        RECT 61.665 168.175 61.835 168.345 ;
        RECT 62.125 168.175 62.295 168.345 ;
        RECT 62.585 168.175 62.755 168.345 ;
        RECT 63.045 168.175 63.215 168.345 ;
        RECT 63.505 168.175 63.675 168.345 ;
        RECT 63.965 168.175 64.135 168.345 ;
        RECT 64.425 168.175 64.595 168.345 ;
        RECT 64.885 168.175 65.055 168.345 ;
        RECT 65.345 168.175 65.515 168.345 ;
        RECT 65.805 168.175 65.975 168.345 ;
        RECT 66.265 168.175 66.435 168.345 ;
        RECT 66.725 168.175 66.895 168.345 ;
        RECT 67.185 168.175 67.355 168.345 ;
        RECT 67.645 168.175 67.815 168.345 ;
        RECT 68.105 168.175 68.275 168.345 ;
        RECT 68.565 168.175 68.735 168.345 ;
        RECT 69.025 168.175 69.195 168.345 ;
        RECT 69.485 168.175 69.655 168.345 ;
        RECT 69.945 168.175 70.115 168.345 ;
        RECT 70.405 168.175 70.575 168.345 ;
        RECT 70.865 168.175 71.035 168.345 ;
        RECT 71.325 168.175 71.495 168.345 ;
        RECT 71.785 168.175 71.955 168.345 ;
        RECT 72.245 168.175 72.415 168.345 ;
        RECT 72.705 168.175 72.875 168.345 ;
        RECT 73.165 168.175 73.335 168.345 ;
        RECT 73.625 168.175 73.795 168.345 ;
        RECT 74.085 168.175 74.255 168.345 ;
        RECT 74.545 168.175 74.715 168.345 ;
        RECT 75.005 168.175 75.175 168.345 ;
        RECT 75.465 168.175 75.635 168.345 ;
        RECT 75.925 168.175 76.095 168.345 ;
        RECT 76.385 168.175 76.555 168.345 ;
        RECT 76.845 168.175 77.015 168.345 ;
        RECT 77.305 168.175 77.475 168.345 ;
        RECT 77.765 168.175 77.935 168.345 ;
        RECT 78.225 168.175 78.395 168.345 ;
        RECT 78.685 168.175 78.855 168.345 ;
        RECT 79.145 168.175 79.315 168.345 ;
        RECT 79.605 168.175 79.775 168.345 ;
        RECT 80.065 168.175 80.235 168.345 ;
        RECT 80.525 168.175 80.695 168.345 ;
        RECT 80.985 168.175 81.155 168.345 ;
        RECT 81.445 168.175 81.615 168.345 ;
        RECT 81.905 168.175 82.075 168.345 ;
        RECT 82.365 168.175 82.535 168.345 ;
        RECT 82.825 168.175 82.995 168.345 ;
        RECT 83.285 168.175 83.455 168.345 ;
        RECT 83.745 168.175 83.915 168.345 ;
        RECT 84.205 168.175 84.375 168.345 ;
        RECT 84.665 168.175 84.835 168.345 ;
        RECT 85.125 168.175 85.295 168.345 ;
        RECT 85.585 168.175 85.755 168.345 ;
        RECT 86.045 168.175 86.215 168.345 ;
        RECT 86.505 168.175 86.675 168.345 ;
        RECT 86.965 168.175 87.135 168.345 ;
        RECT 87.425 168.175 87.595 168.345 ;
        RECT 87.885 168.175 88.055 168.345 ;
        RECT 88.345 168.175 88.515 168.345 ;
        RECT 88.805 168.175 88.975 168.345 ;
        RECT 89.265 168.175 89.435 168.345 ;
        RECT 89.725 168.175 89.895 168.345 ;
        RECT 90.185 168.175 90.355 168.345 ;
        RECT 90.645 168.175 90.815 168.345 ;
        RECT 91.105 168.175 91.275 168.345 ;
        RECT 91.565 168.175 91.735 168.345 ;
        RECT 92.025 168.175 92.195 168.345 ;
        RECT 55.225 167.665 55.395 167.835 ;
        RECT 53.845 166.645 54.015 166.815 ;
        RECT 54.305 166.645 54.475 166.815 ;
        RECT 60.745 166.985 60.915 167.155 ;
        RECT 58.445 166.645 58.615 166.815 ;
        RECT 59.955 166.645 60.125 166.815 ;
        RECT 57.525 165.965 57.695 166.135 ;
        RECT 61.665 166.305 61.835 166.475 ;
        RECT 63.505 166.305 63.675 166.475 ;
        RECT 72.245 165.965 72.415 166.135 ;
        RECT 77.765 167.325 77.935 167.495 ;
        RECT 75.465 166.645 75.635 166.815 ;
        RECT 76.385 166.645 76.555 166.815 ;
        RECT 76.845 166.645 77.015 166.815 ;
        RECT 78.255 166.645 78.425 166.815 ;
        RECT 77.765 166.305 77.935 166.475 ;
        RECT 79.145 166.645 79.315 166.815 ;
        RECT 78.685 166.305 78.855 166.475 ;
        RECT 18.425 165.455 18.595 165.625 ;
        RECT 18.885 165.455 19.055 165.625 ;
        RECT 19.345 165.455 19.515 165.625 ;
        RECT 19.805 165.455 19.975 165.625 ;
        RECT 20.265 165.455 20.435 165.625 ;
        RECT 20.725 165.455 20.895 165.625 ;
        RECT 21.185 165.455 21.355 165.625 ;
        RECT 21.645 165.455 21.815 165.625 ;
        RECT 22.105 165.455 22.275 165.625 ;
        RECT 22.565 165.455 22.735 165.625 ;
        RECT 23.025 165.455 23.195 165.625 ;
        RECT 23.485 165.455 23.655 165.625 ;
        RECT 23.945 165.455 24.115 165.625 ;
        RECT 24.405 165.455 24.575 165.625 ;
        RECT 24.865 165.455 25.035 165.625 ;
        RECT 25.325 165.455 25.495 165.625 ;
        RECT 25.785 165.455 25.955 165.625 ;
        RECT 26.245 165.455 26.415 165.625 ;
        RECT 26.705 165.455 26.875 165.625 ;
        RECT 27.165 165.455 27.335 165.625 ;
        RECT 27.625 165.455 27.795 165.625 ;
        RECT 28.085 165.455 28.255 165.625 ;
        RECT 28.545 165.455 28.715 165.625 ;
        RECT 29.005 165.455 29.175 165.625 ;
        RECT 29.465 165.455 29.635 165.625 ;
        RECT 29.925 165.455 30.095 165.625 ;
        RECT 30.385 165.455 30.555 165.625 ;
        RECT 30.845 165.455 31.015 165.625 ;
        RECT 31.305 165.455 31.475 165.625 ;
        RECT 31.765 165.455 31.935 165.625 ;
        RECT 32.225 165.455 32.395 165.625 ;
        RECT 32.685 165.455 32.855 165.625 ;
        RECT 33.145 165.455 33.315 165.625 ;
        RECT 33.605 165.455 33.775 165.625 ;
        RECT 34.065 165.455 34.235 165.625 ;
        RECT 34.525 165.455 34.695 165.625 ;
        RECT 34.985 165.455 35.155 165.625 ;
        RECT 35.445 165.455 35.615 165.625 ;
        RECT 35.905 165.455 36.075 165.625 ;
        RECT 36.365 165.455 36.535 165.625 ;
        RECT 36.825 165.455 36.995 165.625 ;
        RECT 37.285 165.455 37.455 165.625 ;
        RECT 37.745 165.455 37.915 165.625 ;
        RECT 38.205 165.455 38.375 165.625 ;
        RECT 38.665 165.455 38.835 165.625 ;
        RECT 39.125 165.455 39.295 165.625 ;
        RECT 39.585 165.455 39.755 165.625 ;
        RECT 40.045 165.455 40.215 165.625 ;
        RECT 40.505 165.455 40.675 165.625 ;
        RECT 40.965 165.455 41.135 165.625 ;
        RECT 41.425 165.455 41.595 165.625 ;
        RECT 41.885 165.455 42.055 165.625 ;
        RECT 42.345 165.455 42.515 165.625 ;
        RECT 42.805 165.455 42.975 165.625 ;
        RECT 43.265 165.455 43.435 165.625 ;
        RECT 43.725 165.455 43.895 165.625 ;
        RECT 44.185 165.455 44.355 165.625 ;
        RECT 44.645 165.455 44.815 165.625 ;
        RECT 45.105 165.455 45.275 165.625 ;
        RECT 45.565 165.455 45.735 165.625 ;
        RECT 46.025 165.455 46.195 165.625 ;
        RECT 46.485 165.455 46.655 165.625 ;
        RECT 46.945 165.455 47.115 165.625 ;
        RECT 47.405 165.455 47.575 165.625 ;
        RECT 47.865 165.455 48.035 165.625 ;
        RECT 48.325 165.455 48.495 165.625 ;
        RECT 48.785 165.455 48.955 165.625 ;
        RECT 49.245 165.455 49.415 165.625 ;
        RECT 49.705 165.455 49.875 165.625 ;
        RECT 50.165 165.455 50.335 165.625 ;
        RECT 50.625 165.455 50.795 165.625 ;
        RECT 51.085 165.455 51.255 165.625 ;
        RECT 51.545 165.455 51.715 165.625 ;
        RECT 52.005 165.455 52.175 165.625 ;
        RECT 52.465 165.455 52.635 165.625 ;
        RECT 52.925 165.455 53.095 165.625 ;
        RECT 53.385 165.455 53.555 165.625 ;
        RECT 53.845 165.455 54.015 165.625 ;
        RECT 54.305 165.455 54.475 165.625 ;
        RECT 54.765 165.455 54.935 165.625 ;
        RECT 55.225 165.455 55.395 165.625 ;
        RECT 55.685 165.455 55.855 165.625 ;
        RECT 56.145 165.455 56.315 165.625 ;
        RECT 56.605 165.455 56.775 165.625 ;
        RECT 57.065 165.455 57.235 165.625 ;
        RECT 57.525 165.455 57.695 165.625 ;
        RECT 57.985 165.455 58.155 165.625 ;
        RECT 58.445 165.455 58.615 165.625 ;
        RECT 58.905 165.455 59.075 165.625 ;
        RECT 59.365 165.455 59.535 165.625 ;
        RECT 59.825 165.455 59.995 165.625 ;
        RECT 60.285 165.455 60.455 165.625 ;
        RECT 60.745 165.455 60.915 165.625 ;
        RECT 61.205 165.455 61.375 165.625 ;
        RECT 61.665 165.455 61.835 165.625 ;
        RECT 62.125 165.455 62.295 165.625 ;
        RECT 62.585 165.455 62.755 165.625 ;
        RECT 63.045 165.455 63.215 165.625 ;
        RECT 63.505 165.455 63.675 165.625 ;
        RECT 63.965 165.455 64.135 165.625 ;
        RECT 64.425 165.455 64.595 165.625 ;
        RECT 64.885 165.455 65.055 165.625 ;
        RECT 65.345 165.455 65.515 165.625 ;
        RECT 65.805 165.455 65.975 165.625 ;
        RECT 66.265 165.455 66.435 165.625 ;
        RECT 66.725 165.455 66.895 165.625 ;
        RECT 67.185 165.455 67.355 165.625 ;
        RECT 67.645 165.455 67.815 165.625 ;
        RECT 68.105 165.455 68.275 165.625 ;
        RECT 68.565 165.455 68.735 165.625 ;
        RECT 69.025 165.455 69.195 165.625 ;
        RECT 69.485 165.455 69.655 165.625 ;
        RECT 69.945 165.455 70.115 165.625 ;
        RECT 70.405 165.455 70.575 165.625 ;
        RECT 70.865 165.455 71.035 165.625 ;
        RECT 71.325 165.455 71.495 165.625 ;
        RECT 71.785 165.455 71.955 165.625 ;
        RECT 72.245 165.455 72.415 165.625 ;
        RECT 72.705 165.455 72.875 165.625 ;
        RECT 73.165 165.455 73.335 165.625 ;
        RECT 73.625 165.455 73.795 165.625 ;
        RECT 74.085 165.455 74.255 165.625 ;
        RECT 74.545 165.455 74.715 165.625 ;
        RECT 75.005 165.455 75.175 165.625 ;
        RECT 75.465 165.455 75.635 165.625 ;
        RECT 75.925 165.455 76.095 165.625 ;
        RECT 76.385 165.455 76.555 165.625 ;
        RECT 76.845 165.455 77.015 165.625 ;
        RECT 77.305 165.455 77.475 165.625 ;
        RECT 77.765 165.455 77.935 165.625 ;
        RECT 78.225 165.455 78.395 165.625 ;
        RECT 78.685 165.455 78.855 165.625 ;
        RECT 79.145 165.455 79.315 165.625 ;
        RECT 79.605 165.455 79.775 165.625 ;
        RECT 80.065 165.455 80.235 165.625 ;
        RECT 80.525 165.455 80.695 165.625 ;
        RECT 80.985 165.455 81.155 165.625 ;
        RECT 81.445 165.455 81.615 165.625 ;
        RECT 81.905 165.455 82.075 165.625 ;
        RECT 82.365 165.455 82.535 165.625 ;
        RECT 82.825 165.455 82.995 165.625 ;
        RECT 83.285 165.455 83.455 165.625 ;
        RECT 83.745 165.455 83.915 165.625 ;
        RECT 84.205 165.455 84.375 165.625 ;
        RECT 84.665 165.455 84.835 165.625 ;
        RECT 85.125 165.455 85.295 165.625 ;
        RECT 85.585 165.455 85.755 165.625 ;
        RECT 86.045 165.455 86.215 165.625 ;
        RECT 86.505 165.455 86.675 165.625 ;
        RECT 86.965 165.455 87.135 165.625 ;
        RECT 87.425 165.455 87.595 165.625 ;
        RECT 87.885 165.455 88.055 165.625 ;
        RECT 88.345 165.455 88.515 165.625 ;
        RECT 88.805 165.455 88.975 165.625 ;
        RECT 89.265 165.455 89.435 165.625 ;
        RECT 89.725 165.455 89.895 165.625 ;
        RECT 90.185 165.455 90.355 165.625 ;
        RECT 90.645 165.455 90.815 165.625 ;
        RECT 91.105 165.455 91.275 165.625 ;
        RECT 91.565 165.455 91.735 165.625 ;
        RECT 92.025 165.455 92.195 165.625 ;
        RECT 48.325 164.945 48.495 165.115 ;
        RECT 49.165 164.945 49.335 165.115 ;
        RECT 38.665 164.265 38.835 164.435 ;
        RECT 39.585 164.265 39.755 164.435 ;
        RECT 38.665 163.245 38.835 163.415 ;
        RECT 45.565 164.265 45.735 164.435 ;
        RECT 44.645 163.925 44.815 164.095 ;
        RECT 46.485 164.265 46.655 164.435 ;
        RECT 46.945 164.265 47.115 164.435 ;
        RECT 46.025 163.585 46.195 163.755 ;
        RECT 47.865 164.265 48.035 164.435 ;
        RECT 50.165 164.605 50.335 164.775 ;
        RECT 56.145 164.945 56.315 165.115 ;
        RECT 51.545 164.265 51.715 164.435 ;
        RECT 52.925 164.265 53.095 164.435 ;
        RECT 52.465 163.925 52.635 164.095 ;
        RECT 53.845 164.265 54.015 164.435 ;
        RECT 54.305 164.265 54.475 164.435 ;
        RECT 50.625 163.585 50.795 163.755 ;
        RECT 49.245 163.245 49.415 163.415 ;
        RECT 55.225 164.265 55.395 164.435 ;
        RECT 57.525 164.265 57.695 164.435 ;
        RECT 56.605 163.925 56.775 164.095 ;
        RECT 58.905 164.945 59.075 165.115 ;
        RECT 58.445 163.245 58.615 163.415 ;
        RECT 61.215 163.925 61.385 164.095 ;
        RECT 61.650 163.585 61.820 163.755 ;
        RECT 63.735 163.925 63.905 164.095 ;
        RECT 63.220 163.585 63.390 163.755 ;
        RECT 64.470 164.265 64.640 164.435 ;
        RECT 64.925 163.925 65.095 164.095 ;
        RECT 69.485 164.945 69.655 165.115 ;
        RECT 65.805 164.265 65.975 164.435 ;
        RECT 67.185 164.265 67.355 164.435 ;
        RECT 68.565 164.265 68.735 164.435 ;
        RECT 67.645 163.925 67.815 164.095 ;
        RECT 65.320 163.585 65.490 163.755 ;
        RECT 70.405 164.265 70.575 164.435 ;
        RECT 70.890 163.585 71.060 163.755 ;
        RECT 71.285 163.925 71.455 164.095 ;
        RECT 71.630 164.605 71.800 164.775 ;
        RECT 72.475 163.925 72.645 164.095 ;
        RECT 72.990 163.585 73.160 163.755 ;
        RECT 74.560 163.585 74.730 163.755 ;
        RECT 74.995 163.925 75.165 164.095 ;
        RECT 77.305 164.945 77.475 165.115 ;
        RECT 77.765 163.925 77.935 164.095 ;
        RECT 78.685 164.265 78.855 164.435 ;
        RECT 79.145 164.265 79.315 164.435 ;
        RECT 80.985 164.265 81.155 164.435 ;
        RECT 78.225 163.245 78.395 163.415 ;
        RECT 82.365 164.265 82.535 164.435 ;
        RECT 81.905 163.925 82.075 164.095 ;
        RECT 81.445 163.245 81.615 163.415 ;
        RECT 82.830 163.585 83.000 163.755 ;
        RECT 83.290 164.605 83.460 164.775 ;
        RECT 83.745 163.925 83.915 164.095 ;
        RECT 84.690 164.605 84.860 164.775 ;
        RECT 86.530 164.605 86.700 164.775 ;
        RECT 85.150 163.585 85.320 163.755 ;
        RECT 86.530 163.585 86.700 163.755 ;
        RECT 90.185 163.245 90.355 163.415 ;
        RECT 18.425 162.735 18.595 162.905 ;
        RECT 18.885 162.735 19.055 162.905 ;
        RECT 19.345 162.735 19.515 162.905 ;
        RECT 19.805 162.735 19.975 162.905 ;
        RECT 20.265 162.735 20.435 162.905 ;
        RECT 20.725 162.735 20.895 162.905 ;
        RECT 21.185 162.735 21.355 162.905 ;
        RECT 21.645 162.735 21.815 162.905 ;
        RECT 22.105 162.735 22.275 162.905 ;
        RECT 22.565 162.735 22.735 162.905 ;
        RECT 23.025 162.735 23.195 162.905 ;
        RECT 23.485 162.735 23.655 162.905 ;
        RECT 23.945 162.735 24.115 162.905 ;
        RECT 24.405 162.735 24.575 162.905 ;
        RECT 24.865 162.735 25.035 162.905 ;
        RECT 25.325 162.735 25.495 162.905 ;
        RECT 25.785 162.735 25.955 162.905 ;
        RECT 26.245 162.735 26.415 162.905 ;
        RECT 26.705 162.735 26.875 162.905 ;
        RECT 27.165 162.735 27.335 162.905 ;
        RECT 27.625 162.735 27.795 162.905 ;
        RECT 28.085 162.735 28.255 162.905 ;
        RECT 28.545 162.735 28.715 162.905 ;
        RECT 29.005 162.735 29.175 162.905 ;
        RECT 29.465 162.735 29.635 162.905 ;
        RECT 29.925 162.735 30.095 162.905 ;
        RECT 30.385 162.735 30.555 162.905 ;
        RECT 30.845 162.735 31.015 162.905 ;
        RECT 31.305 162.735 31.475 162.905 ;
        RECT 31.765 162.735 31.935 162.905 ;
        RECT 32.225 162.735 32.395 162.905 ;
        RECT 32.685 162.735 32.855 162.905 ;
        RECT 33.145 162.735 33.315 162.905 ;
        RECT 33.605 162.735 33.775 162.905 ;
        RECT 34.065 162.735 34.235 162.905 ;
        RECT 34.525 162.735 34.695 162.905 ;
        RECT 34.985 162.735 35.155 162.905 ;
        RECT 35.445 162.735 35.615 162.905 ;
        RECT 35.905 162.735 36.075 162.905 ;
        RECT 36.365 162.735 36.535 162.905 ;
        RECT 36.825 162.735 36.995 162.905 ;
        RECT 37.285 162.735 37.455 162.905 ;
        RECT 37.745 162.735 37.915 162.905 ;
        RECT 38.205 162.735 38.375 162.905 ;
        RECT 38.665 162.735 38.835 162.905 ;
        RECT 39.125 162.735 39.295 162.905 ;
        RECT 39.585 162.735 39.755 162.905 ;
        RECT 40.045 162.735 40.215 162.905 ;
        RECT 40.505 162.735 40.675 162.905 ;
        RECT 40.965 162.735 41.135 162.905 ;
        RECT 41.425 162.735 41.595 162.905 ;
        RECT 41.885 162.735 42.055 162.905 ;
        RECT 42.345 162.735 42.515 162.905 ;
        RECT 42.805 162.735 42.975 162.905 ;
        RECT 43.265 162.735 43.435 162.905 ;
        RECT 43.725 162.735 43.895 162.905 ;
        RECT 44.185 162.735 44.355 162.905 ;
        RECT 44.645 162.735 44.815 162.905 ;
        RECT 45.105 162.735 45.275 162.905 ;
        RECT 45.565 162.735 45.735 162.905 ;
        RECT 46.025 162.735 46.195 162.905 ;
        RECT 46.485 162.735 46.655 162.905 ;
        RECT 46.945 162.735 47.115 162.905 ;
        RECT 47.405 162.735 47.575 162.905 ;
        RECT 47.865 162.735 48.035 162.905 ;
        RECT 48.325 162.735 48.495 162.905 ;
        RECT 48.785 162.735 48.955 162.905 ;
        RECT 49.245 162.735 49.415 162.905 ;
        RECT 49.705 162.735 49.875 162.905 ;
        RECT 50.165 162.735 50.335 162.905 ;
        RECT 50.625 162.735 50.795 162.905 ;
        RECT 51.085 162.735 51.255 162.905 ;
        RECT 51.545 162.735 51.715 162.905 ;
        RECT 52.005 162.735 52.175 162.905 ;
        RECT 52.465 162.735 52.635 162.905 ;
        RECT 52.925 162.735 53.095 162.905 ;
        RECT 53.385 162.735 53.555 162.905 ;
        RECT 53.845 162.735 54.015 162.905 ;
        RECT 54.305 162.735 54.475 162.905 ;
        RECT 54.765 162.735 54.935 162.905 ;
        RECT 55.225 162.735 55.395 162.905 ;
        RECT 55.685 162.735 55.855 162.905 ;
        RECT 56.145 162.735 56.315 162.905 ;
        RECT 56.605 162.735 56.775 162.905 ;
        RECT 57.065 162.735 57.235 162.905 ;
        RECT 57.525 162.735 57.695 162.905 ;
        RECT 57.985 162.735 58.155 162.905 ;
        RECT 58.445 162.735 58.615 162.905 ;
        RECT 58.905 162.735 59.075 162.905 ;
        RECT 59.365 162.735 59.535 162.905 ;
        RECT 59.825 162.735 59.995 162.905 ;
        RECT 60.285 162.735 60.455 162.905 ;
        RECT 60.745 162.735 60.915 162.905 ;
        RECT 61.205 162.735 61.375 162.905 ;
        RECT 61.665 162.735 61.835 162.905 ;
        RECT 62.125 162.735 62.295 162.905 ;
        RECT 62.585 162.735 62.755 162.905 ;
        RECT 63.045 162.735 63.215 162.905 ;
        RECT 63.505 162.735 63.675 162.905 ;
        RECT 63.965 162.735 64.135 162.905 ;
        RECT 64.425 162.735 64.595 162.905 ;
        RECT 64.885 162.735 65.055 162.905 ;
        RECT 65.345 162.735 65.515 162.905 ;
        RECT 65.805 162.735 65.975 162.905 ;
        RECT 66.265 162.735 66.435 162.905 ;
        RECT 66.725 162.735 66.895 162.905 ;
        RECT 67.185 162.735 67.355 162.905 ;
        RECT 67.645 162.735 67.815 162.905 ;
        RECT 68.105 162.735 68.275 162.905 ;
        RECT 68.565 162.735 68.735 162.905 ;
        RECT 69.025 162.735 69.195 162.905 ;
        RECT 69.485 162.735 69.655 162.905 ;
        RECT 69.945 162.735 70.115 162.905 ;
        RECT 70.405 162.735 70.575 162.905 ;
        RECT 70.865 162.735 71.035 162.905 ;
        RECT 71.325 162.735 71.495 162.905 ;
        RECT 71.785 162.735 71.955 162.905 ;
        RECT 72.245 162.735 72.415 162.905 ;
        RECT 72.705 162.735 72.875 162.905 ;
        RECT 73.165 162.735 73.335 162.905 ;
        RECT 73.625 162.735 73.795 162.905 ;
        RECT 74.085 162.735 74.255 162.905 ;
        RECT 74.545 162.735 74.715 162.905 ;
        RECT 75.005 162.735 75.175 162.905 ;
        RECT 75.465 162.735 75.635 162.905 ;
        RECT 75.925 162.735 76.095 162.905 ;
        RECT 76.385 162.735 76.555 162.905 ;
        RECT 76.845 162.735 77.015 162.905 ;
        RECT 77.305 162.735 77.475 162.905 ;
        RECT 77.765 162.735 77.935 162.905 ;
        RECT 78.225 162.735 78.395 162.905 ;
        RECT 78.685 162.735 78.855 162.905 ;
        RECT 79.145 162.735 79.315 162.905 ;
        RECT 79.605 162.735 79.775 162.905 ;
        RECT 80.065 162.735 80.235 162.905 ;
        RECT 80.525 162.735 80.695 162.905 ;
        RECT 80.985 162.735 81.155 162.905 ;
        RECT 81.445 162.735 81.615 162.905 ;
        RECT 81.905 162.735 82.075 162.905 ;
        RECT 82.365 162.735 82.535 162.905 ;
        RECT 82.825 162.735 82.995 162.905 ;
        RECT 83.285 162.735 83.455 162.905 ;
        RECT 83.745 162.735 83.915 162.905 ;
        RECT 84.205 162.735 84.375 162.905 ;
        RECT 84.665 162.735 84.835 162.905 ;
        RECT 85.125 162.735 85.295 162.905 ;
        RECT 85.585 162.735 85.755 162.905 ;
        RECT 86.045 162.735 86.215 162.905 ;
        RECT 86.505 162.735 86.675 162.905 ;
        RECT 86.965 162.735 87.135 162.905 ;
        RECT 87.425 162.735 87.595 162.905 ;
        RECT 87.885 162.735 88.055 162.905 ;
        RECT 88.345 162.735 88.515 162.905 ;
        RECT 88.805 162.735 88.975 162.905 ;
        RECT 89.265 162.735 89.435 162.905 ;
        RECT 89.725 162.735 89.895 162.905 ;
        RECT 90.185 162.735 90.355 162.905 ;
        RECT 90.645 162.735 90.815 162.905 ;
        RECT 91.105 162.735 91.275 162.905 ;
        RECT 91.565 162.735 91.735 162.905 ;
        RECT 92.025 162.735 92.195 162.905 ;
        RECT 36.850 161.885 37.020 162.055 ;
        RECT 36.365 161.205 36.535 161.375 ;
        RECT 37.245 161.545 37.415 161.715 ;
        RECT 37.700 160.865 37.870 161.035 ;
        RECT 38.950 161.885 39.120 162.055 ;
        RECT 38.435 161.545 38.605 161.715 ;
        RECT 40.520 161.885 40.690 162.055 ;
        RECT 40.955 161.545 41.125 161.715 ;
        RECT 43.265 161.885 43.435 162.055 ;
        RECT 47.405 162.225 47.575 162.395 ;
        RECT 46.945 161.205 47.115 161.375 ;
        RECT 52.465 162.225 52.635 162.395 ;
        RECT 51.545 161.885 51.715 162.055 ;
        RECT 52.235 161.035 52.405 161.205 ;
        RECT 53.845 161.205 54.015 161.375 ;
        RECT 53.385 160.865 53.555 161.035 ;
        RECT 54.765 161.205 54.935 161.375 ;
        RECT 54.305 160.525 54.475 160.695 ;
        RECT 59.365 161.545 59.535 161.715 ;
        RECT 61.205 162.225 61.375 162.395 ;
        RECT 57.985 160.865 58.155 161.035 ;
        RECT 60.285 161.205 60.455 161.375 ;
        RECT 68.565 162.225 68.735 162.395 ;
        RECT 68.565 160.865 68.735 161.035 ;
        RECT 69.945 161.205 70.115 161.375 ;
        RECT 69.485 160.525 69.655 160.695 ;
        RECT 76.845 162.225 77.015 162.395 ;
        RECT 79.145 161.885 79.315 162.055 ;
        RECT 76.335 161.205 76.505 161.375 ;
        RECT 77.305 161.205 77.475 161.375 ;
        RECT 77.765 161.205 77.935 161.375 ;
        RECT 78.225 161.205 78.395 161.375 ;
        RECT 79.145 161.205 79.315 161.375 ;
        RECT 83.285 162.225 83.455 162.395 ;
        RECT 83.285 161.205 83.455 161.375 ;
        RECT 84.665 161.205 84.835 161.375 ;
        RECT 84.205 160.525 84.375 160.695 ;
        RECT 18.425 160.015 18.595 160.185 ;
        RECT 18.885 160.015 19.055 160.185 ;
        RECT 19.345 160.015 19.515 160.185 ;
        RECT 19.805 160.015 19.975 160.185 ;
        RECT 20.265 160.015 20.435 160.185 ;
        RECT 20.725 160.015 20.895 160.185 ;
        RECT 21.185 160.015 21.355 160.185 ;
        RECT 21.645 160.015 21.815 160.185 ;
        RECT 22.105 160.015 22.275 160.185 ;
        RECT 22.565 160.015 22.735 160.185 ;
        RECT 23.025 160.015 23.195 160.185 ;
        RECT 23.485 160.015 23.655 160.185 ;
        RECT 23.945 160.015 24.115 160.185 ;
        RECT 24.405 160.015 24.575 160.185 ;
        RECT 24.865 160.015 25.035 160.185 ;
        RECT 25.325 160.015 25.495 160.185 ;
        RECT 25.785 160.015 25.955 160.185 ;
        RECT 26.245 160.015 26.415 160.185 ;
        RECT 26.705 160.015 26.875 160.185 ;
        RECT 27.165 160.015 27.335 160.185 ;
        RECT 27.625 160.015 27.795 160.185 ;
        RECT 28.085 160.015 28.255 160.185 ;
        RECT 28.545 160.015 28.715 160.185 ;
        RECT 29.005 160.015 29.175 160.185 ;
        RECT 29.465 160.015 29.635 160.185 ;
        RECT 29.925 160.015 30.095 160.185 ;
        RECT 30.385 160.015 30.555 160.185 ;
        RECT 30.845 160.015 31.015 160.185 ;
        RECT 31.305 160.015 31.475 160.185 ;
        RECT 31.765 160.015 31.935 160.185 ;
        RECT 32.225 160.015 32.395 160.185 ;
        RECT 32.685 160.015 32.855 160.185 ;
        RECT 33.145 160.015 33.315 160.185 ;
        RECT 33.605 160.015 33.775 160.185 ;
        RECT 34.065 160.015 34.235 160.185 ;
        RECT 34.525 160.015 34.695 160.185 ;
        RECT 34.985 160.015 35.155 160.185 ;
        RECT 35.445 160.015 35.615 160.185 ;
        RECT 35.905 160.015 36.075 160.185 ;
        RECT 36.365 160.015 36.535 160.185 ;
        RECT 36.825 160.015 36.995 160.185 ;
        RECT 37.285 160.015 37.455 160.185 ;
        RECT 37.745 160.015 37.915 160.185 ;
        RECT 38.205 160.015 38.375 160.185 ;
        RECT 38.665 160.015 38.835 160.185 ;
        RECT 39.125 160.015 39.295 160.185 ;
        RECT 39.585 160.015 39.755 160.185 ;
        RECT 40.045 160.015 40.215 160.185 ;
        RECT 40.505 160.015 40.675 160.185 ;
        RECT 40.965 160.015 41.135 160.185 ;
        RECT 41.425 160.015 41.595 160.185 ;
        RECT 41.885 160.015 42.055 160.185 ;
        RECT 42.345 160.015 42.515 160.185 ;
        RECT 42.805 160.015 42.975 160.185 ;
        RECT 43.265 160.015 43.435 160.185 ;
        RECT 43.725 160.015 43.895 160.185 ;
        RECT 44.185 160.015 44.355 160.185 ;
        RECT 44.645 160.015 44.815 160.185 ;
        RECT 45.105 160.015 45.275 160.185 ;
        RECT 45.565 160.015 45.735 160.185 ;
        RECT 46.025 160.015 46.195 160.185 ;
        RECT 46.485 160.015 46.655 160.185 ;
        RECT 46.945 160.015 47.115 160.185 ;
        RECT 47.405 160.015 47.575 160.185 ;
        RECT 47.865 160.015 48.035 160.185 ;
        RECT 48.325 160.015 48.495 160.185 ;
        RECT 48.785 160.015 48.955 160.185 ;
        RECT 49.245 160.015 49.415 160.185 ;
        RECT 49.705 160.015 49.875 160.185 ;
        RECT 50.165 160.015 50.335 160.185 ;
        RECT 50.625 160.015 50.795 160.185 ;
        RECT 51.085 160.015 51.255 160.185 ;
        RECT 51.545 160.015 51.715 160.185 ;
        RECT 52.005 160.015 52.175 160.185 ;
        RECT 52.465 160.015 52.635 160.185 ;
        RECT 52.925 160.015 53.095 160.185 ;
        RECT 53.385 160.015 53.555 160.185 ;
        RECT 53.845 160.015 54.015 160.185 ;
        RECT 54.305 160.015 54.475 160.185 ;
        RECT 54.765 160.015 54.935 160.185 ;
        RECT 55.225 160.015 55.395 160.185 ;
        RECT 55.685 160.015 55.855 160.185 ;
        RECT 56.145 160.015 56.315 160.185 ;
        RECT 56.605 160.015 56.775 160.185 ;
        RECT 57.065 160.015 57.235 160.185 ;
        RECT 57.525 160.015 57.695 160.185 ;
        RECT 57.985 160.015 58.155 160.185 ;
        RECT 58.445 160.015 58.615 160.185 ;
        RECT 58.905 160.015 59.075 160.185 ;
        RECT 59.365 160.015 59.535 160.185 ;
        RECT 59.825 160.015 59.995 160.185 ;
        RECT 60.285 160.015 60.455 160.185 ;
        RECT 60.745 160.015 60.915 160.185 ;
        RECT 61.205 160.015 61.375 160.185 ;
        RECT 61.665 160.015 61.835 160.185 ;
        RECT 62.125 160.015 62.295 160.185 ;
        RECT 62.585 160.015 62.755 160.185 ;
        RECT 63.045 160.015 63.215 160.185 ;
        RECT 63.505 160.015 63.675 160.185 ;
        RECT 63.965 160.015 64.135 160.185 ;
        RECT 64.425 160.015 64.595 160.185 ;
        RECT 64.885 160.015 65.055 160.185 ;
        RECT 65.345 160.015 65.515 160.185 ;
        RECT 65.805 160.015 65.975 160.185 ;
        RECT 66.265 160.015 66.435 160.185 ;
        RECT 66.725 160.015 66.895 160.185 ;
        RECT 67.185 160.015 67.355 160.185 ;
        RECT 67.645 160.015 67.815 160.185 ;
        RECT 68.105 160.015 68.275 160.185 ;
        RECT 68.565 160.015 68.735 160.185 ;
        RECT 69.025 160.015 69.195 160.185 ;
        RECT 69.485 160.015 69.655 160.185 ;
        RECT 69.945 160.015 70.115 160.185 ;
        RECT 70.405 160.015 70.575 160.185 ;
        RECT 70.865 160.015 71.035 160.185 ;
        RECT 71.325 160.015 71.495 160.185 ;
        RECT 71.785 160.015 71.955 160.185 ;
        RECT 72.245 160.015 72.415 160.185 ;
        RECT 72.705 160.015 72.875 160.185 ;
        RECT 73.165 160.015 73.335 160.185 ;
        RECT 73.625 160.015 73.795 160.185 ;
        RECT 74.085 160.015 74.255 160.185 ;
        RECT 74.545 160.015 74.715 160.185 ;
        RECT 75.005 160.015 75.175 160.185 ;
        RECT 75.465 160.015 75.635 160.185 ;
        RECT 75.925 160.015 76.095 160.185 ;
        RECT 76.385 160.015 76.555 160.185 ;
        RECT 76.845 160.015 77.015 160.185 ;
        RECT 77.305 160.015 77.475 160.185 ;
        RECT 77.765 160.015 77.935 160.185 ;
        RECT 78.225 160.015 78.395 160.185 ;
        RECT 78.685 160.015 78.855 160.185 ;
        RECT 79.145 160.015 79.315 160.185 ;
        RECT 79.605 160.015 79.775 160.185 ;
        RECT 80.065 160.015 80.235 160.185 ;
        RECT 80.525 160.015 80.695 160.185 ;
        RECT 80.985 160.015 81.155 160.185 ;
        RECT 81.445 160.015 81.615 160.185 ;
        RECT 81.905 160.015 82.075 160.185 ;
        RECT 82.365 160.015 82.535 160.185 ;
        RECT 82.825 160.015 82.995 160.185 ;
        RECT 83.285 160.015 83.455 160.185 ;
        RECT 83.745 160.015 83.915 160.185 ;
        RECT 84.205 160.015 84.375 160.185 ;
        RECT 84.665 160.015 84.835 160.185 ;
        RECT 85.125 160.015 85.295 160.185 ;
        RECT 85.585 160.015 85.755 160.185 ;
        RECT 86.045 160.015 86.215 160.185 ;
        RECT 86.505 160.015 86.675 160.185 ;
        RECT 86.965 160.015 87.135 160.185 ;
        RECT 87.425 160.015 87.595 160.185 ;
        RECT 87.885 160.015 88.055 160.185 ;
        RECT 88.345 160.015 88.515 160.185 ;
        RECT 88.805 160.015 88.975 160.185 ;
        RECT 89.265 160.015 89.435 160.185 ;
        RECT 89.725 160.015 89.895 160.185 ;
        RECT 90.185 160.015 90.355 160.185 ;
        RECT 90.645 160.015 90.815 160.185 ;
        RECT 91.105 160.015 91.275 160.185 ;
        RECT 91.565 160.015 91.735 160.185 ;
        RECT 92.025 160.015 92.195 160.185 ;
        RECT 36.825 158.485 36.995 158.655 ;
        RECT 37.310 158.145 37.480 158.315 ;
        RECT 37.705 158.485 37.875 158.655 ;
        RECT 38.160 158.825 38.330 158.995 ;
        RECT 38.895 158.485 39.065 158.655 ;
        RECT 39.410 158.145 39.580 158.315 ;
        RECT 40.980 158.145 41.150 158.315 ;
        RECT 41.415 158.485 41.585 158.655 ;
        RECT 43.725 157.805 43.895 157.975 ;
        RECT 53.385 159.165 53.555 159.335 ;
        RECT 54.765 158.825 54.935 158.995 ;
        RECT 46.945 158.145 47.115 158.315 ;
        RECT 55.685 157.805 55.855 157.975 ;
        RECT 70.405 159.165 70.575 159.335 ;
        RECT 79.145 158.825 79.315 158.995 ;
        RECT 79.605 158.825 79.775 158.995 ;
        RECT 80.070 158.145 80.240 158.315 ;
        RECT 80.530 159.165 80.700 159.335 ;
        RECT 80.985 158.485 81.155 158.655 ;
        RECT 81.930 159.165 82.100 159.335 ;
        RECT 83.770 159.165 83.940 159.335 ;
        RECT 82.390 158.145 82.560 158.315 ;
        RECT 83.770 158.145 83.940 158.315 ;
        RECT 87.425 157.805 87.595 157.975 ;
        RECT 18.425 157.295 18.595 157.465 ;
        RECT 18.885 157.295 19.055 157.465 ;
        RECT 19.345 157.295 19.515 157.465 ;
        RECT 19.805 157.295 19.975 157.465 ;
        RECT 20.265 157.295 20.435 157.465 ;
        RECT 20.725 157.295 20.895 157.465 ;
        RECT 21.185 157.295 21.355 157.465 ;
        RECT 21.645 157.295 21.815 157.465 ;
        RECT 22.105 157.295 22.275 157.465 ;
        RECT 22.565 157.295 22.735 157.465 ;
        RECT 23.025 157.295 23.195 157.465 ;
        RECT 23.485 157.295 23.655 157.465 ;
        RECT 23.945 157.295 24.115 157.465 ;
        RECT 24.405 157.295 24.575 157.465 ;
        RECT 24.865 157.295 25.035 157.465 ;
        RECT 25.325 157.295 25.495 157.465 ;
        RECT 25.785 157.295 25.955 157.465 ;
        RECT 26.245 157.295 26.415 157.465 ;
        RECT 26.705 157.295 26.875 157.465 ;
        RECT 27.165 157.295 27.335 157.465 ;
        RECT 27.625 157.295 27.795 157.465 ;
        RECT 28.085 157.295 28.255 157.465 ;
        RECT 28.545 157.295 28.715 157.465 ;
        RECT 29.005 157.295 29.175 157.465 ;
        RECT 29.465 157.295 29.635 157.465 ;
        RECT 29.925 157.295 30.095 157.465 ;
        RECT 30.385 157.295 30.555 157.465 ;
        RECT 30.845 157.295 31.015 157.465 ;
        RECT 31.305 157.295 31.475 157.465 ;
        RECT 31.765 157.295 31.935 157.465 ;
        RECT 32.225 157.295 32.395 157.465 ;
        RECT 32.685 157.295 32.855 157.465 ;
        RECT 33.145 157.295 33.315 157.465 ;
        RECT 33.605 157.295 33.775 157.465 ;
        RECT 34.065 157.295 34.235 157.465 ;
        RECT 34.525 157.295 34.695 157.465 ;
        RECT 34.985 157.295 35.155 157.465 ;
        RECT 35.445 157.295 35.615 157.465 ;
        RECT 35.905 157.295 36.075 157.465 ;
        RECT 36.365 157.295 36.535 157.465 ;
        RECT 36.825 157.295 36.995 157.465 ;
        RECT 37.285 157.295 37.455 157.465 ;
        RECT 37.745 157.295 37.915 157.465 ;
        RECT 38.205 157.295 38.375 157.465 ;
        RECT 38.665 157.295 38.835 157.465 ;
        RECT 39.125 157.295 39.295 157.465 ;
        RECT 39.585 157.295 39.755 157.465 ;
        RECT 40.045 157.295 40.215 157.465 ;
        RECT 40.505 157.295 40.675 157.465 ;
        RECT 40.965 157.295 41.135 157.465 ;
        RECT 41.425 157.295 41.595 157.465 ;
        RECT 41.885 157.295 42.055 157.465 ;
        RECT 42.345 157.295 42.515 157.465 ;
        RECT 42.805 157.295 42.975 157.465 ;
        RECT 43.265 157.295 43.435 157.465 ;
        RECT 43.725 157.295 43.895 157.465 ;
        RECT 44.185 157.295 44.355 157.465 ;
        RECT 44.645 157.295 44.815 157.465 ;
        RECT 45.105 157.295 45.275 157.465 ;
        RECT 45.565 157.295 45.735 157.465 ;
        RECT 46.025 157.295 46.195 157.465 ;
        RECT 46.485 157.295 46.655 157.465 ;
        RECT 46.945 157.295 47.115 157.465 ;
        RECT 47.405 157.295 47.575 157.465 ;
        RECT 47.865 157.295 48.035 157.465 ;
        RECT 48.325 157.295 48.495 157.465 ;
        RECT 48.785 157.295 48.955 157.465 ;
        RECT 49.245 157.295 49.415 157.465 ;
        RECT 49.705 157.295 49.875 157.465 ;
        RECT 50.165 157.295 50.335 157.465 ;
        RECT 50.625 157.295 50.795 157.465 ;
        RECT 51.085 157.295 51.255 157.465 ;
        RECT 51.545 157.295 51.715 157.465 ;
        RECT 52.005 157.295 52.175 157.465 ;
        RECT 52.465 157.295 52.635 157.465 ;
        RECT 52.925 157.295 53.095 157.465 ;
        RECT 53.385 157.295 53.555 157.465 ;
        RECT 53.845 157.295 54.015 157.465 ;
        RECT 54.305 157.295 54.475 157.465 ;
        RECT 54.765 157.295 54.935 157.465 ;
        RECT 55.225 157.295 55.395 157.465 ;
        RECT 55.685 157.295 55.855 157.465 ;
        RECT 56.145 157.295 56.315 157.465 ;
        RECT 56.605 157.295 56.775 157.465 ;
        RECT 57.065 157.295 57.235 157.465 ;
        RECT 57.525 157.295 57.695 157.465 ;
        RECT 57.985 157.295 58.155 157.465 ;
        RECT 58.445 157.295 58.615 157.465 ;
        RECT 58.905 157.295 59.075 157.465 ;
        RECT 59.365 157.295 59.535 157.465 ;
        RECT 59.825 157.295 59.995 157.465 ;
        RECT 60.285 157.295 60.455 157.465 ;
        RECT 60.745 157.295 60.915 157.465 ;
        RECT 61.205 157.295 61.375 157.465 ;
        RECT 61.665 157.295 61.835 157.465 ;
        RECT 62.125 157.295 62.295 157.465 ;
        RECT 62.585 157.295 62.755 157.465 ;
        RECT 63.045 157.295 63.215 157.465 ;
        RECT 63.505 157.295 63.675 157.465 ;
        RECT 63.965 157.295 64.135 157.465 ;
        RECT 64.425 157.295 64.595 157.465 ;
        RECT 64.885 157.295 65.055 157.465 ;
        RECT 65.345 157.295 65.515 157.465 ;
        RECT 65.805 157.295 65.975 157.465 ;
        RECT 66.265 157.295 66.435 157.465 ;
        RECT 66.725 157.295 66.895 157.465 ;
        RECT 67.185 157.295 67.355 157.465 ;
        RECT 67.645 157.295 67.815 157.465 ;
        RECT 68.105 157.295 68.275 157.465 ;
        RECT 68.565 157.295 68.735 157.465 ;
        RECT 69.025 157.295 69.195 157.465 ;
        RECT 69.485 157.295 69.655 157.465 ;
        RECT 69.945 157.295 70.115 157.465 ;
        RECT 70.405 157.295 70.575 157.465 ;
        RECT 70.865 157.295 71.035 157.465 ;
        RECT 71.325 157.295 71.495 157.465 ;
        RECT 71.785 157.295 71.955 157.465 ;
        RECT 72.245 157.295 72.415 157.465 ;
        RECT 72.705 157.295 72.875 157.465 ;
        RECT 73.165 157.295 73.335 157.465 ;
        RECT 73.625 157.295 73.795 157.465 ;
        RECT 74.085 157.295 74.255 157.465 ;
        RECT 74.545 157.295 74.715 157.465 ;
        RECT 75.005 157.295 75.175 157.465 ;
        RECT 75.465 157.295 75.635 157.465 ;
        RECT 75.925 157.295 76.095 157.465 ;
        RECT 76.385 157.295 76.555 157.465 ;
        RECT 76.845 157.295 77.015 157.465 ;
        RECT 77.305 157.295 77.475 157.465 ;
        RECT 77.765 157.295 77.935 157.465 ;
        RECT 78.225 157.295 78.395 157.465 ;
        RECT 78.685 157.295 78.855 157.465 ;
        RECT 79.145 157.295 79.315 157.465 ;
        RECT 79.605 157.295 79.775 157.465 ;
        RECT 80.065 157.295 80.235 157.465 ;
        RECT 80.525 157.295 80.695 157.465 ;
        RECT 80.985 157.295 81.155 157.465 ;
        RECT 81.445 157.295 81.615 157.465 ;
        RECT 81.905 157.295 82.075 157.465 ;
        RECT 82.365 157.295 82.535 157.465 ;
        RECT 82.825 157.295 82.995 157.465 ;
        RECT 83.285 157.295 83.455 157.465 ;
        RECT 83.745 157.295 83.915 157.465 ;
        RECT 84.205 157.295 84.375 157.465 ;
        RECT 84.665 157.295 84.835 157.465 ;
        RECT 85.125 157.295 85.295 157.465 ;
        RECT 85.585 157.295 85.755 157.465 ;
        RECT 86.045 157.295 86.215 157.465 ;
        RECT 86.505 157.295 86.675 157.465 ;
        RECT 86.965 157.295 87.135 157.465 ;
        RECT 87.425 157.295 87.595 157.465 ;
        RECT 87.885 157.295 88.055 157.465 ;
        RECT 88.345 157.295 88.515 157.465 ;
        RECT 88.805 157.295 88.975 157.465 ;
        RECT 89.265 157.295 89.435 157.465 ;
        RECT 89.725 157.295 89.895 157.465 ;
        RECT 90.185 157.295 90.355 157.465 ;
        RECT 90.645 157.295 90.815 157.465 ;
        RECT 91.105 157.295 91.275 157.465 ;
        RECT 91.565 157.295 91.735 157.465 ;
        RECT 92.025 157.295 92.195 157.465 ;
        RECT 45.565 156.785 45.735 156.955 ;
        RECT 44.645 155.765 44.815 155.935 ;
        RECT 45.565 155.765 45.735 155.935 ;
        RECT 46.945 155.765 47.115 155.935 ;
        RECT 47.405 155.765 47.575 155.935 ;
        RECT 46.485 155.085 46.655 155.255 ;
        RECT 50.165 156.105 50.335 156.275 ;
        RECT 52.005 156.105 52.175 156.275 ;
        RECT 52.925 155.765 53.095 155.935 ;
        RECT 53.385 155.085 53.555 155.255 ;
        RECT 53.845 155.085 54.015 155.255 ;
        RECT 54.765 155.425 54.935 155.595 ;
        RECT 59.390 156.445 59.560 156.615 ;
        RECT 57.525 155.765 57.695 155.935 ;
        RECT 58.905 156.105 59.075 156.275 ;
        RECT 58.445 155.765 58.615 155.935 ;
        RECT 57.985 155.425 58.155 155.595 ;
        RECT 59.785 156.105 59.955 156.275 ;
        RECT 60.130 155.425 60.300 155.595 ;
        RECT 61.490 156.445 61.660 156.615 ;
        RECT 60.975 156.105 61.145 156.275 ;
        RECT 63.060 156.445 63.230 156.615 ;
        RECT 63.495 156.105 63.665 156.275 ;
        RECT 66.265 156.105 66.435 156.275 ;
        RECT 67.185 155.765 67.355 155.935 ;
        RECT 67.645 155.765 67.815 155.935 ;
        RECT 68.105 156.105 68.275 156.275 ;
        RECT 68.565 156.105 68.735 156.275 ;
        RECT 69.485 155.765 69.655 155.935 ;
        RECT 69.945 155.765 70.115 155.935 ;
        RECT 65.805 155.085 65.975 155.255 ;
        RECT 73.165 155.085 73.335 155.255 ;
        RECT 74.545 155.765 74.715 155.935 ;
        RECT 75.005 155.765 75.175 155.935 ;
        RECT 75.465 156.105 75.635 156.275 ;
        RECT 75.925 156.105 76.095 156.275 ;
        RECT 76.845 155.765 77.015 155.935 ;
        RECT 77.305 155.765 77.475 155.935 ;
        RECT 73.625 155.085 73.795 155.255 ;
        RECT 80.525 156.105 80.695 156.275 ;
        RECT 82.365 156.445 82.535 156.615 ;
        RECT 80.985 155.765 81.155 155.935 ;
        RECT 81.445 155.085 81.615 155.255 ;
        RECT 83.285 155.765 83.455 155.935 ;
        RECT 82.365 155.425 82.535 155.595 ;
        RECT 83.745 155.085 83.915 155.255 ;
        RECT 18.425 154.575 18.595 154.745 ;
        RECT 18.885 154.575 19.055 154.745 ;
        RECT 19.345 154.575 19.515 154.745 ;
        RECT 19.805 154.575 19.975 154.745 ;
        RECT 20.265 154.575 20.435 154.745 ;
        RECT 20.725 154.575 20.895 154.745 ;
        RECT 21.185 154.575 21.355 154.745 ;
        RECT 21.645 154.575 21.815 154.745 ;
        RECT 22.105 154.575 22.275 154.745 ;
        RECT 22.565 154.575 22.735 154.745 ;
        RECT 23.025 154.575 23.195 154.745 ;
        RECT 23.485 154.575 23.655 154.745 ;
        RECT 23.945 154.575 24.115 154.745 ;
        RECT 24.405 154.575 24.575 154.745 ;
        RECT 24.865 154.575 25.035 154.745 ;
        RECT 25.325 154.575 25.495 154.745 ;
        RECT 25.785 154.575 25.955 154.745 ;
        RECT 26.245 154.575 26.415 154.745 ;
        RECT 26.705 154.575 26.875 154.745 ;
        RECT 27.165 154.575 27.335 154.745 ;
        RECT 27.625 154.575 27.795 154.745 ;
        RECT 28.085 154.575 28.255 154.745 ;
        RECT 28.545 154.575 28.715 154.745 ;
        RECT 29.005 154.575 29.175 154.745 ;
        RECT 29.465 154.575 29.635 154.745 ;
        RECT 29.925 154.575 30.095 154.745 ;
        RECT 30.385 154.575 30.555 154.745 ;
        RECT 30.845 154.575 31.015 154.745 ;
        RECT 31.305 154.575 31.475 154.745 ;
        RECT 31.765 154.575 31.935 154.745 ;
        RECT 32.225 154.575 32.395 154.745 ;
        RECT 32.685 154.575 32.855 154.745 ;
        RECT 33.145 154.575 33.315 154.745 ;
        RECT 33.605 154.575 33.775 154.745 ;
        RECT 34.065 154.575 34.235 154.745 ;
        RECT 34.525 154.575 34.695 154.745 ;
        RECT 34.985 154.575 35.155 154.745 ;
        RECT 35.445 154.575 35.615 154.745 ;
        RECT 35.905 154.575 36.075 154.745 ;
        RECT 36.365 154.575 36.535 154.745 ;
        RECT 36.825 154.575 36.995 154.745 ;
        RECT 37.285 154.575 37.455 154.745 ;
        RECT 37.745 154.575 37.915 154.745 ;
        RECT 38.205 154.575 38.375 154.745 ;
        RECT 38.665 154.575 38.835 154.745 ;
        RECT 39.125 154.575 39.295 154.745 ;
        RECT 39.585 154.575 39.755 154.745 ;
        RECT 40.045 154.575 40.215 154.745 ;
        RECT 40.505 154.575 40.675 154.745 ;
        RECT 40.965 154.575 41.135 154.745 ;
        RECT 41.425 154.575 41.595 154.745 ;
        RECT 41.885 154.575 42.055 154.745 ;
        RECT 42.345 154.575 42.515 154.745 ;
        RECT 42.805 154.575 42.975 154.745 ;
        RECT 43.265 154.575 43.435 154.745 ;
        RECT 43.725 154.575 43.895 154.745 ;
        RECT 44.185 154.575 44.355 154.745 ;
        RECT 44.645 154.575 44.815 154.745 ;
        RECT 45.105 154.575 45.275 154.745 ;
        RECT 45.565 154.575 45.735 154.745 ;
        RECT 46.025 154.575 46.195 154.745 ;
        RECT 46.485 154.575 46.655 154.745 ;
        RECT 46.945 154.575 47.115 154.745 ;
        RECT 47.405 154.575 47.575 154.745 ;
        RECT 47.865 154.575 48.035 154.745 ;
        RECT 48.325 154.575 48.495 154.745 ;
        RECT 48.785 154.575 48.955 154.745 ;
        RECT 49.245 154.575 49.415 154.745 ;
        RECT 49.705 154.575 49.875 154.745 ;
        RECT 50.165 154.575 50.335 154.745 ;
        RECT 50.625 154.575 50.795 154.745 ;
        RECT 51.085 154.575 51.255 154.745 ;
        RECT 51.545 154.575 51.715 154.745 ;
        RECT 52.005 154.575 52.175 154.745 ;
        RECT 52.465 154.575 52.635 154.745 ;
        RECT 52.925 154.575 53.095 154.745 ;
        RECT 53.385 154.575 53.555 154.745 ;
        RECT 53.845 154.575 54.015 154.745 ;
        RECT 54.305 154.575 54.475 154.745 ;
        RECT 54.765 154.575 54.935 154.745 ;
        RECT 55.225 154.575 55.395 154.745 ;
        RECT 55.685 154.575 55.855 154.745 ;
        RECT 56.145 154.575 56.315 154.745 ;
        RECT 56.605 154.575 56.775 154.745 ;
        RECT 57.065 154.575 57.235 154.745 ;
        RECT 57.525 154.575 57.695 154.745 ;
        RECT 57.985 154.575 58.155 154.745 ;
        RECT 58.445 154.575 58.615 154.745 ;
        RECT 58.905 154.575 59.075 154.745 ;
        RECT 59.365 154.575 59.535 154.745 ;
        RECT 59.825 154.575 59.995 154.745 ;
        RECT 60.285 154.575 60.455 154.745 ;
        RECT 60.745 154.575 60.915 154.745 ;
        RECT 61.205 154.575 61.375 154.745 ;
        RECT 61.665 154.575 61.835 154.745 ;
        RECT 62.125 154.575 62.295 154.745 ;
        RECT 62.585 154.575 62.755 154.745 ;
        RECT 63.045 154.575 63.215 154.745 ;
        RECT 63.505 154.575 63.675 154.745 ;
        RECT 63.965 154.575 64.135 154.745 ;
        RECT 64.425 154.575 64.595 154.745 ;
        RECT 64.885 154.575 65.055 154.745 ;
        RECT 65.345 154.575 65.515 154.745 ;
        RECT 65.805 154.575 65.975 154.745 ;
        RECT 66.265 154.575 66.435 154.745 ;
        RECT 66.725 154.575 66.895 154.745 ;
        RECT 67.185 154.575 67.355 154.745 ;
        RECT 67.645 154.575 67.815 154.745 ;
        RECT 68.105 154.575 68.275 154.745 ;
        RECT 68.565 154.575 68.735 154.745 ;
        RECT 69.025 154.575 69.195 154.745 ;
        RECT 69.485 154.575 69.655 154.745 ;
        RECT 69.945 154.575 70.115 154.745 ;
        RECT 70.405 154.575 70.575 154.745 ;
        RECT 70.865 154.575 71.035 154.745 ;
        RECT 71.325 154.575 71.495 154.745 ;
        RECT 71.785 154.575 71.955 154.745 ;
        RECT 72.245 154.575 72.415 154.745 ;
        RECT 72.705 154.575 72.875 154.745 ;
        RECT 73.165 154.575 73.335 154.745 ;
        RECT 73.625 154.575 73.795 154.745 ;
        RECT 74.085 154.575 74.255 154.745 ;
        RECT 74.545 154.575 74.715 154.745 ;
        RECT 75.005 154.575 75.175 154.745 ;
        RECT 75.465 154.575 75.635 154.745 ;
        RECT 75.925 154.575 76.095 154.745 ;
        RECT 76.385 154.575 76.555 154.745 ;
        RECT 76.845 154.575 77.015 154.745 ;
        RECT 77.305 154.575 77.475 154.745 ;
        RECT 77.765 154.575 77.935 154.745 ;
        RECT 78.225 154.575 78.395 154.745 ;
        RECT 78.685 154.575 78.855 154.745 ;
        RECT 79.145 154.575 79.315 154.745 ;
        RECT 79.605 154.575 79.775 154.745 ;
        RECT 80.065 154.575 80.235 154.745 ;
        RECT 80.525 154.575 80.695 154.745 ;
        RECT 80.985 154.575 81.155 154.745 ;
        RECT 81.445 154.575 81.615 154.745 ;
        RECT 81.905 154.575 82.075 154.745 ;
        RECT 82.365 154.575 82.535 154.745 ;
        RECT 82.825 154.575 82.995 154.745 ;
        RECT 83.285 154.575 83.455 154.745 ;
        RECT 83.745 154.575 83.915 154.745 ;
        RECT 84.205 154.575 84.375 154.745 ;
        RECT 84.665 154.575 84.835 154.745 ;
        RECT 85.125 154.575 85.295 154.745 ;
        RECT 85.585 154.575 85.755 154.745 ;
        RECT 86.045 154.575 86.215 154.745 ;
        RECT 86.505 154.575 86.675 154.745 ;
        RECT 86.965 154.575 87.135 154.745 ;
        RECT 87.425 154.575 87.595 154.745 ;
        RECT 87.885 154.575 88.055 154.745 ;
        RECT 88.345 154.575 88.515 154.745 ;
        RECT 88.805 154.575 88.975 154.745 ;
        RECT 89.265 154.575 89.435 154.745 ;
        RECT 89.725 154.575 89.895 154.745 ;
        RECT 90.185 154.575 90.355 154.745 ;
        RECT 90.645 154.575 90.815 154.745 ;
        RECT 91.105 154.575 91.275 154.745 ;
        RECT 91.565 154.575 91.735 154.745 ;
        RECT 92.025 154.575 92.195 154.745 ;
        RECT 41.885 153.385 42.055 153.555 ;
        RECT 42.805 153.725 42.975 153.895 ;
        RECT 46.485 154.065 46.655 154.235 ;
        RECT 43.265 153.385 43.435 153.555 ;
        RECT 41.885 152.365 42.055 152.535 ;
        RECT 47.405 153.385 47.575 153.555 ;
        RECT 48.325 153.045 48.495 153.215 ;
        RECT 48.785 153.385 48.955 153.555 ;
        RECT 47.865 152.705 48.035 152.875 ;
        RECT 49.705 153.385 49.875 153.555 ;
        RECT 53.385 154.065 53.555 154.235 ;
        RECT 51.545 153.385 51.715 153.555 ;
        RECT 52.925 153.385 53.095 153.555 ;
        RECT 50.165 152.365 50.335 152.535 ;
        RECT 51.545 152.365 51.715 152.535 ;
        RECT 54.305 153.385 54.475 153.555 ;
        RECT 54.765 153.725 54.935 153.895 ;
        RECT 55.225 153.385 55.395 153.555 ;
        RECT 56.605 154.065 56.775 154.235 ;
        RECT 56.145 153.045 56.315 153.215 ;
        RECT 57.525 153.385 57.695 153.555 ;
        RECT 58.445 153.045 58.615 153.215 ;
        RECT 67.645 154.065 67.815 154.235 ;
        RECT 66.265 153.385 66.435 153.555 ;
        RECT 67.185 153.385 67.355 153.555 ;
        RECT 67.185 152.705 67.355 152.875 ;
        RECT 68.485 153.725 68.655 153.895 ;
        RECT 69.485 153.725 69.655 153.895 ;
        RECT 68.565 152.365 68.735 152.535 ;
        RECT 70.405 153.045 70.575 153.215 ;
        RECT 71.325 153.725 71.495 153.895 ;
        RECT 71.785 154.065 71.955 154.235 ;
        RECT 72.245 154.065 72.415 154.235 ;
        RECT 74.085 153.385 74.255 153.555 ;
        RECT 73.165 152.705 73.335 152.875 ;
        RECT 75.465 153.385 75.635 153.555 ;
        RECT 74.545 152.705 74.715 152.875 ;
        RECT 75.950 152.705 76.120 152.875 ;
        RECT 76.345 153.045 76.515 153.215 ;
        RECT 76.690 153.725 76.860 153.895 ;
        RECT 77.535 153.045 77.705 153.215 ;
        RECT 78.050 152.705 78.220 152.875 ;
        RECT 79.620 152.705 79.790 152.875 ;
        RECT 80.055 153.045 80.225 153.215 ;
        RECT 82.365 154.065 82.535 154.235 ;
        RECT 18.425 151.855 18.595 152.025 ;
        RECT 18.885 151.855 19.055 152.025 ;
        RECT 19.345 151.855 19.515 152.025 ;
        RECT 19.805 151.855 19.975 152.025 ;
        RECT 20.265 151.855 20.435 152.025 ;
        RECT 20.725 151.855 20.895 152.025 ;
        RECT 21.185 151.855 21.355 152.025 ;
        RECT 21.645 151.855 21.815 152.025 ;
        RECT 22.105 151.855 22.275 152.025 ;
        RECT 22.565 151.855 22.735 152.025 ;
        RECT 23.025 151.855 23.195 152.025 ;
        RECT 23.485 151.855 23.655 152.025 ;
        RECT 23.945 151.855 24.115 152.025 ;
        RECT 24.405 151.855 24.575 152.025 ;
        RECT 24.865 151.855 25.035 152.025 ;
        RECT 25.325 151.855 25.495 152.025 ;
        RECT 25.785 151.855 25.955 152.025 ;
        RECT 26.245 151.855 26.415 152.025 ;
        RECT 26.705 151.855 26.875 152.025 ;
        RECT 27.165 151.855 27.335 152.025 ;
        RECT 27.625 151.855 27.795 152.025 ;
        RECT 28.085 151.855 28.255 152.025 ;
        RECT 28.545 151.855 28.715 152.025 ;
        RECT 29.005 151.855 29.175 152.025 ;
        RECT 29.465 151.855 29.635 152.025 ;
        RECT 29.925 151.855 30.095 152.025 ;
        RECT 30.385 151.855 30.555 152.025 ;
        RECT 30.845 151.855 31.015 152.025 ;
        RECT 31.305 151.855 31.475 152.025 ;
        RECT 31.765 151.855 31.935 152.025 ;
        RECT 32.225 151.855 32.395 152.025 ;
        RECT 32.685 151.855 32.855 152.025 ;
        RECT 33.145 151.855 33.315 152.025 ;
        RECT 33.605 151.855 33.775 152.025 ;
        RECT 34.065 151.855 34.235 152.025 ;
        RECT 34.525 151.855 34.695 152.025 ;
        RECT 34.985 151.855 35.155 152.025 ;
        RECT 35.445 151.855 35.615 152.025 ;
        RECT 35.905 151.855 36.075 152.025 ;
        RECT 36.365 151.855 36.535 152.025 ;
        RECT 36.825 151.855 36.995 152.025 ;
        RECT 37.285 151.855 37.455 152.025 ;
        RECT 37.745 151.855 37.915 152.025 ;
        RECT 38.205 151.855 38.375 152.025 ;
        RECT 38.665 151.855 38.835 152.025 ;
        RECT 39.125 151.855 39.295 152.025 ;
        RECT 39.585 151.855 39.755 152.025 ;
        RECT 40.045 151.855 40.215 152.025 ;
        RECT 40.505 151.855 40.675 152.025 ;
        RECT 40.965 151.855 41.135 152.025 ;
        RECT 41.425 151.855 41.595 152.025 ;
        RECT 41.885 151.855 42.055 152.025 ;
        RECT 42.345 151.855 42.515 152.025 ;
        RECT 42.805 151.855 42.975 152.025 ;
        RECT 43.265 151.855 43.435 152.025 ;
        RECT 43.725 151.855 43.895 152.025 ;
        RECT 44.185 151.855 44.355 152.025 ;
        RECT 44.645 151.855 44.815 152.025 ;
        RECT 45.105 151.855 45.275 152.025 ;
        RECT 45.565 151.855 45.735 152.025 ;
        RECT 46.025 151.855 46.195 152.025 ;
        RECT 46.485 151.855 46.655 152.025 ;
        RECT 46.945 151.855 47.115 152.025 ;
        RECT 47.405 151.855 47.575 152.025 ;
        RECT 47.865 151.855 48.035 152.025 ;
        RECT 48.325 151.855 48.495 152.025 ;
        RECT 48.785 151.855 48.955 152.025 ;
        RECT 49.245 151.855 49.415 152.025 ;
        RECT 49.705 151.855 49.875 152.025 ;
        RECT 50.165 151.855 50.335 152.025 ;
        RECT 50.625 151.855 50.795 152.025 ;
        RECT 51.085 151.855 51.255 152.025 ;
        RECT 51.545 151.855 51.715 152.025 ;
        RECT 52.005 151.855 52.175 152.025 ;
        RECT 52.465 151.855 52.635 152.025 ;
        RECT 52.925 151.855 53.095 152.025 ;
        RECT 53.385 151.855 53.555 152.025 ;
        RECT 53.845 151.855 54.015 152.025 ;
        RECT 54.305 151.855 54.475 152.025 ;
        RECT 54.765 151.855 54.935 152.025 ;
        RECT 55.225 151.855 55.395 152.025 ;
        RECT 55.685 151.855 55.855 152.025 ;
        RECT 56.145 151.855 56.315 152.025 ;
        RECT 56.605 151.855 56.775 152.025 ;
        RECT 57.065 151.855 57.235 152.025 ;
        RECT 57.525 151.855 57.695 152.025 ;
        RECT 57.985 151.855 58.155 152.025 ;
        RECT 58.445 151.855 58.615 152.025 ;
        RECT 58.905 151.855 59.075 152.025 ;
        RECT 59.365 151.855 59.535 152.025 ;
        RECT 59.825 151.855 59.995 152.025 ;
        RECT 60.285 151.855 60.455 152.025 ;
        RECT 60.745 151.855 60.915 152.025 ;
        RECT 61.205 151.855 61.375 152.025 ;
        RECT 61.665 151.855 61.835 152.025 ;
        RECT 62.125 151.855 62.295 152.025 ;
        RECT 62.585 151.855 62.755 152.025 ;
        RECT 63.045 151.855 63.215 152.025 ;
        RECT 63.505 151.855 63.675 152.025 ;
        RECT 63.965 151.855 64.135 152.025 ;
        RECT 64.425 151.855 64.595 152.025 ;
        RECT 64.885 151.855 65.055 152.025 ;
        RECT 65.345 151.855 65.515 152.025 ;
        RECT 65.805 151.855 65.975 152.025 ;
        RECT 66.265 151.855 66.435 152.025 ;
        RECT 66.725 151.855 66.895 152.025 ;
        RECT 67.185 151.855 67.355 152.025 ;
        RECT 67.645 151.855 67.815 152.025 ;
        RECT 68.105 151.855 68.275 152.025 ;
        RECT 68.565 151.855 68.735 152.025 ;
        RECT 69.025 151.855 69.195 152.025 ;
        RECT 69.485 151.855 69.655 152.025 ;
        RECT 69.945 151.855 70.115 152.025 ;
        RECT 70.405 151.855 70.575 152.025 ;
        RECT 70.865 151.855 71.035 152.025 ;
        RECT 71.325 151.855 71.495 152.025 ;
        RECT 71.785 151.855 71.955 152.025 ;
        RECT 72.245 151.855 72.415 152.025 ;
        RECT 72.705 151.855 72.875 152.025 ;
        RECT 73.165 151.855 73.335 152.025 ;
        RECT 73.625 151.855 73.795 152.025 ;
        RECT 74.085 151.855 74.255 152.025 ;
        RECT 74.545 151.855 74.715 152.025 ;
        RECT 75.005 151.855 75.175 152.025 ;
        RECT 75.465 151.855 75.635 152.025 ;
        RECT 75.925 151.855 76.095 152.025 ;
        RECT 76.385 151.855 76.555 152.025 ;
        RECT 76.845 151.855 77.015 152.025 ;
        RECT 77.305 151.855 77.475 152.025 ;
        RECT 77.765 151.855 77.935 152.025 ;
        RECT 78.225 151.855 78.395 152.025 ;
        RECT 78.685 151.855 78.855 152.025 ;
        RECT 79.145 151.855 79.315 152.025 ;
        RECT 79.605 151.855 79.775 152.025 ;
        RECT 80.065 151.855 80.235 152.025 ;
        RECT 80.525 151.855 80.695 152.025 ;
        RECT 80.985 151.855 81.155 152.025 ;
        RECT 81.445 151.855 81.615 152.025 ;
        RECT 81.905 151.855 82.075 152.025 ;
        RECT 82.365 151.855 82.535 152.025 ;
        RECT 82.825 151.855 82.995 152.025 ;
        RECT 83.285 151.855 83.455 152.025 ;
        RECT 83.745 151.855 83.915 152.025 ;
        RECT 84.205 151.855 84.375 152.025 ;
        RECT 84.665 151.855 84.835 152.025 ;
        RECT 85.125 151.855 85.295 152.025 ;
        RECT 85.585 151.855 85.755 152.025 ;
        RECT 86.045 151.855 86.215 152.025 ;
        RECT 86.505 151.855 86.675 152.025 ;
        RECT 86.965 151.855 87.135 152.025 ;
        RECT 87.425 151.855 87.595 152.025 ;
        RECT 87.885 151.855 88.055 152.025 ;
        RECT 88.345 151.855 88.515 152.025 ;
        RECT 88.805 151.855 88.975 152.025 ;
        RECT 89.265 151.855 89.435 152.025 ;
        RECT 89.725 151.855 89.895 152.025 ;
        RECT 90.185 151.855 90.355 152.025 ;
        RECT 90.645 151.855 90.815 152.025 ;
        RECT 91.105 151.855 91.275 152.025 ;
        RECT 91.565 151.855 91.735 152.025 ;
        RECT 92.025 151.855 92.195 152.025 ;
        RECT 37.310 151.005 37.480 151.175 ;
        RECT 36.825 150.325 36.995 150.495 ;
        RECT 37.705 150.665 37.875 150.835 ;
        RECT 38.160 150.325 38.330 150.495 ;
        RECT 39.410 151.005 39.580 151.175 ;
        RECT 38.895 150.665 39.065 150.835 ;
        RECT 40.980 151.005 41.150 151.175 ;
        RECT 41.415 150.665 41.585 150.835 ;
        RECT 43.725 151.005 43.895 151.175 ;
        RECT 45.105 150.665 45.275 150.835 ;
        RECT 48.785 151.345 48.955 151.515 ;
        RECT 50.165 151.345 50.335 151.515 ;
        RECT 47.865 150.325 48.035 150.495 ;
        RECT 48.325 150.325 48.495 150.495 ;
        RECT 49.200 150.325 49.370 150.495 ;
        RECT 51.085 150.325 51.255 150.495 ;
        RECT 51.545 150.325 51.715 150.495 ;
        RECT 52.005 150.325 52.175 150.495 ;
        RECT 52.465 150.665 52.635 150.835 ;
        RECT 60.285 151.005 60.455 151.175 ;
        RECT 60.285 149.985 60.455 150.155 ;
        RECT 61.665 150.325 61.835 150.495 ;
        RECT 62.125 150.325 62.295 150.495 ;
        RECT 63.045 150.325 63.215 150.495 ;
        RECT 61.205 149.645 61.375 149.815 ;
        RECT 62.585 149.645 62.755 149.815 ;
        RECT 70.865 150.665 71.035 150.835 ;
        RECT 70.405 150.325 70.575 150.495 ;
        RECT 72.245 149.645 72.415 149.815 ;
        RECT 74.085 151.345 74.255 151.515 ;
        RECT 74.085 150.325 74.255 150.495 ;
        RECT 75.005 150.325 75.175 150.495 ;
        RECT 18.425 149.135 18.595 149.305 ;
        RECT 18.885 149.135 19.055 149.305 ;
        RECT 19.345 149.135 19.515 149.305 ;
        RECT 19.805 149.135 19.975 149.305 ;
        RECT 20.265 149.135 20.435 149.305 ;
        RECT 20.725 149.135 20.895 149.305 ;
        RECT 21.185 149.135 21.355 149.305 ;
        RECT 21.645 149.135 21.815 149.305 ;
        RECT 22.105 149.135 22.275 149.305 ;
        RECT 22.565 149.135 22.735 149.305 ;
        RECT 23.025 149.135 23.195 149.305 ;
        RECT 23.485 149.135 23.655 149.305 ;
        RECT 23.945 149.135 24.115 149.305 ;
        RECT 24.405 149.135 24.575 149.305 ;
        RECT 24.865 149.135 25.035 149.305 ;
        RECT 25.325 149.135 25.495 149.305 ;
        RECT 25.785 149.135 25.955 149.305 ;
        RECT 26.245 149.135 26.415 149.305 ;
        RECT 26.705 149.135 26.875 149.305 ;
        RECT 27.165 149.135 27.335 149.305 ;
        RECT 27.625 149.135 27.795 149.305 ;
        RECT 28.085 149.135 28.255 149.305 ;
        RECT 28.545 149.135 28.715 149.305 ;
        RECT 29.005 149.135 29.175 149.305 ;
        RECT 29.465 149.135 29.635 149.305 ;
        RECT 29.925 149.135 30.095 149.305 ;
        RECT 30.385 149.135 30.555 149.305 ;
        RECT 30.845 149.135 31.015 149.305 ;
        RECT 31.305 149.135 31.475 149.305 ;
        RECT 31.765 149.135 31.935 149.305 ;
        RECT 32.225 149.135 32.395 149.305 ;
        RECT 32.685 149.135 32.855 149.305 ;
        RECT 33.145 149.135 33.315 149.305 ;
        RECT 33.605 149.135 33.775 149.305 ;
        RECT 34.065 149.135 34.235 149.305 ;
        RECT 34.525 149.135 34.695 149.305 ;
        RECT 34.985 149.135 35.155 149.305 ;
        RECT 35.445 149.135 35.615 149.305 ;
        RECT 35.905 149.135 36.075 149.305 ;
        RECT 36.365 149.135 36.535 149.305 ;
        RECT 36.825 149.135 36.995 149.305 ;
        RECT 37.285 149.135 37.455 149.305 ;
        RECT 37.745 149.135 37.915 149.305 ;
        RECT 38.205 149.135 38.375 149.305 ;
        RECT 38.665 149.135 38.835 149.305 ;
        RECT 39.125 149.135 39.295 149.305 ;
        RECT 39.585 149.135 39.755 149.305 ;
        RECT 40.045 149.135 40.215 149.305 ;
        RECT 40.505 149.135 40.675 149.305 ;
        RECT 40.965 149.135 41.135 149.305 ;
        RECT 41.425 149.135 41.595 149.305 ;
        RECT 41.885 149.135 42.055 149.305 ;
        RECT 42.345 149.135 42.515 149.305 ;
        RECT 42.805 149.135 42.975 149.305 ;
        RECT 43.265 149.135 43.435 149.305 ;
        RECT 43.725 149.135 43.895 149.305 ;
        RECT 44.185 149.135 44.355 149.305 ;
        RECT 44.645 149.135 44.815 149.305 ;
        RECT 45.105 149.135 45.275 149.305 ;
        RECT 45.565 149.135 45.735 149.305 ;
        RECT 46.025 149.135 46.195 149.305 ;
        RECT 46.485 149.135 46.655 149.305 ;
        RECT 46.945 149.135 47.115 149.305 ;
        RECT 47.405 149.135 47.575 149.305 ;
        RECT 47.865 149.135 48.035 149.305 ;
        RECT 48.325 149.135 48.495 149.305 ;
        RECT 48.785 149.135 48.955 149.305 ;
        RECT 49.245 149.135 49.415 149.305 ;
        RECT 49.705 149.135 49.875 149.305 ;
        RECT 50.165 149.135 50.335 149.305 ;
        RECT 50.625 149.135 50.795 149.305 ;
        RECT 51.085 149.135 51.255 149.305 ;
        RECT 51.545 149.135 51.715 149.305 ;
        RECT 52.005 149.135 52.175 149.305 ;
        RECT 52.465 149.135 52.635 149.305 ;
        RECT 52.925 149.135 53.095 149.305 ;
        RECT 53.385 149.135 53.555 149.305 ;
        RECT 53.845 149.135 54.015 149.305 ;
        RECT 54.305 149.135 54.475 149.305 ;
        RECT 54.765 149.135 54.935 149.305 ;
        RECT 55.225 149.135 55.395 149.305 ;
        RECT 55.685 149.135 55.855 149.305 ;
        RECT 56.145 149.135 56.315 149.305 ;
        RECT 56.605 149.135 56.775 149.305 ;
        RECT 57.065 149.135 57.235 149.305 ;
        RECT 57.525 149.135 57.695 149.305 ;
        RECT 57.985 149.135 58.155 149.305 ;
        RECT 58.445 149.135 58.615 149.305 ;
        RECT 58.905 149.135 59.075 149.305 ;
        RECT 59.365 149.135 59.535 149.305 ;
        RECT 59.825 149.135 59.995 149.305 ;
        RECT 60.285 149.135 60.455 149.305 ;
        RECT 60.745 149.135 60.915 149.305 ;
        RECT 61.205 149.135 61.375 149.305 ;
        RECT 61.665 149.135 61.835 149.305 ;
        RECT 62.125 149.135 62.295 149.305 ;
        RECT 62.585 149.135 62.755 149.305 ;
        RECT 63.045 149.135 63.215 149.305 ;
        RECT 63.505 149.135 63.675 149.305 ;
        RECT 63.965 149.135 64.135 149.305 ;
        RECT 64.425 149.135 64.595 149.305 ;
        RECT 64.885 149.135 65.055 149.305 ;
        RECT 65.345 149.135 65.515 149.305 ;
        RECT 65.805 149.135 65.975 149.305 ;
        RECT 66.265 149.135 66.435 149.305 ;
        RECT 66.725 149.135 66.895 149.305 ;
        RECT 67.185 149.135 67.355 149.305 ;
        RECT 67.645 149.135 67.815 149.305 ;
        RECT 68.105 149.135 68.275 149.305 ;
        RECT 68.565 149.135 68.735 149.305 ;
        RECT 69.025 149.135 69.195 149.305 ;
        RECT 69.485 149.135 69.655 149.305 ;
        RECT 69.945 149.135 70.115 149.305 ;
        RECT 70.405 149.135 70.575 149.305 ;
        RECT 70.865 149.135 71.035 149.305 ;
        RECT 71.325 149.135 71.495 149.305 ;
        RECT 71.785 149.135 71.955 149.305 ;
        RECT 72.245 149.135 72.415 149.305 ;
        RECT 72.705 149.135 72.875 149.305 ;
        RECT 73.165 149.135 73.335 149.305 ;
        RECT 73.625 149.135 73.795 149.305 ;
        RECT 74.085 149.135 74.255 149.305 ;
        RECT 74.545 149.135 74.715 149.305 ;
        RECT 75.005 149.135 75.175 149.305 ;
        RECT 75.465 149.135 75.635 149.305 ;
        RECT 75.925 149.135 76.095 149.305 ;
        RECT 76.385 149.135 76.555 149.305 ;
        RECT 76.845 149.135 77.015 149.305 ;
        RECT 77.305 149.135 77.475 149.305 ;
        RECT 77.765 149.135 77.935 149.305 ;
        RECT 78.225 149.135 78.395 149.305 ;
        RECT 78.685 149.135 78.855 149.305 ;
        RECT 79.145 149.135 79.315 149.305 ;
        RECT 79.605 149.135 79.775 149.305 ;
        RECT 80.065 149.135 80.235 149.305 ;
        RECT 80.525 149.135 80.695 149.305 ;
        RECT 80.985 149.135 81.155 149.305 ;
        RECT 81.445 149.135 81.615 149.305 ;
        RECT 81.905 149.135 82.075 149.305 ;
        RECT 82.365 149.135 82.535 149.305 ;
        RECT 82.825 149.135 82.995 149.305 ;
        RECT 83.285 149.135 83.455 149.305 ;
        RECT 83.745 149.135 83.915 149.305 ;
        RECT 84.205 149.135 84.375 149.305 ;
        RECT 84.665 149.135 84.835 149.305 ;
        RECT 85.125 149.135 85.295 149.305 ;
        RECT 85.585 149.135 85.755 149.305 ;
        RECT 86.045 149.135 86.215 149.305 ;
        RECT 86.505 149.135 86.675 149.305 ;
        RECT 86.965 149.135 87.135 149.305 ;
        RECT 87.425 149.135 87.595 149.305 ;
        RECT 87.885 149.135 88.055 149.305 ;
        RECT 88.345 149.135 88.515 149.305 ;
        RECT 88.805 149.135 88.975 149.305 ;
        RECT 89.265 149.135 89.435 149.305 ;
        RECT 89.725 149.135 89.895 149.305 ;
        RECT 90.185 149.135 90.355 149.305 ;
        RECT 90.645 149.135 90.815 149.305 ;
        RECT 91.105 149.135 91.275 149.305 ;
        RECT 91.565 149.135 91.735 149.305 ;
        RECT 92.025 149.135 92.195 149.305 ;
        RECT 54.305 148.285 54.475 148.455 ;
        RECT 56.145 148.625 56.315 148.795 ;
        RECT 53.845 147.945 54.015 148.115 ;
        RECT 54.805 147.945 54.975 148.115 ;
        RECT 55.685 147.945 55.855 148.115 ;
        RECT 56.605 147.945 56.775 148.115 ;
        RECT 57.065 147.945 57.235 148.115 ;
        RECT 63.505 148.625 63.675 148.795 ;
        RECT 65.345 148.625 65.515 148.795 ;
        RECT 60.745 147.945 60.915 148.115 ;
        RECT 62.585 147.945 62.755 148.115 ;
        RECT 61.205 146.925 61.375 147.095 ;
        RECT 65.805 148.285 65.975 148.455 ;
        RECT 73.165 147.945 73.335 148.115 ;
        RECT 70.405 146.925 70.575 147.095 ;
        RECT 73.625 147.605 73.795 147.775 ;
        RECT 18.425 146.415 18.595 146.585 ;
        RECT 18.885 146.415 19.055 146.585 ;
        RECT 19.345 146.415 19.515 146.585 ;
        RECT 19.805 146.415 19.975 146.585 ;
        RECT 20.265 146.415 20.435 146.585 ;
        RECT 20.725 146.415 20.895 146.585 ;
        RECT 21.185 146.415 21.355 146.585 ;
        RECT 21.645 146.415 21.815 146.585 ;
        RECT 22.105 146.415 22.275 146.585 ;
        RECT 22.565 146.415 22.735 146.585 ;
        RECT 23.025 146.415 23.195 146.585 ;
        RECT 23.485 146.415 23.655 146.585 ;
        RECT 23.945 146.415 24.115 146.585 ;
        RECT 24.405 146.415 24.575 146.585 ;
        RECT 24.865 146.415 25.035 146.585 ;
        RECT 25.325 146.415 25.495 146.585 ;
        RECT 25.785 146.415 25.955 146.585 ;
        RECT 26.245 146.415 26.415 146.585 ;
        RECT 26.705 146.415 26.875 146.585 ;
        RECT 27.165 146.415 27.335 146.585 ;
        RECT 27.625 146.415 27.795 146.585 ;
        RECT 28.085 146.415 28.255 146.585 ;
        RECT 28.545 146.415 28.715 146.585 ;
        RECT 29.005 146.415 29.175 146.585 ;
        RECT 29.465 146.415 29.635 146.585 ;
        RECT 29.925 146.415 30.095 146.585 ;
        RECT 30.385 146.415 30.555 146.585 ;
        RECT 30.845 146.415 31.015 146.585 ;
        RECT 31.305 146.415 31.475 146.585 ;
        RECT 31.765 146.415 31.935 146.585 ;
        RECT 32.225 146.415 32.395 146.585 ;
        RECT 32.685 146.415 32.855 146.585 ;
        RECT 33.145 146.415 33.315 146.585 ;
        RECT 33.605 146.415 33.775 146.585 ;
        RECT 34.065 146.415 34.235 146.585 ;
        RECT 34.525 146.415 34.695 146.585 ;
        RECT 34.985 146.415 35.155 146.585 ;
        RECT 35.445 146.415 35.615 146.585 ;
        RECT 35.905 146.415 36.075 146.585 ;
        RECT 36.365 146.415 36.535 146.585 ;
        RECT 36.825 146.415 36.995 146.585 ;
        RECT 37.285 146.415 37.455 146.585 ;
        RECT 37.745 146.415 37.915 146.585 ;
        RECT 38.205 146.415 38.375 146.585 ;
        RECT 38.665 146.415 38.835 146.585 ;
        RECT 39.125 146.415 39.295 146.585 ;
        RECT 39.585 146.415 39.755 146.585 ;
        RECT 40.045 146.415 40.215 146.585 ;
        RECT 40.505 146.415 40.675 146.585 ;
        RECT 40.965 146.415 41.135 146.585 ;
        RECT 41.425 146.415 41.595 146.585 ;
        RECT 41.885 146.415 42.055 146.585 ;
        RECT 42.345 146.415 42.515 146.585 ;
        RECT 42.805 146.415 42.975 146.585 ;
        RECT 43.265 146.415 43.435 146.585 ;
        RECT 43.725 146.415 43.895 146.585 ;
        RECT 44.185 146.415 44.355 146.585 ;
        RECT 44.645 146.415 44.815 146.585 ;
        RECT 45.105 146.415 45.275 146.585 ;
        RECT 45.565 146.415 45.735 146.585 ;
        RECT 46.025 146.415 46.195 146.585 ;
        RECT 46.485 146.415 46.655 146.585 ;
        RECT 46.945 146.415 47.115 146.585 ;
        RECT 47.405 146.415 47.575 146.585 ;
        RECT 47.865 146.415 48.035 146.585 ;
        RECT 48.325 146.415 48.495 146.585 ;
        RECT 48.785 146.415 48.955 146.585 ;
        RECT 49.245 146.415 49.415 146.585 ;
        RECT 49.705 146.415 49.875 146.585 ;
        RECT 50.165 146.415 50.335 146.585 ;
        RECT 50.625 146.415 50.795 146.585 ;
        RECT 51.085 146.415 51.255 146.585 ;
        RECT 51.545 146.415 51.715 146.585 ;
        RECT 52.005 146.415 52.175 146.585 ;
        RECT 52.465 146.415 52.635 146.585 ;
        RECT 52.925 146.415 53.095 146.585 ;
        RECT 53.385 146.415 53.555 146.585 ;
        RECT 53.845 146.415 54.015 146.585 ;
        RECT 54.305 146.415 54.475 146.585 ;
        RECT 54.765 146.415 54.935 146.585 ;
        RECT 55.225 146.415 55.395 146.585 ;
        RECT 55.685 146.415 55.855 146.585 ;
        RECT 56.145 146.415 56.315 146.585 ;
        RECT 56.605 146.415 56.775 146.585 ;
        RECT 57.065 146.415 57.235 146.585 ;
        RECT 57.525 146.415 57.695 146.585 ;
        RECT 57.985 146.415 58.155 146.585 ;
        RECT 58.445 146.415 58.615 146.585 ;
        RECT 58.905 146.415 59.075 146.585 ;
        RECT 59.365 146.415 59.535 146.585 ;
        RECT 59.825 146.415 59.995 146.585 ;
        RECT 60.285 146.415 60.455 146.585 ;
        RECT 60.745 146.415 60.915 146.585 ;
        RECT 61.205 146.415 61.375 146.585 ;
        RECT 61.665 146.415 61.835 146.585 ;
        RECT 62.125 146.415 62.295 146.585 ;
        RECT 62.585 146.415 62.755 146.585 ;
        RECT 63.045 146.415 63.215 146.585 ;
        RECT 63.505 146.415 63.675 146.585 ;
        RECT 63.965 146.415 64.135 146.585 ;
        RECT 64.425 146.415 64.595 146.585 ;
        RECT 64.885 146.415 65.055 146.585 ;
        RECT 65.345 146.415 65.515 146.585 ;
        RECT 65.805 146.415 65.975 146.585 ;
        RECT 66.265 146.415 66.435 146.585 ;
        RECT 66.725 146.415 66.895 146.585 ;
        RECT 67.185 146.415 67.355 146.585 ;
        RECT 67.645 146.415 67.815 146.585 ;
        RECT 68.105 146.415 68.275 146.585 ;
        RECT 68.565 146.415 68.735 146.585 ;
        RECT 69.025 146.415 69.195 146.585 ;
        RECT 69.485 146.415 69.655 146.585 ;
        RECT 69.945 146.415 70.115 146.585 ;
        RECT 70.405 146.415 70.575 146.585 ;
        RECT 70.865 146.415 71.035 146.585 ;
        RECT 71.325 146.415 71.495 146.585 ;
        RECT 71.785 146.415 71.955 146.585 ;
        RECT 72.245 146.415 72.415 146.585 ;
        RECT 72.705 146.415 72.875 146.585 ;
        RECT 73.165 146.415 73.335 146.585 ;
        RECT 73.625 146.415 73.795 146.585 ;
        RECT 74.085 146.415 74.255 146.585 ;
        RECT 74.545 146.415 74.715 146.585 ;
        RECT 75.005 146.415 75.175 146.585 ;
        RECT 75.465 146.415 75.635 146.585 ;
        RECT 75.925 146.415 76.095 146.585 ;
        RECT 76.385 146.415 76.555 146.585 ;
        RECT 76.845 146.415 77.015 146.585 ;
        RECT 77.305 146.415 77.475 146.585 ;
        RECT 77.765 146.415 77.935 146.585 ;
        RECT 78.225 146.415 78.395 146.585 ;
        RECT 78.685 146.415 78.855 146.585 ;
        RECT 79.145 146.415 79.315 146.585 ;
        RECT 79.605 146.415 79.775 146.585 ;
        RECT 80.065 146.415 80.235 146.585 ;
        RECT 80.525 146.415 80.695 146.585 ;
        RECT 80.985 146.415 81.155 146.585 ;
        RECT 81.445 146.415 81.615 146.585 ;
        RECT 81.905 146.415 82.075 146.585 ;
        RECT 82.365 146.415 82.535 146.585 ;
        RECT 82.825 146.415 82.995 146.585 ;
        RECT 83.285 146.415 83.455 146.585 ;
        RECT 83.745 146.415 83.915 146.585 ;
        RECT 84.205 146.415 84.375 146.585 ;
        RECT 84.665 146.415 84.835 146.585 ;
        RECT 85.125 146.415 85.295 146.585 ;
        RECT 85.585 146.415 85.755 146.585 ;
        RECT 86.045 146.415 86.215 146.585 ;
        RECT 86.505 146.415 86.675 146.585 ;
        RECT 86.965 146.415 87.135 146.585 ;
        RECT 87.425 146.415 87.595 146.585 ;
        RECT 87.885 146.415 88.055 146.585 ;
        RECT 88.345 146.415 88.515 146.585 ;
        RECT 88.805 146.415 88.975 146.585 ;
        RECT 89.265 146.415 89.435 146.585 ;
        RECT 89.725 146.415 89.895 146.585 ;
        RECT 90.185 146.415 90.355 146.585 ;
        RECT 90.645 146.415 90.815 146.585 ;
        RECT 91.105 146.415 91.275 146.585 ;
        RECT 91.565 146.415 91.735 146.585 ;
        RECT 92.025 146.415 92.195 146.585 ;
        RECT 43.290 145.565 43.460 145.735 ;
        RECT 42.805 145.225 42.975 145.395 ;
        RECT 43.685 145.225 43.855 145.395 ;
        RECT 44.140 144.545 44.310 144.715 ;
        RECT 45.390 145.565 45.560 145.735 ;
        RECT 44.875 145.225 45.045 145.395 ;
        RECT 46.960 145.565 47.130 145.735 ;
        RECT 47.395 145.225 47.565 145.395 ;
        RECT 50.790 144.885 50.960 145.055 ;
        RECT 49.705 144.205 49.875 144.375 ;
        RECT 50.165 144.205 50.335 144.375 ;
        RECT 52.925 145.225 53.095 145.395 ;
        RECT 53.845 145.225 54.015 145.395 ;
        RECT 53.385 144.885 53.555 145.055 ;
        RECT 55.225 145.225 55.395 145.395 ;
        RECT 55.685 144.885 55.855 145.055 ;
        RECT 57.525 145.905 57.695 146.075 ;
        RECT 59.835 145.225 60.005 145.395 ;
        RECT 60.270 145.565 60.440 145.735 ;
        RECT 61.840 145.565 62.010 145.735 ;
        RECT 62.355 145.225 62.525 145.395 ;
        RECT 63.090 144.885 63.260 145.055 ;
        RECT 63.545 145.225 63.715 145.395 ;
        RECT 63.940 145.565 64.110 145.735 ;
        RECT 65.830 145.565 66.000 145.735 ;
        RECT 64.425 144.885 64.595 145.055 ;
        RECT 65.345 144.885 65.515 145.055 ;
        RECT 66.225 145.225 66.395 145.395 ;
        RECT 66.680 144.545 66.850 144.715 ;
        RECT 67.930 145.565 68.100 145.735 ;
        RECT 67.415 145.225 67.585 145.395 ;
        RECT 69.500 145.565 69.670 145.735 ;
        RECT 69.935 145.225 70.105 145.395 ;
        RECT 72.245 145.905 72.415 146.075 ;
        RECT 18.425 143.695 18.595 143.865 ;
        RECT 18.885 143.695 19.055 143.865 ;
        RECT 19.345 143.695 19.515 143.865 ;
        RECT 19.805 143.695 19.975 143.865 ;
        RECT 20.265 143.695 20.435 143.865 ;
        RECT 20.725 143.695 20.895 143.865 ;
        RECT 21.185 143.695 21.355 143.865 ;
        RECT 21.645 143.695 21.815 143.865 ;
        RECT 22.105 143.695 22.275 143.865 ;
        RECT 22.565 143.695 22.735 143.865 ;
        RECT 23.025 143.695 23.195 143.865 ;
        RECT 23.485 143.695 23.655 143.865 ;
        RECT 23.945 143.695 24.115 143.865 ;
        RECT 24.405 143.695 24.575 143.865 ;
        RECT 24.865 143.695 25.035 143.865 ;
        RECT 25.325 143.695 25.495 143.865 ;
        RECT 25.785 143.695 25.955 143.865 ;
        RECT 26.245 143.695 26.415 143.865 ;
        RECT 26.705 143.695 26.875 143.865 ;
        RECT 27.165 143.695 27.335 143.865 ;
        RECT 27.625 143.695 27.795 143.865 ;
        RECT 28.085 143.695 28.255 143.865 ;
        RECT 28.545 143.695 28.715 143.865 ;
        RECT 29.005 143.695 29.175 143.865 ;
        RECT 29.465 143.695 29.635 143.865 ;
        RECT 29.925 143.695 30.095 143.865 ;
        RECT 30.385 143.695 30.555 143.865 ;
        RECT 30.845 143.695 31.015 143.865 ;
        RECT 31.305 143.695 31.475 143.865 ;
        RECT 31.765 143.695 31.935 143.865 ;
        RECT 32.225 143.695 32.395 143.865 ;
        RECT 32.685 143.695 32.855 143.865 ;
        RECT 33.145 143.695 33.315 143.865 ;
        RECT 33.605 143.695 33.775 143.865 ;
        RECT 34.065 143.695 34.235 143.865 ;
        RECT 34.525 143.695 34.695 143.865 ;
        RECT 34.985 143.695 35.155 143.865 ;
        RECT 35.445 143.695 35.615 143.865 ;
        RECT 35.905 143.695 36.075 143.865 ;
        RECT 36.365 143.695 36.535 143.865 ;
        RECT 36.825 143.695 36.995 143.865 ;
        RECT 37.285 143.695 37.455 143.865 ;
        RECT 37.745 143.695 37.915 143.865 ;
        RECT 38.205 143.695 38.375 143.865 ;
        RECT 38.665 143.695 38.835 143.865 ;
        RECT 39.125 143.695 39.295 143.865 ;
        RECT 39.585 143.695 39.755 143.865 ;
        RECT 40.045 143.695 40.215 143.865 ;
        RECT 40.505 143.695 40.675 143.865 ;
        RECT 40.965 143.695 41.135 143.865 ;
        RECT 41.425 143.695 41.595 143.865 ;
        RECT 41.885 143.695 42.055 143.865 ;
        RECT 42.345 143.695 42.515 143.865 ;
        RECT 42.805 143.695 42.975 143.865 ;
        RECT 43.265 143.695 43.435 143.865 ;
        RECT 43.725 143.695 43.895 143.865 ;
        RECT 44.185 143.695 44.355 143.865 ;
        RECT 44.645 143.695 44.815 143.865 ;
        RECT 45.105 143.695 45.275 143.865 ;
        RECT 45.565 143.695 45.735 143.865 ;
        RECT 46.025 143.695 46.195 143.865 ;
        RECT 46.485 143.695 46.655 143.865 ;
        RECT 46.945 143.695 47.115 143.865 ;
        RECT 47.405 143.695 47.575 143.865 ;
        RECT 47.865 143.695 48.035 143.865 ;
        RECT 48.325 143.695 48.495 143.865 ;
        RECT 48.785 143.695 48.955 143.865 ;
        RECT 49.245 143.695 49.415 143.865 ;
        RECT 49.705 143.695 49.875 143.865 ;
        RECT 50.165 143.695 50.335 143.865 ;
        RECT 50.625 143.695 50.795 143.865 ;
        RECT 51.085 143.695 51.255 143.865 ;
        RECT 51.545 143.695 51.715 143.865 ;
        RECT 52.005 143.695 52.175 143.865 ;
        RECT 52.465 143.695 52.635 143.865 ;
        RECT 52.925 143.695 53.095 143.865 ;
        RECT 53.385 143.695 53.555 143.865 ;
        RECT 53.845 143.695 54.015 143.865 ;
        RECT 54.305 143.695 54.475 143.865 ;
        RECT 54.765 143.695 54.935 143.865 ;
        RECT 55.225 143.695 55.395 143.865 ;
        RECT 55.685 143.695 55.855 143.865 ;
        RECT 56.145 143.695 56.315 143.865 ;
        RECT 56.605 143.695 56.775 143.865 ;
        RECT 57.065 143.695 57.235 143.865 ;
        RECT 57.525 143.695 57.695 143.865 ;
        RECT 57.985 143.695 58.155 143.865 ;
        RECT 58.445 143.695 58.615 143.865 ;
        RECT 58.905 143.695 59.075 143.865 ;
        RECT 59.365 143.695 59.535 143.865 ;
        RECT 59.825 143.695 59.995 143.865 ;
        RECT 60.285 143.695 60.455 143.865 ;
        RECT 60.745 143.695 60.915 143.865 ;
        RECT 61.205 143.695 61.375 143.865 ;
        RECT 61.665 143.695 61.835 143.865 ;
        RECT 62.125 143.695 62.295 143.865 ;
        RECT 62.585 143.695 62.755 143.865 ;
        RECT 63.045 143.695 63.215 143.865 ;
        RECT 63.505 143.695 63.675 143.865 ;
        RECT 63.965 143.695 64.135 143.865 ;
        RECT 64.425 143.695 64.595 143.865 ;
        RECT 64.885 143.695 65.055 143.865 ;
        RECT 65.345 143.695 65.515 143.865 ;
        RECT 65.805 143.695 65.975 143.865 ;
        RECT 66.265 143.695 66.435 143.865 ;
        RECT 66.725 143.695 66.895 143.865 ;
        RECT 67.185 143.695 67.355 143.865 ;
        RECT 67.645 143.695 67.815 143.865 ;
        RECT 68.105 143.695 68.275 143.865 ;
        RECT 68.565 143.695 68.735 143.865 ;
        RECT 69.025 143.695 69.195 143.865 ;
        RECT 69.485 143.695 69.655 143.865 ;
        RECT 69.945 143.695 70.115 143.865 ;
        RECT 70.405 143.695 70.575 143.865 ;
        RECT 70.865 143.695 71.035 143.865 ;
        RECT 71.325 143.695 71.495 143.865 ;
        RECT 71.785 143.695 71.955 143.865 ;
        RECT 72.245 143.695 72.415 143.865 ;
        RECT 72.705 143.695 72.875 143.865 ;
        RECT 73.165 143.695 73.335 143.865 ;
        RECT 73.625 143.695 73.795 143.865 ;
        RECT 74.085 143.695 74.255 143.865 ;
        RECT 74.545 143.695 74.715 143.865 ;
        RECT 75.005 143.695 75.175 143.865 ;
        RECT 75.465 143.695 75.635 143.865 ;
        RECT 75.925 143.695 76.095 143.865 ;
        RECT 76.385 143.695 76.555 143.865 ;
        RECT 76.845 143.695 77.015 143.865 ;
        RECT 77.305 143.695 77.475 143.865 ;
        RECT 77.765 143.695 77.935 143.865 ;
        RECT 78.225 143.695 78.395 143.865 ;
        RECT 78.685 143.695 78.855 143.865 ;
        RECT 79.145 143.695 79.315 143.865 ;
        RECT 79.605 143.695 79.775 143.865 ;
        RECT 80.065 143.695 80.235 143.865 ;
        RECT 80.525 143.695 80.695 143.865 ;
        RECT 80.985 143.695 81.155 143.865 ;
        RECT 81.445 143.695 81.615 143.865 ;
        RECT 81.905 143.695 82.075 143.865 ;
        RECT 82.365 143.695 82.535 143.865 ;
        RECT 82.825 143.695 82.995 143.865 ;
        RECT 83.285 143.695 83.455 143.865 ;
        RECT 83.745 143.695 83.915 143.865 ;
        RECT 84.205 143.695 84.375 143.865 ;
        RECT 84.665 143.695 84.835 143.865 ;
        RECT 85.125 143.695 85.295 143.865 ;
        RECT 85.585 143.695 85.755 143.865 ;
        RECT 86.045 143.695 86.215 143.865 ;
        RECT 86.505 143.695 86.675 143.865 ;
        RECT 86.965 143.695 87.135 143.865 ;
        RECT 87.425 143.695 87.595 143.865 ;
        RECT 87.885 143.695 88.055 143.865 ;
        RECT 88.345 143.695 88.515 143.865 ;
        RECT 88.805 143.695 88.975 143.865 ;
        RECT 89.265 143.695 89.435 143.865 ;
        RECT 89.725 143.695 89.895 143.865 ;
        RECT 90.185 143.695 90.355 143.865 ;
        RECT 90.645 143.695 90.815 143.865 ;
        RECT 91.105 143.695 91.275 143.865 ;
        RECT 91.565 143.695 91.735 143.865 ;
        RECT 92.025 143.695 92.195 143.865 ;
        RECT 45.105 143.185 45.275 143.355 ;
        RECT 44.645 142.505 44.815 142.675 ;
        RECT 45.565 142.505 45.735 142.675 ;
        RECT 67.185 143.185 67.355 143.355 ;
        RECT 66.725 142.505 66.895 142.675 ;
        RECT 67.645 142.505 67.815 142.675 ;
        RECT 18.425 140.975 18.595 141.145 ;
        RECT 18.885 140.975 19.055 141.145 ;
        RECT 19.345 140.975 19.515 141.145 ;
        RECT 19.805 140.975 19.975 141.145 ;
        RECT 20.265 140.975 20.435 141.145 ;
        RECT 20.725 140.975 20.895 141.145 ;
        RECT 21.185 140.975 21.355 141.145 ;
        RECT 21.645 140.975 21.815 141.145 ;
        RECT 22.105 140.975 22.275 141.145 ;
        RECT 22.565 140.975 22.735 141.145 ;
        RECT 23.025 140.975 23.195 141.145 ;
        RECT 23.485 140.975 23.655 141.145 ;
        RECT 23.945 140.975 24.115 141.145 ;
        RECT 24.405 140.975 24.575 141.145 ;
        RECT 24.865 140.975 25.035 141.145 ;
        RECT 25.325 140.975 25.495 141.145 ;
        RECT 25.785 140.975 25.955 141.145 ;
        RECT 26.245 140.975 26.415 141.145 ;
        RECT 26.705 140.975 26.875 141.145 ;
        RECT 27.165 140.975 27.335 141.145 ;
        RECT 27.625 140.975 27.795 141.145 ;
        RECT 28.085 140.975 28.255 141.145 ;
        RECT 28.545 140.975 28.715 141.145 ;
        RECT 29.005 140.975 29.175 141.145 ;
        RECT 29.465 140.975 29.635 141.145 ;
        RECT 29.925 140.975 30.095 141.145 ;
        RECT 30.385 140.975 30.555 141.145 ;
        RECT 30.845 140.975 31.015 141.145 ;
        RECT 31.305 140.975 31.475 141.145 ;
        RECT 31.765 140.975 31.935 141.145 ;
        RECT 32.225 140.975 32.395 141.145 ;
        RECT 32.685 140.975 32.855 141.145 ;
        RECT 33.145 140.975 33.315 141.145 ;
        RECT 33.605 140.975 33.775 141.145 ;
        RECT 34.065 140.975 34.235 141.145 ;
        RECT 34.525 140.975 34.695 141.145 ;
        RECT 34.985 140.975 35.155 141.145 ;
        RECT 35.445 140.975 35.615 141.145 ;
        RECT 35.905 140.975 36.075 141.145 ;
        RECT 36.365 140.975 36.535 141.145 ;
        RECT 36.825 140.975 36.995 141.145 ;
        RECT 37.285 140.975 37.455 141.145 ;
        RECT 37.745 140.975 37.915 141.145 ;
        RECT 38.205 140.975 38.375 141.145 ;
        RECT 38.665 140.975 38.835 141.145 ;
        RECT 39.125 140.975 39.295 141.145 ;
        RECT 39.585 140.975 39.755 141.145 ;
        RECT 40.045 140.975 40.215 141.145 ;
        RECT 40.505 140.975 40.675 141.145 ;
        RECT 40.965 140.975 41.135 141.145 ;
        RECT 41.425 140.975 41.595 141.145 ;
        RECT 41.885 140.975 42.055 141.145 ;
        RECT 42.345 140.975 42.515 141.145 ;
        RECT 42.805 140.975 42.975 141.145 ;
        RECT 43.265 140.975 43.435 141.145 ;
        RECT 43.725 140.975 43.895 141.145 ;
        RECT 44.185 140.975 44.355 141.145 ;
        RECT 44.645 140.975 44.815 141.145 ;
        RECT 45.105 140.975 45.275 141.145 ;
        RECT 45.565 140.975 45.735 141.145 ;
        RECT 46.025 140.975 46.195 141.145 ;
        RECT 46.485 140.975 46.655 141.145 ;
        RECT 46.945 140.975 47.115 141.145 ;
        RECT 47.405 140.975 47.575 141.145 ;
        RECT 47.865 140.975 48.035 141.145 ;
        RECT 48.325 140.975 48.495 141.145 ;
        RECT 48.785 140.975 48.955 141.145 ;
        RECT 49.245 140.975 49.415 141.145 ;
        RECT 49.705 140.975 49.875 141.145 ;
        RECT 50.165 140.975 50.335 141.145 ;
        RECT 50.625 140.975 50.795 141.145 ;
        RECT 51.085 140.975 51.255 141.145 ;
        RECT 51.545 140.975 51.715 141.145 ;
        RECT 52.005 140.975 52.175 141.145 ;
        RECT 52.465 140.975 52.635 141.145 ;
        RECT 52.925 140.975 53.095 141.145 ;
        RECT 53.385 140.975 53.555 141.145 ;
        RECT 53.845 140.975 54.015 141.145 ;
        RECT 54.305 140.975 54.475 141.145 ;
        RECT 54.765 140.975 54.935 141.145 ;
        RECT 55.225 140.975 55.395 141.145 ;
        RECT 55.685 140.975 55.855 141.145 ;
        RECT 56.145 140.975 56.315 141.145 ;
        RECT 56.605 140.975 56.775 141.145 ;
        RECT 57.065 140.975 57.235 141.145 ;
        RECT 57.525 140.975 57.695 141.145 ;
        RECT 57.985 140.975 58.155 141.145 ;
        RECT 58.445 140.975 58.615 141.145 ;
        RECT 58.905 140.975 59.075 141.145 ;
        RECT 59.365 140.975 59.535 141.145 ;
        RECT 59.825 140.975 59.995 141.145 ;
        RECT 60.285 140.975 60.455 141.145 ;
        RECT 60.745 140.975 60.915 141.145 ;
        RECT 61.205 140.975 61.375 141.145 ;
        RECT 61.665 140.975 61.835 141.145 ;
        RECT 62.125 140.975 62.295 141.145 ;
        RECT 62.585 140.975 62.755 141.145 ;
        RECT 63.045 140.975 63.215 141.145 ;
        RECT 63.505 140.975 63.675 141.145 ;
        RECT 63.965 140.975 64.135 141.145 ;
        RECT 64.425 140.975 64.595 141.145 ;
        RECT 64.885 140.975 65.055 141.145 ;
        RECT 65.345 140.975 65.515 141.145 ;
        RECT 65.805 140.975 65.975 141.145 ;
        RECT 66.265 140.975 66.435 141.145 ;
        RECT 66.725 140.975 66.895 141.145 ;
        RECT 67.185 140.975 67.355 141.145 ;
        RECT 67.645 140.975 67.815 141.145 ;
        RECT 68.105 140.975 68.275 141.145 ;
        RECT 68.565 140.975 68.735 141.145 ;
        RECT 69.025 140.975 69.195 141.145 ;
        RECT 69.485 140.975 69.655 141.145 ;
        RECT 69.945 140.975 70.115 141.145 ;
        RECT 70.405 140.975 70.575 141.145 ;
        RECT 70.865 140.975 71.035 141.145 ;
        RECT 71.325 140.975 71.495 141.145 ;
        RECT 71.785 140.975 71.955 141.145 ;
        RECT 72.245 140.975 72.415 141.145 ;
        RECT 72.705 140.975 72.875 141.145 ;
        RECT 73.165 140.975 73.335 141.145 ;
        RECT 73.625 140.975 73.795 141.145 ;
        RECT 74.085 140.975 74.255 141.145 ;
        RECT 74.545 140.975 74.715 141.145 ;
        RECT 75.005 140.975 75.175 141.145 ;
        RECT 75.465 140.975 75.635 141.145 ;
        RECT 75.925 140.975 76.095 141.145 ;
        RECT 76.385 140.975 76.555 141.145 ;
        RECT 76.845 140.975 77.015 141.145 ;
        RECT 77.305 140.975 77.475 141.145 ;
        RECT 77.765 140.975 77.935 141.145 ;
        RECT 78.225 140.975 78.395 141.145 ;
        RECT 78.685 140.975 78.855 141.145 ;
        RECT 79.145 140.975 79.315 141.145 ;
        RECT 79.605 140.975 79.775 141.145 ;
        RECT 80.065 140.975 80.235 141.145 ;
        RECT 80.525 140.975 80.695 141.145 ;
        RECT 80.985 140.975 81.155 141.145 ;
        RECT 81.445 140.975 81.615 141.145 ;
        RECT 81.905 140.975 82.075 141.145 ;
        RECT 82.365 140.975 82.535 141.145 ;
        RECT 82.825 140.975 82.995 141.145 ;
        RECT 83.285 140.975 83.455 141.145 ;
        RECT 83.745 140.975 83.915 141.145 ;
        RECT 84.205 140.975 84.375 141.145 ;
        RECT 84.665 140.975 84.835 141.145 ;
        RECT 85.125 140.975 85.295 141.145 ;
        RECT 85.585 140.975 85.755 141.145 ;
        RECT 86.045 140.975 86.215 141.145 ;
        RECT 86.505 140.975 86.675 141.145 ;
        RECT 86.965 140.975 87.135 141.145 ;
        RECT 87.425 140.975 87.595 141.145 ;
        RECT 87.885 140.975 88.055 141.145 ;
        RECT 88.345 140.975 88.515 141.145 ;
        RECT 88.805 140.975 88.975 141.145 ;
        RECT 89.265 140.975 89.435 141.145 ;
        RECT 89.725 140.975 89.895 141.145 ;
        RECT 90.185 140.975 90.355 141.145 ;
        RECT 90.645 140.975 90.815 141.145 ;
        RECT 91.105 140.975 91.275 141.145 ;
        RECT 91.565 140.975 91.735 141.145 ;
        RECT 92.025 140.975 92.195 141.145 ;
        RECT 18.425 138.255 18.595 138.425 ;
        RECT 18.885 138.255 19.055 138.425 ;
        RECT 19.345 138.255 19.515 138.425 ;
        RECT 19.805 138.255 19.975 138.425 ;
        RECT 20.265 138.255 20.435 138.425 ;
        RECT 20.725 138.255 20.895 138.425 ;
        RECT 21.185 138.255 21.355 138.425 ;
        RECT 21.645 138.255 21.815 138.425 ;
        RECT 22.105 138.255 22.275 138.425 ;
        RECT 22.565 138.255 22.735 138.425 ;
        RECT 23.025 138.255 23.195 138.425 ;
        RECT 23.485 138.255 23.655 138.425 ;
        RECT 23.945 138.255 24.115 138.425 ;
        RECT 24.405 138.255 24.575 138.425 ;
        RECT 24.865 138.255 25.035 138.425 ;
        RECT 25.325 138.255 25.495 138.425 ;
        RECT 25.785 138.255 25.955 138.425 ;
        RECT 26.245 138.255 26.415 138.425 ;
        RECT 26.705 138.255 26.875 138.425 ;
        RECT 27.165 138.255 27.335 138.425 ;
        RECT 27.625 138.255 27.795 138.425 ;
        RECT 28.085 138.255 28.255 138.425 ;
        RECT 28.545 138.255 28.715 138.425 ;
        RECT 29.005 138.255 29.175 138.425 ;
        RECT 29.465 138.255 29.635 138.425 ;
        RECT 29.925 138.255 30.095 138.425 ;
        RECT 30.385 138.255 30.555 138.425 ;
        RECT 30.845 138.255 31.015 138.425 ;
        RECT 31.305 138.255 31.475 138.425 ;
        RECT 31.765 138.255 31.935 138.425 ;
        RECT 32.225 138.255 32.395 138.425 ;
        RECT 32.685 138.255 32.855 138.425 ;
        RECT 33.145 138.255 33.315 138.425 ;
        RECT 33.605 138.255 33.775 138.425 ;
        RECT 34.065 138.255 34.235 138.425 ;
        RECT 34.525 138.255 34.695 138.425 ;
        RECT 34.985 138.255 35.155 138.425 ;
        RECT 35.445 138.255 35.615 138.425 ;
        RECT 35.905 138.255 36.075 138.425 ;
        RECT 36.365 138.255 36.535 138.425 ;
        RECT 36.825 138.255 36.995 138.425 ;
        RECT 37.285 138.255 37.455 138.425 ;
        RECT 37.745 138.255 37.915 138.425 ;
        RECT 38.205 138.255 38.375 138.425 ;
        RECT 38.665 138.255 38.835 138.425 ;
        RECT 39.125 138.255 39.295 138.425 ;
        RECT 39.585 138.255 39.755 138.425 ;
        RECT 40.045 138.255 40.215 138.425 ;
        RECT 40.505 138.255 40.675 138.425 ;
        RECT 40.965 138.255 41.135 138.425 ;
        RECT 41.425 138.255 41.595 138.425 ;
        RECT 41.885 138.255 42.055 138.425 ;
        RECT 42.345 138.255 42.515 138.425 ;
        RECT 42.805 138.255 42.975 138.425 ;
        RECT 43.265 138.255 43.435 138.425 ;
        RECT 43.725 138.255 43.895 138.425 ;
        RECT 44.185 138.255 44.355 138.425 ;
        RECT 44.645 138.255 44.815 138.425 ;
        RECT 45.105 138.255 45.275 138.425 ;
        RECT 45.565 138.255 45.735 138.425 ;
        RECT 46.025 138.255 46.195 138.425 ;
        RECT 46.485 138.255 46.655 138.425 ;
        RECT 46.945 138.255 47.115 138.425 ;
        RECT 47.405 138.255 47.575 138.425 ;
        RECT 47.865 138.255 48.035 138.425 ;
        RECT 48.325 138.255 48.495 138.425 ;
        RECT 48.785 138.255 48.955 138.425 ;
        RECT 49.245 138.255 49.415 138.425 ;
        RECT 49.705 138.255 49.875 138.425 ;
        RECT 50.165 138.255 50.335 138.425 ;
        RECT 50.625 138.255 50.795 138.425 ;
        RECT 51.085 138.255 51.255 138.425 ;
        RECT 51.545 138.255 51.715 138.425 ;
        RECT 52.005 138.255 52.175 138.425 ;
        RECT 52.465 138.255 52.635 138.425 ;
        RECT 52.925 138.255 53.095 138.425 ;
        RECT 53.385 138.255 53.555 138.425 ;
        RECT 53.845 138.255 54.015 138.425 ;
        RECT 54.305 138.255 54.475 138.425 ;
        RECT 54.765 138.255 54.935 138.425 ;
        RECT 55.225 138.255 55.395 138.425 ;
        RECT 55.685 138.255 55.855 138.425 ;
        RECT 56.145 138.255 56.315 138.425 ;
        RECT 56.605 138.255 56.775 138.425 ;
        RECT 57.065 138.255 57.235 138.425 ;
        RECT 57.525 138.255 57.695 138.425 ;
        RECT 57.985 138.255 58.155 138.425 ;
        RECT 58.445 138.255 58.615 138.425 ;
        RECT 58.905 138.255 59.075 138.425 ;
        RECT 59.365 138.255 59.535 138.425 ;
        RECT 59.825 138.255 59.995 138.425 ;
        RECT 60.285 138.255 60.455 138.425 ;
        RECT 60.745 138.255 60.915 138.425 ;
        RECT 61.205 138.255 61.375 138.425 ;
        RECT 61.665 138.255 61.835 138.425 ;
        RECT 62.125 138.255 62.295 138.425 ;
        RECT 62.585 138.255 62.755 138.425 ;
        RECT 63.045 138.255 63.215 138.425 ;
        RECT 63.505 138.255 63.675 138.425 ;
        RECT 63.965 138.255 64.135 138.425 ;
        RECT 64.425 138.255 64.595 138.425 ;
        RECT 64.885 138.255 65.055 138.425 ;
        RECT 65.345 138.255 65.515 138.425 ;
        RECT 65.805 138.255 65.975 138.425 ;
        RECT 66.265 138.255 66.435 138.425 ;
        RECT 66.725 138.255 66.895 138.425 ;
        RECT 67.185 138.255 67.355 138.425 ;
        RECT 67.645 138.255 67.815 138.425 ;
        RECT 68.105 138.255 68.275 138.425 ;
        RECT 68.565 138.255 68.735 138.425 ;
        RECT 69.025 138.255 69.195 138.425 ;
        RECT 69.485 138.255 69.655 138.425 ;
        RECT 69.945 138.255 70.115 138.425 ;
        RECT 70.405 138.255 70.575 138.425 ;
        RECT 70.865 138.255 71.035 138.425 ;
        RECT 71.325 138.255 71.495 138.425 ;
        RECT 71.785 138.255 71.955 138.425 ;
        RECT 72.245 138.255 72.415 138.425 ;
        RECT 72.705 138.255 72.875 138.425 ;
        RECT 73.165 138.255 73.335 138.425 ;
        RECT 73.625 138.255 73.795 138.425 ;
        RECT 74.085 138.255 74.255 138.425 ;
        RECT 74.545 138.255 74.715 138.425 ;
        RECT 75.005 138.255 75.175 138.425 ;
        RECT 75.465 138.255 75.635 138.425 ;
        RECT 75.925 138.255 76.095 138.425 ;
        RECT 76.385 138.255 76.555 138.425 ;
        RECT 76.845 138.255 77.015 138.425 ;
        RECT 77.305 138.255 77.475 138.425 ;
        RECT 77.765 138.255 77.935 138.425 ;
        RECT 78.225 138.255 78.395 138.425 ;
        RECT 78.685 138.255 78.855 138.425 ;
        RECT 79.145 138.255 79.315 138.425 ;
        RECT 79.605 138.255 79.775 138.425 ;
        RECT 80.065 138.255 80.235 138.425 ;
        RECT 80.525 138.255 80.695 138.425 ;
        RECT 80.985 138.255 81.155 138.425 ;
        RECT 81.445 138.255 81.615 138.425 ;
        RECT 81.905 138.255 82.075 138.425 ;
        RECT 82.365 138.255 82.535 138.425 ;
        RECT 82.825 138.255 82.995 138.425 ;
        RECT 83.285 138.255 83.455 138.425 ;
        RECT 83.745 138.255 83.915 138.425 ;
        RECT 84.205 138.255 84.375 138.425 ;
        RECT 84.665 138.255 84.835 138.425 ;
        RECT 85.125 138.255 85.295 138.425 ;
        RECT 85.585 138.255 85.755 138.425 ;
        RECT 86.045 138.255 86.215 138.425 ;
        RECT 86.505 138.255 86.675 138.425 ;
        RECT 86.965 138.255 87.135 138.425 ;
        RECT 87.425 138.255 87.595 138.425 ;
        RECT 87.885 138.255 88.055 138.425 ;
        RECT 88.345 138.255 88.515 138.425 ;
        RECT 88.805 138.255 88.975 138.425 ;
        RECT 89.265 138.255 89.435 138.425 ;
        RECT 89.725 138.255 89.895 138.425 ;
        RECT 90.185 138.255 90.355 138.425 ;
        RECT 90.645 138.255 90.815 138.425 ;
        RECT 91.105 138.255 91.275 138.425 ;
        RECT 91.565 138.255 91.735 138.425 ;
        RECT 92.025 138.255 92.195 138.425 ;
        RECT 18.425 135.535 18.595 135.705 ;
        RECT 18.885 135.535 19.055 135.705 ;
        RECT 19.345 135.535 19.515 135.705 ;
        RECT 19.805 135.535 19.975 135.705 ;
        RECT 20.265 135.535 20.435 135.705 ;
        RECT 20.725 135.535 20.895 135.705 ;
        RECT 21.185 135.535 21.355 135.705 ;
        RECT 21.645 135.535 21.815 135.705 ;
        RECT 22.105 135.535 22.275 135.705 ;
        RECT 22.565 135.535 22.735 135.705 ;
        RECT 23.025 135.535 23.195 135.705 ;
        RECT 23.485 135.535 23.655 135.705 ;
        RECT 23.945 135.535 24.115 135.705 ;
        RECT 24.405 135.535 24.575 135.705 ;
        RECT 24.865 135.535 25.035 135.705 ;
        RECT 25.325 135.535 25.495 135.705 ;
        RECT 25.785 135.535 25.955 135.705 ;
        RECT 26.245 135.535 26.415 135.705 ;
        RECT 26.705 135.535 26.875 135.705 ;
        RECT 27.165 135.535 27.335 135.705 ;
        RECT 27.625 135.535 27.795 135.705 ;
        RECT 28.085 135.535 28.255 135.705 ;
        RECT 28.545 135.535 28.715 135.705 ;
        RECT 29.005 135.535 29.175 135.705 ;
        RECT 29.465 135.535 29.635 135.705 ;
        RECT 29.925 135.535 30.095 135.705 ;
        RECT 30.385 135.535 30.555 135.705 ;
        RECT 30.845 135.535 31.015 135.705 ;
        RECT 31.305 135.535 31.475 135.705 ;
        RECT 31.765 135.535 31.935 135.705 ;
        RECT 32.225 135.535 32.395 135.705 ;
        RECT 32.685 135.535 32.855 135.705 ;
        RECT 33.145 135.535 33.315 135.705 ;
        RECT 33.605 135.535 33.775 135.705 ;
        RECT 34.065 135.535 34.235 135.705 ;
        RECT 34.525 135.535 34.695 135.705 ;
        RECT 34.985 135.535 35.155 135.705 ;
        RECT 35.445 135.535 35.615 135.705 ;
        RECT 35.905 135.535 36.075 135.705 ;
        RECT 36.365 135.535 36.535 135.705 ;
        RECT 36.825 135.535 36.995 135.705 ;
        RECT 37.285 135.535 37.455 135.705 ;
        RECT 37.745 135.535 37.915 135.705 ;
        RECT 38.205 135.535 38.375 135.705 ;
        RECT 38.665 135.535 38.835 135.705 ;
        RECT 39.125 135.535 39.295 135.705 ;
        RECT 39.585 135.535 39.755 135.705 ;
        RECT 40.045 135.535 40.215 135.705 ;
        RECT 40.505 135.535 40.675 135.705 ;
        RECT 40.965 135.535 41.135 135.705 ;
        RECT 41.425 135.535 41.595 135.705 ;
        RECT 41.885 135.535 42.055 135.705 ;
        RECT 42.345 135.535 42.515 135.705 ;
        RECT 42.805 135.535 42.975 135.705 ;
        RECT 43.265 135.535 43.435 135.705 ;
        RECT 43.725 135.535 43.895 135.705 ;
        RECT 44.185 135.535 44.355 135.705 ;
        RECT 44.645 135.535 44.815 135.705 ;
        RECT 45.105 135.535 45.275 135.705 ;
        RECT 45.565 135.535 45.735 135.705 ;
        RECT 46.025 135.535 46.195 135.705 ;
        RECT 46.485 135.535 46.655 135.705 ;
        RECT 46.945 135.535 47.115 135.705 ;
        RECT 47.405 135.535 47.575 135.705 ;
        RECT 47.865 135.535 48.035 135.705 ;
        RECT 48.325 135.535 48.495 135.705 ;
        RECT 48.785 135.535 48.955 135.705 ;
        RECT 49.245 135.535 49.415 135.705 ;
        RECT 49.705 135.535 49.875 135.705 ;
        RECT 50.165 135.535 50.335 135.705 ;
        RECT 50.625 135.535 50.795 135.705 ;
        RECT 51.085 135.535 51.255 135.705 ;
        RECT 51.545 135.535 51.715 135.705 ;
        RECT 52.005 135.535 52.175 135.705 ;
        RECT 52.465 135.535 52.635 135.705 ;
        RECT 52.925 135.535 53.095 135.705 ;
        RECT 53.385 135.535 53.555 135.705 ;
        RECT 53.845 135.535 54.015 135.705 ;
        RECT 54.305 135.535 54.475 135.705 ;
        RECT 54.765 135.535 54.935 135.705 ;
        RECT 55.225 135.535 55.395 135.705 ;
        RECT 55.685 135.535 55.855 135.705 ;
        RECT 56.145 135.535 56.315 135.705 ;
        RECT 56.605 135.535 56.775 135.705 ;
        RECT 57.065 135.535 57.235 135.705 ;
        RECT 57.525 135.535 57.695 135.705 ;
        RECT 57.985 135.535 58.155 135.705 ;
        RECT 58.445 135.535 58.615 135.705 ;
        RECT 58.905 135.535 59.075 135.705 ;
        RECT 59.365 135.535 59.535 135.705 ;
        RECT 59.825 135.535 59.995 135.705 ;
        RECT 60.285 135.535 60.455 135.705 ;
        RECT 60.745 135.535 60.915 135.705 ;
        RECT 61.205 135.535 61.375 135.705 ;
        RECT 61.665 135.535 61.835 135.705 ;
        RECT 62.125 135.535 62.295 135.705 ;
        RECT 62.585 135.535 62.755 135.705 ;
        RECT 63.045 135.535 63.215 135.705 ;
        RECT 63.505 135.535 63.675 135.705 ;
        RECT 63.965 135.535 64.135 135.705 ;
        RECT 64.425 135.535 64.595 135.705 ;
        RECT 64.885 135.535 65.055 135.705 ;
        RECT 65.345 135.535 65.515 135.705 ;
        RECT 65.805 135.535 65.975 135.705 ;
        RECT 66.265 135.535 66.435 135.705 ;
        RECT 66.725 135.535 66.895 135.705 ;
        RECT 67.185 135.535 67.355 135.705 ;
        RECT 67.645 135.535 67.815 135.705 ;
        RECT 68.105 135.535 68.275 135.705 ;
        RECT 68.565 135.535 68.735 135.705 ;
        RECT 69.025 135.535 69.195 135.705 ;
        RECT 69.485 135.535 69.655 135.705 ;
        RECT 69.945 135.535 70.115 135.705 ;
        RECT 70.405 135.535 70.575 135.705 ;
        RECT 70.865 135.535 71.035 135.705 ;
        RECT 71.325 135.535 71.495 135.705 ;
        RECT 71.785 135.535 71.955 135.705 ;
        RECT 72.245 135.535 72.415 135.705 ;
        RECT 72.705 135.535 72.875 135.705 ;
        RECT 73.165 135.535 73.335 135.705 ;
        RECT 73.625 135.535 73.795 135.705 ;
        RECT 74.085 135.535 74.255 135.705 ;
        RECT 74.545 135.535 74.715 135.705 ;
        RECT 75.005 135.535 75.175 135.705 ;
        RECT 75.465 135.535 75.635 135.705 ;
        RECT 75.925 135.535 76.095 135.705 ;
        RECT 76.385 135.535 76.555 135.705 ;
        RECT 76.845 135.535 77.015 135.705 ;
        RECT 77.305 135.535 77.475 135.705 ;
        RECT 77.765 135.535 77.935 135.705 ;
        RECT 78.225 135.535 78.395 135.705 ;
        RECT 78.685 135.535 78.855 135.705 ;
        RECT 79.145 135.535 79.315 135.705 ;
        RECT 79.605 135.535 79.775 135.705 ;
        RECT 80.065 135.535 80.235 135.705 ;
        RECT 80.525 135.535 80.695 135.705 ;
        RECT 80.985 135.535 81.155 135.705 ;
        RECT 81.445 135.535 81.615 135.705 ;
        RECT 81.905 135.535 82.075 135.705 ;
        RECT 82.365 135.535 82.535 135.705 ;
        RECT 82.825 135.535 82.995 135.705 ;
        RECT 83.285 135.535 83.455 135.705 ;
        RECT 83.745 135.535 83.915 135.705 ;
        RECT 84.205 135.535 84.375 135.705 ;
        RECT 84.665 135.535 84.835 135.705 ;
        RECT 85.125 135.535 85.295 135.705 ;
        RECT 85.585 135.535 85.755 135.705 ;
        RECT 86.045 135.535 86.215 135.705 ;
        RECT 86.505 135.535 86.675 135.705 ;
        RECT 86.965 135.535 87.135 135.705 ;
        RECT 87.425 135.535 87.595 135.705 ;
        RECT 87.885 135.535 88.055 135.705 ;
        RECT 88.345 135.535 88.515 135.705 ;
        RECT 88.805 135.535 88.975 135.705 ;
        RECT 89.265 135.535 89.435 135.705 ;
        RECT 89.725 135.535 89.895 135.705 ;
        RECT 90.185 135.535 90.355 135.705 ;
        RECT 90.645 135.535 90.815 135.705 ;
        RECT 91.105 135.535 91.275 135.705 ;
        RECT 91.565 135.535 91.735 135.705 ;
        RECT 92.025 135.535 92.195 135.705 ;
        RECT 18.425 132.815 18.595 132.985 ;
        RECT 18.885 132.815 19.055 132.985 ;
        RECT 19.345 132.815 19.515 132.985 ;
        RECT 19.805 132.815 19.975 132.985 ;
        RECT 20.265 132.815 20.435 132.985 ;
        RECT 20.725 132.815 20.895 132.985 ;
        RECT 21.185 132.815 21.355 132.985 ;
        RECT 21.645 132.815 21.815 132.985 ;
        RECT 22.105 132.815 22.275 132.985 ;
        RECT 22.565 132.815 22.735 132.985 ;
        RECT 23.025 132.815 23.195 132.985 ;
        RECT 23.485 132.815 23.655 132.985 ;
        RECT 23.945 132.815 24.115 132.985 ;
        RECT 24.405 132.815 24.575 132.985 ;
        RECT 24.865 132.815 25.035 132.985 ;
        RECT 25.325 132.815 25.495 132.985 ;
        RECT 25.785 132.815 25.955 132.985 ;
        RECT 26.245 132.815 26.415 132.985 ;
        RECT 26.705 132.815 26.875 132.985 ;
        RECT 27.165 132.815 27.335 132.985 ;
        RECT 27.625 132.815 27.795 132.985 ;
        RECT 28.085 132.815 28.255 132.985 ;
        RECT 28.545 132.815 28.715 132.985 ;
        RECT 29.005 132.815 29.175 132.985 ;
        RECT 29.465 132.815 29.635 132.985 ;
        RECT 29.925 132.815 30.095 132.985 ;
        RECT 30.385 132.815 30.555 132.985 ;
        RECT 30.845 132.815 31.015 132.985 ;
        RECT 31.305 132.815 31.475 132.985 ;
        RECT 31.765 132.815 31.935 132.985 ;
        RECT 32.225 132.815 32.395 132.985 ;
        RECT 32.685 132.815 32.855 132.985 ;
        RECT 33.145 132.815 33.315 132.985 ;
        RECT 33.605 132.815 33.775 132.985 ;
        RECT 34.065 132.815 34.235 132.985 ;
        RECT 34.525 132.815 34.695 132.985 ;
        RECT 34.985 132.815 35.155 132.985 ;
        RECT 35.445 132.815 35.615 132.985 ;
        RECT 35.905 132.815 36.075 132.985 ;
        RECT 36.365 132.815 36.535 132.985 ;
        RECT 36.825 132.815 36.995 132.985 ;
        RECT 37.285 132.815 37.455 132.985 ;
        RECT 37.745 132.815 37.915 132.985 ;
        RECT 38.205 132.815 38.375 132.985 ;
        RECT 38.665 132.815 38.835 132.985 ;
        RECT 39.125 132.815 39.295 132.985 ;
        RECT 39.585 132.815 39.755 132.985 ;
        RECT 40.045 132.815 40.215 132.985 ;
        RECT 40.505 132.815 40.675 132.985 ;
        RECT 40.965 132.815 41.135 132.985 ;
        RECT 41.425 132.815 41.595 132.985 ;
        RECT 41.885 132.815 42.055 132.985 ;
        RECT 42.345 132.815 42.515 132.985 ;
        RECT 42.805 132.815 42.975 132.985 ;
        RECT 43.265 132.815 43.435 132.985 ;
        RECT 43.725 132.815 43.895 132.985 ;
        RECT 44.185 132.815 44.355 132.985 ;
        RECT 44.645 132.815 44.815 132.985 ;
        RECT 45.105 132.815 45.275 132.985 ;
        RECT 45.565 132.815 45.735 132.985 ;
        RECT 46.025 132.815 46.195 132.985 ;
        RECT 46.485 132.815 46.655 132.985 ;
        RECT 46.945 132.815 47.115 132.985 ;
        RECT 47.405 132.815 47.575 132.985 ;
        RECT 47.865 132.815 48.035 132.985 ;
        RECT 48.325 132.815 48.495 132.985 ;
        RECT 48.785 132.815 48.955 132.985 ;
        RECT 49.245 132.815 49.415 132.985 ;
        RECT 49.705 132.815 49.875 132.985 ;
        RECT 50.165 132.815 50.335 132.985 ;
        RECT 50.625 132.815 50.795 132.985 ;
        RECT 51.085 132.815 51.255 132.985 ;
        RECT 51.545 132.815 51.715 132.985 ;
        RECT 52.005 132.815 52.175 132.985 ;
        RECT 52.465 132.815 52.635 132.985 ;
        RECT 52.925 132.815 53.095 132.985 ;
        RECT 53.385 132.815 53.555 132.985 ;
        RECT 53.845 132.815 54.015 132.985 ;
        RECT 54.305 132.815 54.475 132.985 ;
        RECT 54.765 132.815 54.935 132.985 ;
        RECT 55.225 132.815 55.395 132.985 ;
        RECT 55.685 132.815 55.855 132.985 ;
        RECT 56.145 132.815 56.315 132.985 ;
        RECT 56.605 132.815 56.775 132.985 ;
        RECT 57.065 132.815 57.235 132.985 ;
        RECT 57.525 132.815 57.695 132.985 ;
        RECT 57.985 132.815 58.155 132.985 ;
        RECT 58.445 132.815 58.615 132.985 ;
        RECT 58.905 132.815 59.075 132.985 ;
        RECT 59.365 132.815 59.535 132.985 ;
        RECT 59.825 132.815 59.995 132.985 ;
        RECT 60.285 132.815 60.455 132.985 ;
        RECT 60.745 132.815 60.915 132.985 ;
        RECT 61.205 132.815 61.375 132.985 ;
        RECT 61.665 132.815 61.835 132.985 ;
        RECT 62.125 132.815 62.295 132.985 ;
        RECT 62.585 132.815 62.755 132.985 ;
        RECT 63.045 132.815 63.215 132.985 ;
        RECT 63.505 132.815 63.675 132.985 ;
        RECT 63.965 132.815 64.135 132.985 ;
        RECT 64.425 132.815 64.595 132.985 ;
        RECT 64.885 132.815 65.055 132.985 ;
        RECT 65.345 132.815 65.515 132.985 ;
        RECT 65.805 132.815 65.975 132.985 ;
        RECT 66.265 132.815 66.435 132.985 ;
        RECT 66.725 132.815 66.895 132.985 ;
        RECT 67.185 132.815 67.355 132.985 ;
        RECT 67.645 132.815 67.815 132.985 ;
        RECT 68.105 132.815 68.275 132.985 ;
        RECT 68.565 132.815 68.735 132.985 ;
        RECT 69.025 132.815 69.195 132.985 ;
        RECT 69.485 132.815 69.655 132.985 ;
        RECT 69.945 132.815 70.115 132.985 ;
        RECT 70.405 132.815 70.575 132.985 ;
        RECT 70.865 132.815 71.035 132.985 ;
        RECT 71.325 132.815 71.495 132.985 ;
        RECT 71.785 132.815 71.955 132.985 ;
        RECT 72.245 132.815 72.415 132.985 ;
        RECT 72.705 132.815 72.875 132.985 ;
        RECT 73.165 132.815 73.335 132.985 ;
        RECT 73.625 132.815 73.795 132.985 ;
        RECT 74.085 132.815 74.255 132.985 ;
        RECT 74.545 132.815 74.715 132.985 ;
        RECT 75.005 132.815 75.175 132.985 ;
        RECT 75.465 132.815 75.635 132.985 ;
        RECT 75.925 132.815 76.095 132.985 ;
        RECT 76.385 132.815 76.555 132.985 ;
        RECT 76.845 132.815 77.015 132.985 ;
        RECT 77.305 132.815 77.475 132.985 ;
        RECT 77.765 132.815 77.935 132.985 ;
        RECT 78.225 132.815 78.395 132.985 ;
        RECT 78.685 132.815 78.855 132.985 ;
        RECT 79.145 132.815 79.315 132.985 ;
        RECT 79.605 132.815 79.775 132.985 ;
        RECT 80.065 132.815 80.235 132.985 ;
        RECT 80.525 132.815 80.695 132.985 ;
        RECT 80.985 132.815 81.155 132.985 ;
        RECT 81.445 132.815 81.615 132.985 ;
        RECT 81.905 132.815 82.075 132.985 ;
        RECT 82.365 132.815 82.535 132.985 ;
        RECT 82.825 132.815 82.995 132.985 ;
        RECT 83.285 132.815 83.455 132.985 ;
        RECT 83.745 132.815 83.915 132.985 ;
        RECT 84.205 132.815 84.375 132.985 ;
        RECT 84.665 132.815 84.835 132.985 ;
        RECT 85.125 132.815 85.295 132.985 ;
        RECT 85.585 132.815 85.755 132.985 ;
        RECT 86.045 132.815 86.215 132.985 ;
        RECT 86.505 132.815 86.675 132.985 ;
        RECT 86.965 132.815 87.135 132.985 ;
        RECT 87.425 132.815 87.595 132.985 ;
        RECT 87.885 132.815 88.055 132.985 ;
        RECT 88.345 132.815 88.515 132.985 ;
        RECT 88.805 132.815 88.975 132.985 ;
        RECT 89.265 132.815 89.435 132.985 ;
        RECT 89.725 132.815 89.895 132.985 ;
        RECT 90.185 132.815 90.355 132.985 ;
        RECT 90.645 132.815 90.815 132.985 ;
        RECT 91.105 132.815 91.275 132.985 ;
        RECT 91.565 132.815 91.735 132.985 ;
        RECT 92.025 132.815 92.195 132.985 ;
        RECT 106.910 112.075 107.100 114.060 ;
        RECT 106.910 69.920 107.100 71.905 ;
        RECT 110.910 139.075 111.100 141.060 ;
        RECT 110.910 96.920 111.100 98.905 ;
        RECT 113.910 139.075 114.100 141.060 ;
        RECT 113.910 96.920 114.100 98.905 ;
        RECT 116.910 139.075 117.100 141.060 ;
        RECT 116.910 96.920 117.100 98.905 ;
        RECT 119.910 139.075 120.100 141.060 ;
        RECT 119.910 96.920 120.100 98.905 ;
        RECT 122.910 139.075 123.100 141.060 ;
        RECT 122.910 96.920 123.100 98.905 ;
        RECT 125.910 139.075 126.100 141.060 ;
        RECT 125.910 96.920 126.100 98.905 ;
        RECT 128.910 139.075 129.100 141.060 ;
        RECT 128.910 96.920 129.100 98.905 ;
        RECT 131.910 139.075 132.100 141.060 ;
        RECT 131.910 96.920 132.100 98.905 ;
        RECT 110.910 92.075 111.100 94.060 ;
        RECT 110.910 69.920 111.100 71.905 ;
        RECT 113.910 92.075 114.100 94.060 ;
        RECT 113.910 69.920 114.100 71.905 ;
        RECT 116.910 92.075 117.100 94.060 ;
        RECT 116.910 69.920 117.100 71.905 ;
        RECT 119.910 92.075 120.100 94.060 ;
        RECT 119.910 69.920 120.100 71.905 ;
        RECT 122.910 92.075 123.100 94.060 ;
        RECT 122.910 69.920 123.100 71.905 ;
        RECT 125.910 92.075 126.100 94.060 ;
        RECT 125.910 69.920 126.100 71.905 ;
        RECT 128.910 92.075 129.100 94.060 ;
        RECT 128.910 69.920 129.100 71.905 ;
      LAYER met1 ;
        RECT 18.280 206.100 92.340 206.580 ;
        RECT 39.970 205.700 40.290 205.960 ;
        RECT 59.765 205.900 60.055 205.945 ;
        RECT 69.870 205.900 70.190 205.960 ;
        RECT 59.765 205.760 70.190 205.900 ;
        RECT 59.765 205.715 60.055 205.760 ;
        RECT 69.870 205.700 70.190 205.760 ;
        RECT 28.025 205.560 28.315 205.605 ;
        RECT 43.190 205.560 43.510 205.620 ;
        RECT 28.025 205.420 43.510 205.560 ;
        RECT 28.025 205.375 28.315 205.420 ;
        RECT 43.190 205.360 43.510 205.420 ;
        RECT 21.585 205.220 21.875 205.265 ;
        RECT 39.510 205.220 39.830 205.280 ;
        RECT 58.370 205.220 58.690 205.280 ;
        RECT 21.585 205.080 39.280 205.220 ;
        RECT 21.585 205.035 21.875 205.080 ;
        RECT 19.730 204.880 20.050 204.940 ;
        RECT 20.665 204.880 20.955 204.925 ;
        RECT 19.730 204.740 20.955 204.880 ;
        RECT 19.730 204.680 20.050 204.740 ;
        RECT 20.665 204.695 20.955 204.740 ;
        RECT 26.170 204.880 26.490 204.940 ;
        RECT 27.105 204.880 27.395 204.925 ;
        RECT 26.170 204.740 27.395 204.880 ;
        RECT 26.170 204.680 26.490 204.740 ;
        RECT 27.105 204.695 27.395 204.740 ;
        RECT 32.610 204.880 32.930 204.940 ;
        RECT 33.085 204.880 33.375 204.925 ;
        RECT 32.610 204.740 33.375 204.880 ;
        RECT 39.140 204.880 39.280 205.080 ;
        RECT 39.510 205.080 41.580 205.220 ;
        RECT 39.510 205.020 39.830 205.080 ;
        RECT 39.985 204.880 40.275 204.925 ;
        RECT 40.890 204.880 41.210 204.940 ;
        RECT 41.440 204.925 41.580 205.080 ;
        RECT 58.370 205.080 60.900 205.220 ;
        RECT 58.370 205.020 58.690 205.080 ;
        RECT 39.140 204.740 41.210 204.880 ;
        RECT 32.610 204.680 32.930 204.740 ;
        RECT 33.085 204.695 33.375 204.740 ;
        RECT 39.985 204.695 40.275 204.740 ;
        RECT 40.890 204.680 41.210 204.740 ;
        RECT 41.365 204.695 41.655 204.925 ;
        RECT 41.825 204.695 42.115 204.925 ;
        RECT 44.570 204.880 44.890 204.940 ;
        RECT 45.965 204.880 46.255 204.925 ;
        RECT 44.570 204.740 46.255 204.880 ;
        RECT 39.050 204.540 39.370 204.600 ;
        RECT 41.900 204.540 42.040 204.695 ;
        RECT 44.570 204.680 44.890 204.740 ;
        RECT 45.965 204.695 46.255 204.740 ;
        RECT 51.930 204.880 52.250 204.940 ;
        RECT 52.405 204.880 52.695 204.925 ;
        RECT 51.930 204.740 52.695 204.880 ;
        RECT 51.930 204.680 52.250 204.740 ;
        RECT 52.405 204.695 52.695 204.740 ;
        RECT 53.310 204.880 53.630 204.940 ;
        RECT 58.845 204.880 59.135 204.925 ;
        RECT 53.310 204.740 59.135 204.880 ;
        RECT 53.310 204.680 53.630 204.740 ;
        RECT 58.845 204.695 59.135 204.740 ;
        RECT 60.210 204.680 60.530 204.940 ;
        RECT 60.760 204.925 60.900 205.080 ;
        RECT 60.685 204.695 60.975 204.925 ;
        RECT 65.285 204.880 65.575 204.925 ;
        RECT 65.730 204.880 66.050 204.940 ;
        RECT 65.285 204.740 66.050 204.880 ;
        RECT 65.285 204.695 65.575 204.740 ;
        RECT 65.730 204.680 66.050 204.740 ;
        RECT 71.250 204.880 71.570 204.940 ;
        RECT 71.725 204.880 72.015 204.925 ;
        RECT 71.250 204.740 72.015 204.880 ;
        RECT 71.250 204.680 71.570 204.740 ;
        RECT 71.725 204.695 72.015 204.740 ;
        RECT 77.690 204.880 78.010 204.940 ;
        RECT 79.085 204.880 79.375 204.925 ;
        RECT 77.690 204.740 79.375 204.880 ;
        RECT 77.690 204.680 78.010 204.740 ;
        RECT 79.085 204.695 79.375 204.740 ;
        RECT 84.130 204.880 84.450 204.940 ;
        RECT 84.605 204.880 84.895 204.925 ;
        RECT 84.130 204.740 84.895 204.880 ;
        RECT 84.130 204.680 84.450 204.740 ;
        RECT 84.605 204.695 84.895 204.740 ;
        RECT 39.050 204.400 42.040 204.540 ;
        RECT 68.030 204.540 68.350 204.600 ;
        RECT 68.030 204.400 78.380 204.540 ;
        RECT 39.050 204.340 39.370 204.400 ;
        RECT 68.030 204.340 68.350 204.400 ;
        RECT 34.005 204.200 34.295 204.245 ;
        RECT 37.670 204.200 37.990 204.260 ;
        RECT 34.005 204.060 37.990 204.200 ;
        RECT 34.005 204.015 34.295 204.060 ;
        RECT 37.670 204.000 37.990 204.060 ;
        RECT 38.590 204.000 38.910 204.260 ;
        RECT 42.730 204.000 43.050 204.260 ;
        RECT 46.870 204.000 47.190 204.260 ;
        RECT 53.325 204.200 53.615 204.245 ;
        RECT 53.770 204.200 54.090 204.260 ;
        RECT 53.325 204.060 54.090 204.200 ;
        RECT 53.325 204.015 53.615 204.060 ;
        RECT 53.770 204.000 54.090 204.060 ;
        RECT 57.450 204.000 57.770 204.260 ;
        RECT 60.670 204.200 60.990 204.260 ;
        RECT 61.605 204.200 61.895 204.245 ;
        RECT 60.670 204.060 61.895 204.200 ;
        RECT 60.670 204.000 60.990 204.060 ;
        RECT 61.605 204.015 61.895 204.060 ;
        RECT 66.205 204.200 66.495 204.245 ;
        RECT 69.410 204.200 69.730 204.260 ;
        RECT 66.205 204.060 69.730 204.200 ;
        RECT 66.205 204.015 66.495 204.060 ;
        RECT 69.410 204.000 69.730 204.060 ;
        RECT 72.170 204.200 72.490 204.260 ;
        RECT 78.240 204.245 78.380 204.400 ;
        RECT 72.645 204.200 72.935 204.245 ;
        RECT 72.170 204.060 72.935 204.200 ;
        RECT 72.170 204.000 72.490 204.060 ;
        RECT 72.645 204.015 72.935 204.060 ;
        RECT 78.165 204.015 78.455 204.245 ;
        RECT 79.530 204.000 79.850 204.260 ;
        RECT 85.510 204.000 85.830 204.260 ;
        RECT 18.280 203.380 93.120 203.860 ;
        RECT 44.585 203.180 44.875 203.225 ;
        RECT 52.850 203.180 53.170 203.240 ;
        RECT 56.085 203.180 56.375 203.225 ;
        RECT 56.530 203.180 56.850 203.240 ;
        RECT 60.210 203.180 60.530 203.240 ;
        RECT 44.585 203.040 54.920 203.180 ;
        RECT 44.585 202.995 44.875 203.040 ;
        RECT 52.850 202.980 53.170 203.040 ;
        RECT 41.810 202.840 42.130 202.900 ;
        RECT 40.980 202.700 54.460 202.840 ;
        RECT 39.625 202.500 39.915 202.545 ;
        RECT 40.430 202.500 40.750 202.560 ;
        RECT 40.980 202.545 41.120 202.700 ;
        RECT 41.810 202.640 42.130 202.700 ;
        RECT 39.625 202.360 40.750 202.500 ;
        RECT 39.625 202.315 39.915 202.360 ;
        RECT 40.430 202.300 40.750 202.360 ;
        RECT 40.905 202.315 41.195 202.545 ;
        RECT 41.350 202.500 41.670 202.560 ;
        RECT 50.090 202.545 50.410 202.560 ;
        RECT 51.560 202.545 51.700 202.700 ;
        RECT 42.745 202.500 43.035 202.545 ;
        RECT 41.350 202.360 43.035 202.500 ;
        RECT 41.350 202.300 41.670 202.360 ;
        RECT 42.745 202.315 43.035 202.360 ;
        RECT 50.090 202.315 50.440 202.545 ;
        RECT 51.485 202.315 51.775 202.545 ;
        RECT 36.315 202.160 36.605 202.205 ;
        RECT 38.835 202.160 39.125 202.205 ;
        RECT 40.025 202.160 40.315 202.205 ;
        RECT 36.315 202.020 40.315 202.160 ;
        RECT 36.315 201.975 36.605 202.020 ;
        RECT 38.835 201.975 39.125 202.020 ;
        RECT 40.025 201.975 40.315 202.020 ;
        RECT 36.750 201.820 37.040 201.865 ;
        RECT 38.320 201.820 38.610 201.865 ;
        RECT 40.420 201.820 40.710 201.865 ;
        RECT 36.750 201.680 40.710 201.820 ;
        RECT 36.750 201.635 37.040 201.680 ;
        RECT 38.320 201.635 38.610 201.680 ;
        RECT 40.420 201.635 40.710 201.680 ;
        RECT 34.005 201.480 34.295 201.525 ;
        RECT 39.510 201.480 39.830 201.540 ;
        RECT 34.005 201.340 39.830 201.480 ;
        RECT 34.005 201.295 34.295 201.340 ;
        RECT 39.510 201.280 39.830 201.340 ;
        RECT 41.350 201.480 41.670 201.540 ;
        RECT 41.825 201.480 42.115 201.525 ;
        RECT 41.350 201.340 42.115 201.480 ;
        RECT 41.350 201.280 41.670 201.340 ;
        RECT 41.825 201.295 42.115 201.340 ;
        RECT 42.270 201.480 42.590 201.540 ;
        RECT 42.820 201.480 42.960 202.315 ;
        RECT 50.090 202.300 50.410 202.315 ;
        RECT 53.310 202.300 53.630 202.560 ;
        RECT 46.895 202.160 47.185 202.205 ;
        RECT 49.415 202.160 49.705 202.205 ;
        RECT 50.605 202.160 50.895 202.205 ;
        RECT 46.895 202.020 50.895 202.160 ;
        RECT 46.895 201.975 47.185 202.020 ;
        RECT 49.415 201.975 49.705 202.020 ;
        RECT 50.605 201.975 50.895 202.020 ;
        RECT 47.330 201.820 47.620 201.865 ;
        RECT 48.900 201.820 49.190 201.865 ;
        RECT 51.000 201.820 51.290 201.865 ;
        RECT 53.400 201.820 53.540 202.300 ;
        RECT 54.320 202.160 54.460 202.700 ;
        RECT 54.780 202.545 54.920 203.040 ;
        RECT 56.085 203.040 60.530 203.180 ;
        RECT 56.085 202.995 56.375 203.040 ;
        RECT 56.530 202.980 56.850 203.040 ;
        RECT 60.210 202.980 60.530 203.040 ;
        RECT 85.510 202.980 85.830 203.240 ;
        RECT 79.085 202.840 79.375 202.885 ;
        RECT 79.530 202.840 79.850 202.900 ;
        RECT 63.060 202.700 77.460 202.840 ;
        RECT 61.590 202.545 61.910 202.560 ;
        RECT 54.705 202.315 54.995 202.545 ;
        RECT 61.590 202.315 61.940 202.545 ;
        RECT 61.590 202.300 61.910 202.315 ;
        RECT 63.060 202.220 63.200 202.700 ;
        RECT 77.320 202.545 77.460 202.700 ;
        RECT 79.085 202.700 79.850 202.840 ;
        RECT 79.085 202.655 79.375 202.700 ;
        RECT 79.530 202.640 79.850 202.700 ;
        RECT 81.365 202.840 82.015 202.885 ;
        RECT 84.965 202.840 85.255 202.885 ;
        RECT 81.365 202.700 85.255 202.840 ;
        RECT 81.365 202.655 82.015 202.700 ;
        RECT 84.665 202.655 85.255 202.700 ;
        RECT 69.425 202.500 69.715 202.545 ;
        RECT 75.910 202.500 76.200 202.545 ;
        RECT 69.425 202.360 76.200 202.500 ;
        RECT 69.425 202.315 69.715 202.360 ;
        RECT 75.910 202.315 76.200 202.360 ;
        RECT 77.245 202.500 77.535 202.545 ;
        RECT 77.690 202.500 78.010 202.560 ;
        RECT 77.245 202.360 78.010 202.500 ;
        RECT 77.245 202.315 77.535 202.360 ;
        RECT 77.690 202.300 78.010 202.360 ;
        RECT 78.170 202.500 78.460 202.545 ;
        RECT 80.005 202.500 80.295 202.545 ;
        RECT 83.585 202.500 83.875 202.545 ;
        RECT 78.170 202.360 83.875 202.500 ;
        RECT 78.170 202.315 78.460 202.360 ;
        RECT 80.005 202.315 80.295 202.360 ;
        RECT 83.585 202.315 83.875 202.360 ;
        RECT 84.665 202.340 84.955 202.655 ;
        RECT 85.600 202.500 85.740 202.980 ;
        RECT 87.365 202.500 87.655 202.545 ;
        RECT 85.600 202.360 87.655 202.500 ;
        RECT 57.910 202.160 58.230 202.220 ;
        RECT 54.320 202.020 58.230 202.160 ;
        RECT 57.910 201.960 58.230 202.020 ;
        RECT 58.395 202.160 58.685 202.205 ;
        RECT 60.915 202.160 61.205 202.205 ;
        RECT 62.105 202.160 62.395 202.205 ;
        RECT 58.395 202.020 62.395 202.160 ;
        RECT 58.395 201.975 58.685 202.020 ;
        RECT 60.915 201.975 61.205 202.020 ;
        RECT 62.105 201.975 62.395 202.020 ;
        RECT 62.970 201.960 63.290 202.220 ;
        RECT 66.190 201.960 66.510 202.220 ;
        RECT 66.650 202.160 66.970 202.220 ;
        RECT 68.045 202.160 68.335 202.205 ;
        RECT 66.650 202.020 68.335 202.160 ;
        RECT 66.650 201.960 66.970 202.020 ;
        RECT 68.045 201.975 68.335 202.020 ;
        RECT 68.505 202.160 68.795 202.205 ;
        RECT 72.170 202.160 72.490 202.220 ;
        RECT 68.505 202.020 72.490 202.160 ;
        RECT 68.505 201.975 68.795 202.020 ;
        RECT 72.170 201.960 72.490 202.020 ;
        RECT 72.655 202.160 72.945 202.205 ;
        RECT 75.175 202.160 75.465 202.205 ;
        RECT 76.365 202.160 76.655 202.205 ;
        RECT 72.655 202.020 76.655 202.160 ;
        RECT 84.680 202.160 84.820 202.340 ;
        RECT 87.365 202.315 87.655 202.360 ;
        RECT 87.825 202.160 88.115 202.205 ;
        RECT 84.680 202.020 88.115 202.160 ;
        RECT 72.655 201.975 72.945 202.020 ;
        RECT 75.175 201.975 75.465 202.020 ;
        RECT 76.365 201.975 76.655 202.020 ;
        RECT 87.825 201.975 88.115 202.020 ;
        RECT 47.330 201.680 51.290 201.820 ;
        RECT 47.330 201.635 47.620 201.680 ;
        RECT 48.900 201.635 49.190 201.680 ;
        RECT 51.000 201.635 51.290 201.680 ;
        RECT 51.560 201.680 53.540 201.820 ;
        RECT 58.830 201.820 59.120 201.865 ;
        RECT 60.400 201.820 60.690 201.865 ;
        RECT 62.500 201.820 62.790 201.865 ;
        RECT 58.830 201.680 62.790 201.820 ;
        RECT 51.560 201.480 51.700 201.680 ;
        RECT 58.830 201.635 59.120 201.680 ;
        RECT 60.400 201.635 60.690 201.680 ;
        RECT 62.500 201.635 62.790 201.680 ;
        RECT 73.090 201.820 73.380 201.865 ;
        RECT 74.660 201.820 74.950 201.865 ;
        RECT 76.760 201.820 77.050 201.865 ;
        RECT 73.090 201.680 77.050 201.820 ;
        RECT 73.090 201.635 73.380 201.680 ;
        RECT 74.660 201.635 74.950 201.680 ;
        RECT 76.760 201.635 77.050 201.680 ;
        RECT 78.575 201.820 78.865 201.865 ;
        RECT 80.465 201.820 80.755 201.865 ;
        RECT 83.585 201.820 83.875 201.865 ;
        RECT 78.575 201.680 83.875 201.820 ;
        RECT 78.575 201.635 78.865 201.680 ;
        RECT 80.465 201.635 80.755 201.680 ;
        RECT 83.585 201.635 83.875 201.680 ;
        RECT 42.270 201.340 51.700 201.480 ;
        RECT 42.270 201.280 42.590 201.340 ;
        RECT 51.930 201.280 52.250 201.540 ;
        RECT 52.390 201.480 52.710 201.540 ;
        RECT 52.865 201.480 53.155 201.525 ;
        RECT 52.390 201.340 53.155 201.480 ;
        RECT 52.390 201.280 52.710 201.340 ;
        RECT 52.865 201.295 53.155 201.340 ;
        RECT 61.130 201.480 61.450 201.540 ;
        RECT 70.330 201.480 70.650 201.540 ;
        RECT 61.130 201.340 70.650 201.480 ;
        RECT 61.130 201.280 61.450 201.340 ;
        RECT 70.330 201.280 70.650 201.340 ;
        RECT 86.430 201.280 86.750 201.540 ;
        RECT 18.280 200.660 92.340 201.140 ;
        RECT 39.970 200.260 40.290 200.520 ;
        RECT 40.430 200.260 40.750 200.520 ;
        RECT 50.090 200.460 50.410 200.520 ;
        RECT 50.565 200.460 50.855 200.505 ;
        RECT 50.090 200.320 50.855 200.460 ;
        RECT 50.090 200.260 50.410 200.320 ;
        RECT 50.565 200.275 50.855 200.320 ;
        RECT 61.590 200.260 61.910 200.520 ;
        RECT 66.190 200.460 66.510 200.520 ;
        RECT 67.585 200.460 67.875 200.505 ;
        RECT 66.190 200.320 67.875 200.460 ;
        RECT 66.190 200.260 66.510 200.320 ;
        RECT 67.585 200.275 67.875 200.320 ;
        RECT 69.870 200.460 70.190 200.520 ;
        RECT 70.790 200.460 71.110 200.520 ;
        RECT 71.725 200.460 72.015 200.505 ;
        RECT 69.870 200.320 72.015 200.460 ;
        RECT 69.870 200.260 70.190 200.320 ;
        RECT 70.790 200.260 71.110 200.320 ;
        RECT 71.725 200.275 72.015 200.320 ;
        RECT 75.850 200.460 76.170 200.520 ;
        RECT 85.050 200.460 85.370 200.520 ;
        RECT 75.850 200.320 85.370 200.460 ;
        RECT 75.850 200.260 76.170 200.320 ;
        RECT 85.050 200.260 85.370 200.320 ;
        RECT 40.060 200.120 40.200 200.260 ;
        RECT 46.410 200.120 46.730 200.180 ;
        RECT 59.290 200.120 59.610 200.180 ;
        RECT 69.410 200.120 69.730 200.180 ;
        RECT 40.060 199.980 46.730 200.120 ;
        RECT 46.410 199.920 46.730 199.980 ;
        RECT 46.960 199.980 60.440 200.120 ;
        RECT 37.225 199.780 37.515 199.825 ;
        RECT 38.590 199.780 38.910 199.840 ;
        RECT 41.350 199.780 41.670 199.840 ;
        RECT 37.225 199.640 38.910 199.780 ;
        RECT 37.225 199.595 37.515 199.640 ;
        RECT 38.590 199.580 38.910 199.640 ;
        RECT 39.140 199.640 43.190 199.780 ;
        RECT 38.130 199.440 38.450 199.500 ;
        RECT 39.140 199.485 39.280 199.640 ;
        RECT 41.350 199.580 41.670 199.640 ;
        RECT 39.065 199.440 39.355 199.485 ;
        RECT 38.130 199.300 39.355 199.440 ;
        RECT 38.130 199.240 38.450 199.300 ;
        RECT 39.065 199.255 39.355 199.300 ;
        RECT 39.525 199.255 39.815 199.485 ;
        RECT 43.050 199.440 43.190 199.640 ;
        RECT 46.960 199.440 47.100 199.980 ;
        RECT 59.290 199.920 59.610 199.980 ;
        RECT 47.345 199.780 47.635 199.825 ;
        RECT 51.930 199.780 52.250 199.840 ;
        RECT 47.345 199.640 52.250 199.780 ;
        RECT 47.345 199.595 47.635 199.640 ;
        RECT 51.930 199.580 52.250 199.640 ;
        RECT 57.450 199.780 57.770 199.840 ;
        RECT 58.385 199.780 58.675 199.825 ;
        RECT 57.450 199.640 58.675 199.780 ;
        RECT 57.450 199.580 57.770 199.640 ;
        RECT 58.385 199.595 58.675 199.640 ;
        RECT 49.185 199.440 49.475 199.485 ;
        RECT 43.050 199.300 49.475 199.440 ;
        RECT 49.185 199.255 49.475 199.300 ;
        RECT 49.645 199.440 49.935 199.485 ;
        RECT 53.770 199.440 54.090 199.500 ;
        RECT 59.750 199.440 60.070 199.500 ;
        RECT 60.300 199.485 60.440 199.980 ;
        RECT 60.760 199.980 69.730 200.120 ;
        RECT 60.760 199.485 60.900 199.980 ;
        RECT 69.410 199.920 69.730 199.980 ;
        RECT 79.990 199.920 80.310 200.180 ;
        RECT 86.430 199.780 86.750 199.840 ;
        RECT 73.180 199.640 88.500 199.780 ;
        RECT 49.645 199.300 60.070 199.440 ;
        RECT 49.645 199.255 49.935 199.300 ;
        RECT 39.600 199.100 39.740 199.255 ;
        RECT 53.770 199.240 54.090 199.300 ;
        RECT 59.750 199.240 60.070 199.300 ;
        RECT 60.225 199.255 60.515 199.485 ;
        RECT 60.685 199.255 60.975 199.485 ;
        RECT 66.650 199.440 66.970 199.500 ;
        RECT 70.330 199.485 70.650 199.500 ;
        RECT 68.505 199.440 68.795 199.485 ;
        RECT 70.315 199.440 70.650 199.485 ;
        RECT 66.650 199.300 68.795 199.440 ;
        RECT 70.135 199.300 70.650 199.440 ;
        RECT 66.650 199.240 66.970 199.300 ;
        RECT 68.505 199.255 68.795 199.300 ;
        RECT 70.315 199.255 70.650 199.300 ;
        RECT 70.330 199.240 70.650 199.255 ;
        RECT 42.730 199.100 43.050 199.160 ;
        RECT 72.630 199.100 72.950 199.160 ;
        RECT 73.180 199.145 73.320 199.640 ;
        RECT 86.430 199.580 86.750 199.640 ;
        RECT 74.930 199.240 75.250 199.500 ;
        RECT 75.850 199.240 76.170 199.500 ;
        RECT 76.310 199.240 76.630 199.500 ;
        RECT 77.230 199.240 77.550 199.500 ;
        RECT 78.610 199.240 78.930 199.500 ;
        RECT 87.810 199.240 88.130 199.500 ;
        RECT 88.360 199.485 88.500 199.640 ;
        RECT 88.285 199.255 88.575 199.485 ;
        RECT 91.030 199.240 91.350 199.500 ;
        RECT 39.600 198.960 72.950 199.100 ;
        RECT 42.730 198.900 43.050 198.960 ;
        RECT 72.630 198.900 72.950 198.960 ;
        RECT 73.105 198.915 73.395 199.145 ;
        RECT 75.405 199.100 75.695 199.145 ;
        RECT 79.085 199.100 79.375 199.145 ;
        RECT 75.405 198.960 79.375 199.100 ;
        RECT 75.405 198.915 75.695 198.960 ;
        RECT 79.085 198.915 79.375 198.960 ;
        RECT 80.005 199.100 80.295 199.145 ;
        RECT 80.450 199.100 80.770 199.160 ;
        RECT 80.005 198.960 80.770 199.100 ;
        RECT 87.900 199.100 88.040 199.240 ;
        RECT 91.120 199.100 91.260 199.240 ;
        RECT 87.900 198.960 91.260 199.100 ;
        RECT 80.005 198.915 80.295 198.960 ;
        RECT 46.410 198.760 46.730 198.820 ;
        RECT 52.390 198.760 52.710 198.820 ;
        RECT 53.770 198.760 54.090 198.820 ;
        RECT 73.180 198.760 73.320 198.915 ;
        RECT 80.450 198.900 80.770 198.960 ;
        RECT 46.410 198.620 73.320 198.760 ;
        RECT 46.410 198.560 46.730 198.620 ;
        RECT 52.390 198.560 52.710 198.620 ;
        RECT 53.770 198.560 54.090 198.620 ;
        RECT 76.770 198.560 77.090 198.820 ;
        RECT 79.530 198.760 79.850 198.820 ;
        RECT 84.605 198.760 84.895 198.805 ;
        RECT 79.530 198.620 84.895 198.760 ;
        RECT 79.530 198.560 79.850 198.620 ;
        RECT 84.605 198.575 84.895 198.620 ;
        RECT 88.730 198.560 89.050 198.820 ;
        RECT 18.280 197.940 93.120 198.420 ;
        RECT 74.930 197.740 75.250 197.800 ;
        RECT 76.325 197.740 76.615 197.785 ;
        RECT 74.930 197.600 76.615 197.740 ;
        RECT 74.930 197.540 75.250 197.600 ;
        RECT 76.325 197.555 76.615 197.600 ;
        RECT 76.770 197.540 77.090 197.800 ;
        RECT 77.690 197.540 78.010 197.800 ;
        RECT 78.610 197.740 78.930 197.800 ;
        RECT 79.085 197.740 79.375 197.785 ;
        RECT 78.610 197.600 79.375 197.740 ;
        RECT 78.610 197.540 78.930 197.600 ;
        RECT 79.085 197.555 79.375 197.600 ;
        RECT 90.125 197.740 90.415 197.785 ;
        RECT 91.030 197.740 91.350 197.800 ;
        RECT 90.125 197.600 91.350 197.740 ;
        RECT 90.125 197.555 90.415 197.600 ;
        RECT 91.030 197.540 91.350 197.600 ;
        RECT 75.850 197.400 76.170 197.460 ;
        RECT 56.620 197.260 76.170 197.400 ;
        RECT 37.225 197.060 37.515 197.105 ;
        RECT 38.130 197.060 38.450 197.120 ;
        RECT 45.965 197.060 46.255 197.105 ;
        RECT 56.620 197.060 56.760 197.260 ;
        RECT 75.850 197.200 76.170 197.260 ;
        RECT 37.225 196.920 38.450 197.060 ;
        RECT 37.225 196.875 37.515 196.920 ;
        RECT 38.130 196.860 38.450 196.920 ;
        RECT 43.050 196.920 46.255 197.060 ;
        RECT 34.925 196.720 35.215 196.765 ;
        RECT 36.290 196.720 36.610 196.780 ;
        RECT 34.925 196.580 36.610 196.720 ;
        RECT 34.925 196.535 35.215 196.580 ;
        RECT 36.290 196.520 36.610 196.580 ;
        RECT 36.765 196.535 37.055 196.765 ;
        RECT 38.220 196.720 38.360 196.860 ;
        RECT 43.050 196.720 43.190 196.920 ;
        RECT 45.965 196.875 46.255 196.920 ;
        RECT 47.420 196.920 56.760 197.060 ;
        RECT 57.105 197.060 57.395 197.105 ;
        RECT 58.830 197.060 59.150 197.120 ;
        RECT 62.050 197.105 62.370 197.120 ;
        RECT 57.105 196.920 59.150 197.060 ;
        RECT 38.220 196.580 43.190 196.720 ;
        RECT 45.505 196.680 45.795 196.765 ;
        RECT 46.870 196.720 47.190 196.780 ;
        RECT 47.420 196.720 47.560 196.920 ;
        RECT 57.105 196.875 57.395 196.920 ;
        RECT 58.830 196.860 59.150 196.920 ;
        RECT 62.020 196.875 62.370 197.105 ;
        RECT 73.795 197.060 74.085 197.105 ;
        RECT 62.050 196.860 62.370 196.875 ;
        RECT 65.820 196.920 74.085 197.060 ;
        RECT 46.500 196.680 47.560 196.720 ;
        RECT 45.505 196.580 47.560 196.680 ;
        RECT 45.505 196.540 46.640 196.580 ;
        RECT 45.505 196.535 45.795 196.540 ;
        RECT 36.840 196.380 36.980 196.535 ;
        RECT 46.870 196.520 47.190 196.580 ;
        RECT 47.790 196.520 48.110 196.780 ;
        RECT 53.795 196.720 54.085 196.765 ;
        RECT 56.315 196.720 56.605 196.765 ;
        RECT 57.505 196.720 57.795 196.765 ;
        RECT 53.795 196.580 57.795 196.720 ;
        RECT 53.795 196.535 54.085 196.580 ;
        RECT 56.315 196.535 56.605 196.580 ;
        RECT 57.505 196.535 57.795 196.580 ;
        RECT 58.370 196.720 58.690 196.780 ;
        RECT 60.685 196.720 60.975 196.765 ;
        RECT 58.370 196.580 60.975 196.720 ;
        RECT 58.370 196.520 58.690 196.580 ;
        RECT 60.685 196.535 60.975 196.580 ;
        RECT 61.565 196.720 61.855 196.765 ;
        RECT 62.755 196.720 63.045 196.765 ;
        RECT 65.275 196.720 65.565 196.765 ;
        RECT 61.565 196.580 65.565 196.720 ;
        RECT 61.565 196.535 61.855 196.580 ;
        RECT 62.755 196.535 63.045 196.580 ;
        RECT 65.275 196.535 65.565 196.580 ;
        RECT 37.210 196.380 37.530 196.440 ;
        RECT 54.230 196.380 54.520 196.425 ;
        RECT 55.800 196.380 56.090 196.425 ;
        RECT 57.900 196.380 58.190 196.425 ;
        RECT 36.840 196.240 54.000 196.380 ;
        RECT 37.210 196.180 37.530 196.240 ;
        RECT 38.130 195.840 38.450 196.100 ;
        RECT 44.570 195.840 44.890 196.100 ;
        RECT 51.485 196.040 51.775 196.085 ;
        RECT 52.390 196.040 52.710 196.100 ;
        RECT 51.485 195.900 52.710 196.040 ;
        RECT 53.860 196.040 54.000 196.240 ;
        RECT 54.230 196.240 58.190 196.380 ;
        RECT 54.230 196.195 54.520 196.240 ;
        RECT 55.800 196.195 56.090 196.240 ;
        RECT 57.900 196.195 58.190 196.240 ;
        RECT 61.170 196.380 61.460 196.425 ;
        RECT 63.270 196.380 63.560 196.425 ;
        RECT 64.840 196.380 65.130 196.425 ;
        RECT 61.170 196.240 65.130 196.380 ;
        RECT 61.170 196.195 61.460 196.240 ;
        RECT 63.270 196.195 63.560 196.240 ;
        RECT 64.840 196.195 65.130 196.240 ;
        RECT 65.820 196.040 65.960 196.920 ;
        RECT 73.795 196.875 74.085 196.920 ;
        RECT 74.470 196.860 74.790 197.120 ;
        RECT 74.930 196.860 75.250 197.120 ;
        RECT 75.405 197.060 75.695 197.105 ;
        RECT 76.860 197.060 77.000 197.540 ;
        RECT 77.780 197.400 77.920 197.540 ;
        RECT 81.830 197.400 82.150 197.460 ;
        RECT 83.230 197.400 83.520 197.445 ;
        RECT 84.630 197.400 84.920 197.445 ;
        RECT 86.470 197.400 86.760 197.445 ;
        RECT 77.780 197.260 82.520 197.400 ;
        RECT 81.830 197.200 82.150 197.260 ;
        RECT 75.405 196.920 77.000 197.060 ;
        RECT 77.230 197.060 77.550 197.120 ;
        RECT 77.705 197.060 77.995 197.105 ;
        RECT 77.230 196.920 77.995 197.060 ;
        RECT 75.405 196.875 75.695 196.920 ;
        RECT 77.230 196.860 77.550 196.920 ;
        RECT 77.705 196.875 77.995 196.920 ;
        RECT 79.530 196.860 79.850 197.120 ;
        RECT 79.990 196.860 80.310 197.120 ;
        RECT 82.380 197.105 82.520 197.260 ;
        RECT 83.230 197.260 86.760 197.400 ;
        RECT 83.230 197.215 83.520 197.260 ;
        RECT 84.630 197.215 84.920 197.260 ;
        RECT 86.470 197.215 86.760 197.260 ;
        RECT 82.305 196.875 82.595 197.105 ;
        RECT 71.710 196.720 72.030 196.780 ;
        RECT 73.105 196.720 73.395 196.765 ;
        RECT 71.710 196.580 73.395 196.720 ;
        RECT 71.710 196.520 72.030 196.580 ;
        RECT 73.105 196.535 73.395 196.580 ;
        RECT 79.085 196.720 79.375 196.765 ;
        RECT 79.620 196.720 79.760 196.860 ;
        RECT 79.085 196.580 79.760 196.720 ;
        RECT 80.080 196.720 80.220 196.860 ;
        RECT 83.685 196.720 83.975 196.765 ;
        RECT 80.080 196.580 83.975 196.720 ;
        RECT 79.085 196.535 79.375 196.580 ;
        RECT 83.685 196.535 83.975 196.580 ;
        RECT 82.770 196.380 83.060 196.425 ;
        RECT 85.090 196.380 85.380 196.425 ;
        RECT 86.470 196.380 86.760 196.425 ;
        RECT 82.770 196.240 86.760 196.380 ;
        RECT 82.770 196.195 83.060 196.240 ;
        RECT 85.090 196.195 85.380 196.240 ;
        RECT 86.470 196.195 86.760 196.240 ;
        RECT 53.860 195.900 65.960 196.040 ;
        RECT 51.485 195.855 51.775 195.900 ;
        RECT 52.390 195.840 52.710 195.900 ;
        RECT 67.570 195.840 67.890 196.100 ;
        RECT 78.150 195.840 78.470 196.100 ;
        RECT 18.280 195.220 92.340 195.700 ;
        RECT 47.790 195.020 48.110 195.080 ;
        RECT 49.185 195.020 49.475 195.065 ;
        RECT 47.790 194.880 49.475 195.020 ;
        RECT 47.790 194.820 48.110 194.880 ;
        RECT 49.185 194.835 49.475 194.880 ;
        RECT 51.025 195.020 51.315 195.065 ;
        RECT 51.930 195.020 52.250 195.080 ;
        RECT 51.025 194.880 52.250 195.020 ;
        RECT 51.025 194.835 51.315 194.880 ;
        RECT 51.930 194.820 52.250 194.880 ;
        RECT 53.310 194.820 53.630 195.080 ;
        RECT 53.770 195.020 54.090 195.080 ;
        RECT 54.245 195.020 54.535 195.065 ;
        RECT 53.770 194.880 54.535 195.020 ;
        RECT 53.770 194.820 54.090 194.880 ;
        RECT 54.245 194.835 54.535 194.880 ;
        RECT 58.830 195.020 59.150 195.080 ;
        RECT 60.685 195.020 60.975 195.065 ;
        RECT 58.830 194.880 60.975 195.020 ;
        RECT 58.830 194.820 59.150 194.880 ;
        RECT 60.685 194.835 60.975 194.880 ;
        RECT 62.050 195.020 62.370 195.080 ;
        RECT 65.285 195.020 65.575 195.065 ;
        RECT 62.050 194.880 65.575 195.020 ;
        RECT 62.050 194.820 62.370 194.880 ;
        RECT 65.285 194.835 65.575 194.880 ;
        RECT 68.950 195.020 69.270 195.080 ;
        RECT 69.885 195.020 70.175 195.065 ;
        RECT 70.790 195.020 71.110 195.080 ;
        RECT 68.950 194.880 71.110 195.020 ;
        RECT 68.950 194.820 69.270 194.880 ;
        RECT 69.885 194.835 70.175 194.880 ;
        RECT 70.790 194.820 71.110 194.880 ;
        RECT 74.470 195.020 74.790 195.080 ;
        RECT 74.470 194.880 80.220 195.020 ;
        RECT 74.470 194.820 74.790 194.880 ;
        RECT 34.450 194.680 34.740 194.725 ;
        RECT 36.020 194.680 36.310 194.725 ;
        RECT 38.120 194.680 38.410 194.725 ;
        RECT 34.450 194.540 38.410 194.680 ;
        RECT 34.450 194.495 34.740 194.540 ;
        RECT 36.020 194.495 36.310 194.540 ;
        RECT 38.120 194.495 38.410 194.540 ;
        RECT 42.310 194.680 42.600 194.725 ;
        RECT 44.410 194.680 44.700 194.725 ;
        RECT 45.980 194.680 46.270 194.725 ;
        RECT 53.400 194.680 53.540 194.820 ;
        RECT 69.040 194.680 69.180 194.820 ;
        RECT 42.310 194.540 46.270 194.680 ;
        RECT 42.310 194.495 42.600 194.540 ;
        RECT 44.410 194.495 44.700 194.540 ;
        RECT 45.980 194.495 46.270 194.540 ;
        RECT 50.640 194.540 55.380 194.680 ;
        RECT 34.015 194.340 34.305 194.385 ;
        RECT 36.535 194.340 36.825 194.385 ;
        RECT 37.725 194.340 38.015 194.385 ;
        RECT 34.015 194.200 38.015 194.340 ;
        RECT 34.015 194.155 34.305 194.200 ;
        RECT 36.535 194.155 36.825 194.200 ;
        RECT 37.725 194.155 38.015 194.200 ;
        RECT 38.605 194.340 38.895 194.385 ;
        RECT 41.810 194.340 42.130 194.400 ;
        RECT 50.640 194.385 50.780 194.540 ;
        RECT 38.605 194.200 42.130 194.340 ;
        RECT 38.605 194.155 38.895 194.200 ;
        RECT 41.810 194.140 42.130 194.200 ;
        RECT 42.705 194.340 42.995 194.385 ;
        RECT 43.895 194.340 44.185 194.385 ;
        RECT 46.415 194.340 46.705 194.385 ;
        RECT 42.705 194.200 46.705 194.340 ;
        RECT 42.705 194.155 42.995 194.200 ;
        RECT 43.895 194.155 44.185 194.200 ;
        RECT 46.415 194.155 46.705 194.200 ;
        RECT 50.565 194.155 50.855 194.385 ;
        RECT 52.390 194.340 52.710 194.400 ;
        RECT 55.240 194.385 55.380 194.540 ;
        RECT 58.920 194.540 69.180 194.680 ;
        RECT 51.100 194.200 52.160 194.340 ;
        RECT 37.325 194.000 37.615 194.045 ;
        RECT 38.130 194.000 38.450 194.060 ;
        RECT 37.325 193.860 38.450 194.000 ;
        RECT 37.325 193.815 37.615 193.860 ;
        RECT 38.130 193.800 38.450 193.860 ;
        RECT 43.160 194.000 43.450 194.045 ;
        RECT 44.570 194.000 44.890 194.060 ;
        RECT 51.100 194.045 51.240 194.200 ;
        RECT 43.160 193.860 44.890 194.000 ;
        RECT 43.160 193.815 43.450 193.860 ;
        RECT 44.570 193.800 44.890 193.860 ;
        RECT 50.995 193.815 51.285 194.045 ;
        RECT 51.485 193.815 51.775 194.045 ;
        RECT 52.020 194.000 52.160 194.200 ;
        RECT 52.390 194.200 54.000 194.340 ;
        RECT 52.390 194.140 52.710 194.200 ;
        RECT 53.860 194.045 54.000 194.200 ;
        RECT 55.165 194.155 55.455 194.385 ;
        RECT 52.020 193.860 53.540 194.000 ;
        RECT 51.560 193.660 51.700 193.815 ;
        RECT 50.180 193.520 51.700 193.660 ;
        RECT 53.400 193.660 53.540 193.860 ;
        RECT 53.785 193.815 54.075 194.045 ;
        RECT 58.920 193.660 59.060 194.540 ;
        RECT 59.290 194.340 59.610 194.400 ;
        RECT 66.650 194.340 66.970 194.400 ;
        RECT 59.290 194.200 66.970 194.340 ;
        RECT 59.290 194.140 59.610 194.200 ;
        RECT 66.650 194.140 66.970 194.200 ;
        RECT 67.660 194.200 70.790 194.340 ;
        RECT 59.765 194.000 60.055 194.045 ;
        RECT 60.670 194.000 60.990 194.060 ;
        RECT 59.765 193.860 60.990 194.000 ;
        RECT 59.765 193.815 60.055 193.860 ;
        RECT 60.670 193.800 60.990 193.860 ;
        RECT 66.205 193.815 66.495 194.045 ;
        RECT 53.400 193.520 59.060 193.660 ;
        RECT 50.180 193.380 50.320 193.520 ;
        RECT 31.690 193.120 32.010 193.380 ;
        RECT 48.725 193.320 49.015 193.365 ;
        RECT 50.090 193.320 50.410 193.380 ;
        RECT 48.725 193.180 50.410 193.320 ;
        RECT 48.725 193.135 49.015 193.180 ;
        RECT 50.090 193.120 50.410 193.180 ;
        RECT 51.930 193.120 52.250 193.380 ;
        RECT 56.545 193.320 56.835 193.365 ;
        RECT 57.465 193.320 57.755 193.365 ;
        RECT 56.545 193.180 57.755 193.320 ;
        RECT 66.280 193.320 66.420 193.815 ;
        RECT 66.740 193.660 66.880 194.140 ;
        RECT 67.660 194.060 67.800 194.200 ;
        RECT 67.570 193.800 67.890 194.060 ;
        RECT 69.885 193.815 70.175 194.045 ;
        RECT 70.650 194.000 70.790 194.200 ;
        RECT 71.725 194.000 72.015 194.045 ;
        RECT 70.650 193.860 72.015 194.000 ;
        RECT 71.725 193.815 72.015 193.860 ;
        RECT 72.185 193.815 72.475 194.045 ;
        RECT 72.630 194.000 72.950 194.060 ;
        RECT 74.560 194.045 74.700 194.820 ;
        RECT 80.080 194.740 80.220 194.880 ;
        RECT 78.610 194.680 78.930 194.740 ;
        RECT 75.480 194.540 78.930 194.680 ;
        RECT 74.930 194.340 75.250 194.400 ;
        RECT 75.480 194.340 75.620 194.540 ;
        RECT 78.610 194.480 78.930 194.540 ;
        RECT 79.085 194.495 79.375 194.725 ;
        RECT 74.930 194.200 75.620 194.340 ;
        RECT 74.930 194.140 75.250 194.200 ;
        RECT 75.480 194.045 75.620 194.200 ;
        RECT 77.230 194.140 77.550 194.400 ;
        RECT 79.160 194.340 79.300 194.495 ;
        RECT 79.990 194.480 80.310 194.740 ;
        RECT 79.160 194.200 85.740 194.340 ;
        RECT 73.105 194.000 73.395 194.045 ;
        RECT 72.630 193.860 73.395 194.000 ;
        RECT 69.960 193.660 70.100 193.815 ;
        RECT 66.740 193.520 70.100 193.660 ;
        RECT 68.030 193.320 68.350 193.380 ;
        RECT 66.280 193.180 68.350 193.320 ;
        RECT 56.545 193.135 56.835 193.180 ;
        RECT 57.465 193.135 57.755 193.180 ;
        RECT 68.030 193.120 68.350 193.180 ;
        RECT 68.505 193.320 68.795 193.365 ;
        RECT 68.965 193.320 69.255 193.365 ;
        RECT 68.505 193.180 69.255 193.320 ;
        RECT 68.505 193.135 68.795 193.180 ;
        RECT 68.965 193.135 69.255 193.180 ;
        RECT 71.710 193.320 72.030 193.380 ;
        RECT 72.260 193.320 72.400 193.815 ;
        RECT 72.630 193.800 72.950 193.860 ;
        RECT 73.105 193.815 73.395 193.860 ;
        RECT 74.485 193.815 74.775 194.045 ;
        RECT 75.405 193.815 75.695 194.045 ;
        RECT 75.865 193.815 76.155 194.045 ;
        RECT 76.325 194.000 76.615 194.045 ;
        RECT 77.320 194.000 77.460 194.140 ;
        RECT 76.325 193.860 77.460 194.000 ;
        RECT 76.325 193.815 76.615 193.860 ;
        RECT 77.705 193.815 77.995 194.045 ;
        RECT 78.165 194.000 78.455 194.045 ;
        RECT 81.385 194.000 81.675 194.045 ;
        RECT 78.165 193.860 81.675 194.000 ;
        RECT 78.165 193.815 78.455 193.860 ;
        RECT 81.385 193.815 81.675 193.860 ;
        RECT 84.605 193.815 84.895 194.045 ;
        RECT 74.025 193.660 74.315 193.705 ;
        RECT 75.940 193.660 76.080 193.815 ;
        RECT 74.025 193.520 76.080 193.660 ;
        RECT 76.770 193.660 77.090 193.720 ;
        RECT 77.245 193.660 77.535 193.705 ;
        RECT 76.770 193.520 77.535 193.660 ;
        RECT 77.780 193.660 77.920 193.815 ;
        RECT 78.610 193.660 78.930 193.720 ;
        RECT 79.545 193.660 79.835 193.705 ;
        RECT 77.780 193.520 78.380 193.660 ;
        RECT 74.025 193.475 74.315 193.520 ;
        RECT 76.770 193.460 77.090 193.520 ;
        RECT 77.245 193.475 77.535 193.520 ;
        RECT 71.710 193.180 72.400 193.320 ;
        RECT 74.945 193.320 75.235 193.365 ;
        RECT 75.390 193.320 75.710 193.380 ;
        RECT 78.240 193.320 78.380 193.520 ;
        RECT 78.610 193.520 79.835 193.660 ;
        RECT 78.610 193.460 78.930 193.520 ;
        RECT 79.545 193.475 79.835 193.520 ;
        RECT 79.990 193.660 80.310 193.720 ;
        RECT 80.465 193.660 80.755 193.705 ;
        RECT 84.680 193.660 84.820 193.815 ;
        RECT 85.050 193.800 85.370 194.060 ;
        RECT 85.600 194.045 85.740 194.200 ;
        RECT 85.525 193.815 85.815 194.045 ;
        RECT 86.430 194.000 86.750 194.060 ;
        RECT 88.730 194.000 89.050 194.060 ;
        RECT 86.430 193.860 89.050 194.000 ;
        RECT 86.430 193.800 86.750 193.860 ;
        RECT 88.730 193.800 89.050 193.860 ;
        RECT 91.030 193.800 91.350 194.060 ;
        RECT 91.120 193.660 91.260 193.800 ;
        RECT 79.990 193.520 91.260 193.660 ;
        RECT 79.990 193.460 80.310 193.520 ;
        RECT 80.465 193.475 80.755 193.520 ;
        RECT 74.945 193.180 78.380 193.320 ;
        RECT 83.225 193.320 83.515 193.365 ;
        RECT 83.670 193.320 83.990 193.380 ;
        RECT 83.225 193.180 83.990 193.320 ;
        RECT 71.710 193.120 72.030 193.180 ;
        RECT 74.945 193.135 75.235 193.180 ;
        RECT 75.390 193.120 75.710 193.180 ;
        RECT 83.225 193.135 83.515 193.180 ;
        RECT 83.670 193.120 83.990 193.180 ;
        RECT 18.280 192.500 93.120 192.980 ;
        RECT 36.765 192.300 37.055 192.345 ;
        RECT 37.670 192.300 37.990 192.360 ;
        RECT 36.765 192.160 37.990 192.300 ;
        RECT 36.765 192.115 37.055 192.160 ;
        RECT 37.670 192.100 37.990 192.160 ;
        RECT 59.750 192.300 60.070 192.360 ;
        RECT 74.930 192.300 75.250 192.360 ;
        RECT 59.750 192.160 75.250 192.300 ;
        RECT 59.750 192.100 60.070 192.160 ;
        RECT 74.930 192.100 75.250 192.160 ;
        RECT 75.390 192.100 75.710 192.360 ;
        RECT 78.150 192.300 78.470 192.360 ;
        RECT 78.625 192.300 78.915 192.345 ;
        RECT 78.150 192.160 78.915 192.300 ;
        RECT 78.150 192.100 78.470 192.160 ;
        RECT 78.625 192.115 78.915 192.160 ;
        RECT 42.270 191.960 42.590 192.020 ;
        RECT 38.220 191.820 42.590 191.960 ;
        RECT 38.220 191.665 38.360 191.820 ;
        RECT 42.270 191.760 42.590 191.820 ;
        RECT 38.145 191.435 38.435 191.665 ;
        RECT 39.525 191.435 39.815 191.665 ;
        RECT 50.550 191.620 50.870 191.680 ;
        RECT 54.705 191.620 54.995 191.665 ;
        RECT 50.550 191.480 54.995 191.620 ;
        RECT 39.600 191.280 39.740 191.435 ;
        RECT 50.550 191.420 50.870 191.480 ;
        RECT 54.705 191.435 54.995 191.480 ;
        RECT 56.070 191.420 56.390 191.680 ;
        RECT 56.530 191.420 56.850 191.680 ;
        RECT 75.480 191.620 75.620 192.100 ;
        RECT 83.230 191.960 83.520 192.005 ;
        RECT 84.630 191.960 84.920 192.005 ;
        RECT 86.470 191.960 86.760 192.005 ;
        RECT 83.230 191.820 86.760 191.960 ;
        RECT 83.230 191.775 83.520 191.820 ;
        RECT 84.630 191.775 84.920 191.820 ;
        RECT 86.470 191.775 86.760 191.820 ;
        RECT 90.585 191.960 90.875 192.005 ;
        RECT 91.030 191.960 91.350 192.020 ;
        RECT 90.585 191.820 91.350 191.960 ;
        RECT 90.585 191.775 90.875 191.820 ;
        RECT 91.030 191.760 91.350 191.820 ;
        RECT 77.705 191.620 77.995 191.665 ;
        RECT 75.480 191.480 77.995 191.620 ;
        RECT 77.705 191.435 77.995 191.480 ;
        RECT 81.830 191.620 82.150 191.680 ;
        RECT 82.305 191.620 82.595 191.665 ;
        RECT 81.830 191.480 82.595 191.620 ;
        RECT 81.830 191.420 82.150 191.480 ;
        RECT 82.305 191.435 82.595 191.480 ;
        RECT 83.670 191.420 83.990 191.680 ;
        RECT 35.000 191.140 39.740 191.280 ;
        RECT 52.390 191.280 52.710 191.340 ;
        RECT 55.165 191.280 55.455 191.325 ;
        RECT 52.390 191.140 55.455 191.280 ;
        RECT 35.000 190.660 35.140 191.140 ;
        RECT 52.390 191.080 52.710 191.140 ;
        RECT 55.165 191.095 55.455 191.140 ;
        RECT 57.925 191.280 58.215 191.325 ;
        RECT 58.370 191.280 58.690 191.340 ;
        RECT 57.925 191.140 58.690 191.280 ;
        RECT 57.925 191.095 58.215 191.140 ;
        RECT 58.370 191.080 58.690 191.140 ;
        RECT 59.750 191.280 60.070 191.340 ;
        RECT 62.985 191.280 63.275 191.325 ;
        RECT 59.750 191.140 63.275 191.280 ;
        RECT 59.750 191.080 60.070 191.140 ;
        RECT 62.985 191.095 63.275 191.140 ;
        RECT 72.630 191.280 72.950 191.340 ;
        RECT 76.770 191.280 77.090 191.340 ;
        RECT 72.630 191.140 77.090 191.280 ;
        RECT 72.630 191.080 72.950 191.140 ;
        RECT 76.770 191.080 77.090 191.140 ;
        RECT 58.830 190.940 59.150 191.000 ;
        RECT 35.460 190.800 59.150 190.940 ;
        RECT 35.460 190.660 35.600 190.800 ;
        RECT 58.830 190.740 59.150 190.800 ;
        RECT 59.290 190.940 59.610 191.000 ;
        RECT 61.130 190.940 61.450 191.000 ;
        RECT 59.290 190.800 61.450 190.940 ;
        RECT 59.290 190.740 59.610 190.800 ;
        RECT 61.130 190.740 61.450 190.800 ;
        RECT 64.825 190.940 65.115 190.985 ;
        RECT 67.570 190.940 67.890 191.000 ;
        RECT 64.825 190.800 67.890 190.940 ;
        RECT 64.825 190.755 65.115 190.800 ;
        RECT 67.570 190.740 67.890 190.800 ;
        RECT 82.770 190.940 83.060 190.985 ;
        RECT 85.090 190.940 85.380 190.985 ;
        RECT 86.470 190.940 86.760 190.985 ;
        RECT 82.770 190.800 86.760 190.940 ;
        RECT 82.770 190.755 83.060 190.800 ;
        RECT 85.090 190.755 85.380 190.800 ;
        RECT 86.470 190.755 86.760 190.800 ;
        RECT 34.910 190.400 35.230 190.660 ;
        RECT 35.370 190.400 35.690 190.660 ;
        RECT 39.065 190.600 39.355 190.645 ;
        RECT 39.970 190.600 40.290 190.660 ;
        RECT 39.065 190.460 40.290 190.600 ;
        RECT 39.065 190.415 39.355 190.460 ;
        RECT 39.970 190.400 40.290 190.460 ;
        RECT 57.450 190.400 57.770 190.660 ;
        RECT 60.225 190.600 60.515 190.645 ;
        RECT 61.590 190.600 61.910 190.660 ;
        RECT 60.225 190.460 61.910 190.600 ;
        RECT 60.225 190.415 60.515 190.460 ;
        RECT 61.590 190.400 61.910 190.460 ;
        RECT 62.510 190.600 62.830 190.660 ;
        RECT 65.285 190.600 65.575 190.645 ;
        RECT 62.510 190.460 65.575 190.600 ;
        RECT 62.510 190.400 62.830 190.460 ;
        RECT 65.285 190.415 65.575 190.460 ;
        RECT 18.280 189.780 92.340 190.260 ;
        RECT 52.390 189.580 52.710 189.640 ;
        RECT 51.100 189.440 52.710 189.580 ;
        RECT 48.725 189.240 49.015 189.285 ;
        RECT 50.090 189.240 50.410 189.300 ;
        RECT 48.725 189.100 50.410 189.240 ;
        RECT 48.725 189.055 49.015 189.100 ;
        RECT 50.090 189.040 50.410 189.100 ;
        RECT 31.690 188.900 32.010 188.960 ;
        RECT 34.910 188.900 35.230 188.960 ;
        RECT 31.690 188.760 35.230 188.900 ;
        RECT 31.690 188.700 32.010 188.760 ;
        RECT 34.910 188.700 35.230 188.760 ;
        RECT 37.225 188.900 37.515 188.945 ;
        RECT 40.430 188.900 40.750 188.960 ;
        RECT 37.225 188.760 42.960 188.900 ;
        RECT 37.225 188.715 37.515 188.760 ;
        RECT 40.430 188.700 40.750 188.760 ;
        RECT 35.370 188.360 35.690 188.620 ;
        RECT 38.590 188.560 38.910 188.620 ;
        RECT 40.905 188.560 41.195 188.605 ;
        RECT 38.590 188.420 41.195 188.560 ;
        RECT 38.590 188.360 38.910 188.420 ;
        RECT 40.905 188.375 41.195 188.420 ;
        RECT 41.825 188.375 42.115 188.605 ;
        RECT 41.900 188.220 42.040 188.375 ;
        RECT 42.270 188.360 42.590 188.620 ;
        RECT 42.820 188.605 42.960 188.760 ;
        RECT 50.550 188.605 50.870 188.620 ;
        RECT 51.100 188.605 51.240 189.440 ;
        RECT 52.390 189.380 52.710 189.440 ;
        RECT 56.530 189.380 56.850 189.640 ;
        RECT 58.830 189.580 59.150 189.640 ;
        RECT 62.050 189.580 62.370 189.640 ;
        RECT 78.610 189.580 78.930 189.640 ;
        RECT 79.085 189.580 79.375 189.625 ;
        RECT 58.830 189.440 71.480 189.580 ;
        RECT 58.830 189.380 59.150 189.440 ;
        RECT 62.050 189.380 62.370 189.440 ;
        RECT 51.930 189.240 52.250 189.300 ;
        RECT 56.620 189.240 56.760 189.380 ;
        RECT 64.390 189.240 64.680 189.285 ;
        RECT 66.490 189.240 66.780 189.285 ;
        RECT 68.060 189.240 68.350 189.285 ;
        RECT 51.930 189.100 56.300 189.240 ;
        RECT 56.620 189.100 58.140 189.240 ;
        RECT 51.930 189.040 52.250 189.100 ;
        RECT 56.160 188.945 56.300 189.100 ;
        RECT 56.085 188.715 56.375 188.945 ;
        RECT 56.990 188.700 57.310 188.960 ;
        RECT 42.745 188.375 43.035 188.605 ;
        RECT 49.645 188.560 49.935 188.605 ;
        RECT 49.260 188.420 49.935 188.560 ;
        RECT 43.650 188.220 43.970 188.280 ;
        RECT 41.900 188.080 43.970 188.220 ;
        RECT 43.650 188.020 43.970 188.080 ;
        RECT 46.870 188.020 47.190 188.280 ;
        RECT 44.110 187.680 44.430 187.940 ;
        RECT 45.490 187.880 45.810 187.940 ;
        RECT 49.260 187.925 49.400 188.420 ;
        RECT 49.645 188.375 49.935 188.420 ;
        RECT 50.385 188.375 50.870 188.605 ;
        RECT 51.025 188.375 51.315 188.605 ;
        RECT 52.175 188.560 52.465 188.605 ;
        RECT 52.850 188.560 53.170 188.620 ;
        RECT 54.245 188.560 54.535 188.605 ;
        RECT 52.175 188.420 54.535 188.560 ;
        RECT 52.175 188.375 52.465 188.420 ;
        RECT 50.550 188.360 50.870 188.375 ;
        RECT 52.850 188.360 53.170 188.420 ;
        RECT 54.245 188.375 54.535 188.420 ;
        RECT 54.705 188.375 54.995 188.605 ;
        RECT 51.485 188.220 51.775 188.265 ;
        RECT 54.780 188.220 54.920 188.375 ;
        RECT 51.485 188.080 54.920 188.220 ;
        RECT 51.485 188.035 51.775 188.080 ;
        RECT 53.860 187.940 54.000 188.080 ;
        RECT 56.070 188.020 56.390 188.280 ;
        RECT 56.545 188.220 56.835 188.265 ;
        RECT 57.080 188.220 57.220 188.700 ;
        RECT 58.000 188.560 58.140 189.100 ;
        RECT 64.390 189.100 68.350 189.240 ;
        RECT 64.390 189.055 64.680 189.100 ;
        RECT 66.490 189.055 66.780 189.100 ;
        RECT 68.060 189.055 68.350 189.100 ;
        RECT 62.970 188.900 63.290 188.960 ;
        RECT 63.905 188.900 64.195 188.945 ;
        RECT 61.220 188.760 62.740 188.900 ;
        RECT 61.220 188.605 61.360 188.760 ;
        RECT 62.600 188.620 62.740 188.760 ;
        RECT 62.970 188.760 64.195 188.900 ;
        RECT 62.970 188.700 63.290 188.760 ;
        RECT 63.905 188.715 64.195 188.760 ;
        RECT 64.785 188.900 65.075 188.945 ;
        RECT 65.975 188.900 66.265 188.945 ;
        RECT 68.495 188.900 68.785 188.945 ;
        RECT 64.785 188.760 68.785 188.900 ;
        RECT 64.785 188.715 65.075 188.760 ;
        RECT 65.975 188.715 66.265 188.760 ;
        RECT 68.495 188.715 68.785 188.760 ;
        RECT 71.340 188.900 71.480 189.440 ;
        RECT 78.610 189.440 79.375 189.580 ;
        RECT 78.610 189.380 78.930 189.440 ;
        RECT 79.085 189.395 79.375 189.440 ;
        RECT 79.990 189.380 80.310 189.640 ;
        RECT 74.025 188.900 74.315 188.945 ;
        RECT 71.340 188.760 74.315 188.900 ;
        RECT 59.075 188.560 59.365 188.605 ;
        RECT 58.000 188.420 59.365 188.560 ;
        RECT 59.075 188.375 59.365 188.420 ;
        RECT 61.140 188.375 61.430 188.605 ;
        RECT 61.590 188.360 61.910 188.620 ;
        RECT 62.510 188.360 62.830 188.620 ;
        RECT 59.765 188.220 60.055 188.265 ;
        RECT 56.545 188.080 57.220 188.220 ;
        RECT 57.540 188.080 60.055 188.220 ;
        RECT 56.545 188.035 56.835 188.080 ;
        RECT 49.185 187.880 49.475 187.925 ;
        RECT 45.490 187.740 49.475 187.880 ;
        RECT 45.490 187.680 45.810 187.740 ;
        RECT 49.185 187.695 49.475 187.740 ;
        RECT 52.850 187.680 53.170 187.940 ;
        RECT 53.310 187.680 53.630 187.940 ;
        RECT 53.770 187.680 54.090 187.940 ;
        RECT 56.160 187.880 56.300 188.020 ;
        RECT 57.540 187.880 57.680 188.080 ;
        RECT 59.765 188.035 60.055 188.080 ;
        RECT 60.210 188.020 60.530 188.280 ;
        RECT 63.890 188.220 64.210 188.280 ;
        RECT 65.130 188.220 65.420 188.265 ;
        RECT 71.340 188.220 71.480 188.760 ;
        RECT 74.025 188.715 74.315 188.760 ;
        RECT 71.710 188.560 72.030 188.620 ;
        RECT 75.865 188.560 76.155 188.605 ;
        RECT 71.710 188.420 76.155 188.560 ;
        RECT 71.710 188.360 72.030 188.420 ;
        RECT 75.865 188.375 76.155 188.420 ;
        RECT 76.785 188.560 77.075 188.605 ;
        RECT 78.700 188.560 78.840 189.380 ;
        RECT 76.785 188.420 78.840 188.560 ;
        RECT 76.785 188.375 77.075 188.420 ;
        RECT 84.605 188.375 84.895 188.605 ;
        RECT 63.890 188.080 65.420 188.220 ;
        RECT 63.890 188.020 64.210 188.080 ;
        RECT 65.130 188.035 65.420 188.080 ;
        RECT 70.880 188.080 71.480 188.220 ;
        RECT 80.910 188.220 81.230 188.280 ;
        RECT 84.680 188.220 84.820 188.375 ;
        RECT 85.050 188.360 85.370 188.620 ;
        RECT 85.510 188.360 85.830 188.620 ;
        RECT 86.430 188.360 86.750 188.620 ;
        RECT 80.910 188.080 84.820 188.220 ;
        RECT 56.160 187.740 57.680 187.880 ;
        RECT 58.370 187.680 58.690 187.940 ;
        RECT 70.880 187.925 71.020 188.080 ;
        RECT 80.910 188.020 81.230 188.080 ;
        RECT 70.805 187.695 71.095 187.925 ;
        RECT 71.250 187.680 71.570 187.940 ;
        RECT 76.325 187.880 76.615 187.925 ;
        RECT 77.690 187.880 78.010 187.940 ;
        RECT 79.990 187.925 80.310 187.940 ;
        RECT 76.325 187.740 78.010 187.880 ;
        RECT 76.325 187.695 76.615 187.740 ;
        RECT 77.690 187.680 78.010 187.740 ;
        RECT 79.925 187.695 80.310 187.925 ;
        RECT 83.225 187.880 83.515 187.925 ;
        RECT 83.670 187.880 83.990 187.940 ;
        RECT 83.225 187.740 83.990 187.880 ;
        RECT 83.225 187.695 83.515 187.740 ;
        RECT 79.990 187.680 80.310 187.695 ;
        RECT 83.670 187.680 83.990 187.740 ;
        RECT 18.280 187.060 93.120 187.540 ;
        RECT 35.370 186.660 35.690 186.920 ;
        RECT 36.765 186.860 37.055 186.905 ;
        RECT 38.590 186.860 38.910 186.920 ;
        RECT 36.765 186.720 38.910 186.860 ;
        RECT 36.765 186.675 37.055 186.720 ;
        RECT 38.590 186.660 38.910 186.720 ;
        RECT 39.525 186.860 39.815 186.905 ;
        RECT 42.270 186.860 42.590 186.920 ;
        RECT 52.390 186.860 52.710 186.920 ;
        RECT 39.525 186.720 42.590 186.860 ;
        RECT 39.525 186.675 39.815 186.720 ;
        RECT 34.465 186.180 34.755 186.225 ;
        RECT 35.460 186.180 35.600 186.660 ;
        RECT 34.465 186.040 35.600 186.180 ;
        RECT 34.465 185.995 34.755 186.040 ;
        RECT 37.210 185.980 37.530 186.240 ;
        RECT 40.060 186.225 40.200 186.720 ;
        RECT 42.270 186.660 42.590 186.720 ;
        RECT 48.800 186.720 52.710 186.860 ;
        RECT 39.985 185.995 40.275 186.225 ;
        RECT 44.110 186.180 44.430 186.240 ;
        RECT 45.045 186.180 45.335 186.225 ;
        RECT 44.110 186.040 45.335 186.180 ;
        RECT 44.110 185.980 44.430 186.040 ;
        RECT 45.045 185.995 45.335 186.040 ;
        RECT 45.490 185.980 45.810 186.240 ;
        RECT 48.800 186.225 48.940 186.720 ;
        RECT 52.390 186.660 52.710 186.720 ;
        RECT 54.245 186.860 54.535 186.905 ;
        RECT 58.370 186.860 58.690 186.920 ;
        RECT 54.245 186.720 58.690 186.860 ;
        RECT 54.245 186.675 54.535 186.720 ;
        RECT 58.370 186.660 58.690 186.720 ;
        RECT 60.210 186.660 60.530 186.920 ;
        RECT 63.890 186.660 64.210 186.920 ;
        RECT 74.930 186.660 75.250 186.920 ;
        RECT 80.465 186.860 80.755 186.905 ;
        RECT 85.510 186.860 85.830 186.920 ;
        RECT 80.465 186.720 85.830 186.860 ;
        RECT 80.465 186.675 80.755 186.720 ;
        RECT 85.510 186.660 85.830 186.720 ;
        RECT 49.260 186.380 54.000 186.520 ;
        RECT 49.260 186.225 49.400 186.380 ;
        RECT 53.860 186.240 54.000 186.380 ;
        RECT 58.830 186.320 59.150 186.580 ;
        RECT 68.045 186.520 68.335 186.565 ;
        RECT 83.230 186.520 83.520 186.565 ;
        RECT 84.630 186.520 84.920 186.565 ;
        RECT 86.470 186.520 86.760 186.565 ;
        RECT 64.900 186.380 68.335 186.520 ;
        RECT 46.425 185.995 46.715 186.225 ;
        RECT 48.725 185.995 49.015 186.225 ;
        RECT 49.185 185.995 49.475 186.225 ;
        RECT 41.350 185.640 41.670 185.900 ;
        RECT 46.500 185.840 46.640 185.995 ;
        RECT 50.550 185.980 50.870 186.240 ;
        RECT 52.405 186.180 52.695 186.225 ;
        RECT 52.850 186.180 53.170 186.240 ;
        RECT 52.405 186.040 53.170 186.180 ;
        RECT 52.405 185.995 52.695 186.040 ;
        RECT 52.850 185.980 53.170 186.040 ;
        RECT 53.310 185.980 53.630 186.240 ;
        RECT 53.770 185.980 54.090 186.240 ;
        RECT 54.705 186.180 54.995 186.225 ;
        RECT 57.450 186.180 57.770 186.240 ;
        RECT 54.705 186.040 57.770 186.180 ;
        RECT 54.705 185.995 54.995 186.040 ;
        RECT 57.450 185.980 57.770 186.040 ;
        RECT 57.925 186.180 58.215 186.225 ;
        RECT 58.920 186.180 59.060 186.320 ;
        RECT 64.900 186.225 65.040 186.380 ;
        RECT 68.045 186.335 68.335 186.380 ;
        RECT 75.940 186.380 79.760 186.520 ;
        RECT 75.940 186.240 76.080 186.380 ;
        RECT 57.925 186.040 59.060 186.180 ;
        RECT 57.925 185.995 58.215 186.040 ;
        RECT 64.825 185.995 65.115 186.225 ;
        RECT 42.820 185.700 52.160 185.840 ;
        RECT 42.820 185.545 42.960 185.700 ;
        RECT 42.745 185.315 43.035 185.545 ;
        RECT 45.965 185.500 46.255 185.545 ;
        RECT 47.805 185.500 48.095 185.545 ;
        RECT 45.965 185.360 48.095 185.500 ;
        RECT 45.965 185.315 46.255 185.360 ;
        RECT 47.805 185.315 48.095 185.360 ;
        RECT 50.090 185.300 50.410 185.560 ;
        RECT 34.910 184.960 35.230 185.220 ;
        RECT 38.605 185.160 38.895 185.205 ;
        RECT 39.510 185.160 39.830 185.220 ;
        RECT 38.605 185.020 39.830 185.160 ;
        RECT 38.605 184.975 38.895 185.020 ;
        RECT 39.510 184.960 39.830 185.020 ;
        RECT 40.430 184.960 40.750 185.220 ;
        RECT 47.330 184.960 47.650 185.220 ;
        RECT 51.025 185.160 51.315 185.205 ;
        RECT 51.470 185.160 51.790 185.220 ;
        RECT 51.025 185.020 51.790 185.160 ;
        RECT 52.020 185.160 52.160 185.700 ;
        RECT 52.865 185.500 53.155 185.545 ;
        RECT 53.400 185.500 53.540 185.980 ;
        RECT 52.865 185.360 53.540 185.500 ;
        RECT 57.450 185.500 57.770 185.560 ;
        RECT 58.000 185.500 58.140 185.995 ;
        RECT 66.190 185.980 66.510 186.240 ;
        RECT 67.125 185.995 67.415 186.225 ;
        RECT 68.505 186.180 68.795 186.225 ;
        RECT 71.250 186.180 71.570 186.240 ;
        RECT 68.505 186.040 71.570 186.180 ;
        RECT 68.505 185.995 68.795 186.040 ;
        RECT 57.450 185.360 58.140 185.500 ;
        RECT 62.970 185.500 63.290 185.560 ;
        RECT 65.285 185.500 65.575 185.545 ;
        RECT 62.970 185.360 65.575 185.500 ;
        RECT 52.865 185.315 53.155 185.360 ;
        RECT 57.450 185.300 57.770 185.360 ;
        RECT 62.970 185.300 63.290 185.360 ;
        RECT 65.285 185.315 65.575 185.360 ;
        RECT 65.730 185.300 66.050 185.560 ;
        RECT 67.200 185.220 67.340 185.995 ;
        RECT 71.250 185.980 71.570 186.040 ;
        RECT 75.850 185.980 76.170 186.240 ;
        RECT 77.230 185.980 77.550 186.240 ;
        RECT 77.690 186.180 78.010 186.240 ;
        RECT 77.690 186.040 78.205 186.180 ;
        RECT 77.690 185.980 78.010 186.040 ;
        RECT 78.610 185.980 78.930 186.240 ;
        RECT 79.070 185.980 79.390 186.240 ;
        RECT 79.620 186.225 79.760 186.380 ;
        RECT 83.230 186.380 86.760 186.520 ;
        RECT 83.230 186.335 83.520 186.380 ;
        RECT 84.630 186.335 84.920 186.380 ;
        RECT 86.470 186.335 86.760 186.380 ;
        RECT 79.570 185.995 79.860 186.225 ;
        RECT 81.830 186.180 82.150 186.240 ;
        RECT 82.305 186.180 82.595 186.225 ;
        RECT 81.830 186.040 82.595 186.180 ;
        RECT 81.830 185.980 82.150 186.040 ;
        RECT 82.305 185.995 82.595 186.040 ;
        RECT 83.670 185.980 83.990 186.240 ;
        RECT 72.630 185.840 72.950 185.900 ;
        RECT 73.565 185.840 73.855 185.885 ;
        RECT 72.630 185.700 73.855 185.840 ;
        RECT 72.630 185.640 72.950 185.700 ;
        RECT 73.565 185.655 73.855 185.700 ;
        RECT 74.485 185.840 74.775 185.885 ;
        RECT 81.370 185.840 81.690 185.900 ;
        RECT 91.030 185.840 91.350 185.900 ;
        RECT 74.485 185.700 81.690 185.840 ;
        RECT 74.485 185.655 74.775 185.700 ;
        RECT 81.370 185.640 81.690 185.700 ;
        RECT 81.920 185.700 91.350 185.840 ;
        RECT 80.910 185.500 81.230 185.560 ;
        RECT 81.920 185.500 82.060 185.700 ;
        RECT 91.030 185.640 91.350 185.700 ;
        RECT 80.910 185.360 82.060 185.500 ;
        RECT 82.770 185.500 83.060 185.545 ;
        RECT 85.090 185.500 85.380 185.545 ;
        RECT 86.470 185.500 86.760 185.545 ;
        RECT 82.770 185.360 86.760 185.500 ;
        RECT 80.910 185.300 81.230 185.360 ;
        RECT 82.770 185.315 83.060 185.360 ;
        RECT 85.090 185.315 85.380 185.360 ;
        RECT 86.470 185.315 86.760 185.360 ;
        RECT 53.325 185.160 53.615 185.205 ;
        RECT 52.020 185.020 53.615 185.160 ;
        RECT 51.025 184.975 51.315 185.020 ;
        RECT 51.470 184.960 51.790 185.020 ;
        RECT 53.325 184.975 53.615 185.020 ;
        RECT 59.290 184.960 59.610 185.220 ;
        RECT 62.510 185.160 62.830 185.220 ;
        RECT 67.110 185.160 67.430 185.220 ;
        RECT 62.510 185.020 67.430 185.160 ;
        RECT 62.510 184.960 62.830 185.020 ;
        RECT 67.110 184.960 67.430 185.020 ;
        RECT 76.785 185.160 77.075 185.205 ;
        RECT 77.690 185.160 78.010 185.220 ;
        RECT 76.785 185.020 78.010 185.160 ;
        RECT 76.785 184.975 77.075 185.020 ;
        RECT 77.690 184.960 78.010 185.020 ;
        RECT 90.125 185.160 90.415 185.205 ;
        RECT 91.030 185.160 91.350 185.220 ;
        RECT 90.125 185.020 91.350 185.160 ;
        RECT 90.125 184.975 90.415 185.020 ;
        RECT 91.030 184.960 91.350 185.020 ;
        RECT 18.280 184.340 92.340 184.820 ;
        RECT 40.445 184.140 40.735 184.185 ;
        RECT 41.350 184.140 41.670 184.200 ;
        RECT 40.445 184.000 41.670 184.140 ;
        RECT 40.445 183.955 40.735 184.000 ;
        RECT 41.350 183.940 41.670 184.000 ;
        RECT 41.810 184.140 42.130 184.200 ;
        RECT 43.205 184.140 43.495 184.185 ;
        RECT 41.810 184.000 43.495 184.140 ;
        RECT 41.810 183.940 42.130 184.000 ;
        RECT 43.205 183.955 43.495 184.000 ;
        RECT 66.190 184.140 66.510 184.200 ;
        RECT 67.125 184.140 67.415 184.185 ;
        RECT 66.190 184.000 67.415 184.140 ;
        RECT 66.190 183.940 66.510 184.000 ;
        RECT 67.125 183.955 67.415 184.000 ;
        RECT 78.610 183.940 78.930 184.200 ;
        RECT 80.910 184.140 81.230 184.200 ;
        RECT 79.160 184.000 81.230 184.140 ;
        RECT 39.510 183.600 39.830 183.860 ;
        RECT 58.370 183.800 58.690 183.860 ;
        RECT 58.370 183.660 65.960 183.800 ;
        RECT 58.370 183.600 58.690 183.660 ;
        RECT 37.210 183.460 37.530 183.520 ;
        RECT 38.145 183.460 38.435 183.505 ;
        RECT 58.830 183.460 59.150 183.520 ;
        RECT 65.820 183.505 65.960 183.660 ;
        RECT 65.285 183.460 65.575 183.505 ;
        RECT 37.210 183.320 65.575 183.460 ;
        RECT 37.210 183.260 37.530 183.320 ;
        RECT 38.145 183.275 38.435 183.320 ;
        RECT 58.830 183.260 59.150 183.320 ;
        RECT 65.285 183.275 65.575 183.320 ;
        RECT 65.745 183.460 66.035 183.505 ;
        RECT 77.230 183.460 77.550 183.520 ;
        RECT 65.745 183.320 77.550 183.460 ;
        RECT 65.745 183.275 66.035 183.320 ;
        RECT 77.230 183.260 77.550 183.320 ;
        RECT 62.050 183.120 62.370 183.180 ;
        RECT 64.825 183.120 65.115 183.165 ;
        RECT 62.050 182.980 65.115 183.120 ;
        RECT 62.050 182.920 62.370 182.980 ;
        RECT 64.825 182.935 65.115 182.980 ;
        RECT 66.190 182.920 66.510 183.180 ;
        RECT 79.160 183.120 79.300 184.000 ;
        RECT 80.910 183.940 81.230 184.000 ;
        RECT 81.370 184.140 81.690 184.200 ;
        RECT 81.845 184.140 82.135 184.185 ;
        RECT 81.370 184.000 82.135 184.140 ;
        RECT 81.370 183.940 81.690 184.000 ;
        RECT 81.845 183.955 82.135 184.000 ;
        RECT 79.530 183.600 79.850 183.860 ;
        RECT 79.620 183.460 79.760 183.600 ;
        RECT 79.620 183.320 81.600 183.460 ;
        RECT 79.545 183.120 79.835 183.165 ;
        RECT 79.160 182.980 79.835 183.120 ;
        RECT 79.545 182.935 79.835 182.980 ;
        RECT 79.990 183.120 80.310 183.180 ;
        RECT 80.910 183.120 81.230 183.180 ;
        RECT 81.460 183.165 81.600 183.320 ;
        RECT 79.990 182.980 81.230 183.120 ;
        RECT 79.990 182.920 80.310 182.980 ;
        RECT 80.910 182.920 81.230 182.980 ;
        RECT 81.385 182.935 81.675 183.165 ;
        RECT 82.305 182.935 82.595 183.165 ;
        RECT 50.565 182.780 50.855 182.825 ;
        RECT 60.210 182.780 60.530 182.840 ;
        RECT 67.585 182.780 67.875 182.825 ;
        RECT 50.565 182.640 67.875 182.780 ;
        RECT 50.565 182.595 50.855 182.640 ;
        RECT 60.210 182.580 60.530 182.640 ;
        RECT 67.585 182.595 67.875 182.640 ;
        RECT 75.850 182.780 76.170 182.840 ;
        RECT 76.325 182.780 76.615 182.825 ;
        RECT 81.830 182.780 82.150 182.840 ;
        RECT 75.850 182.640 82.150 182.780 ;
        RECT 75.850 182.580 76.170 182.640 ;
        RECT 76.325 182.595 76.615 182.640 ;
        RECT 81.830 182.580 82.150 182.640 ;
        RECT 48.250 182.440 48.570 182.500 ;
        RECT 66.650 182.440 66.970 182.500 ;
        RECT 48.250 182.300 66.970 182.440 ;
        RECT 48.250 182.240 48.570 182.300 ;
        RECT 66.650 182.240 66.970 182.300 ;
        RECT 79.990 182.440 80.310 182.500 ;
        RECT 80.465 182.440 80.755 182.485 ;
        RECT 79.990 182.300 80.755 182.440 ;
        RECT 79.990 182.240 80.310 182.300 ;
        RECT 80.465 182.255 80.755 182.300 ;
        RECT 80.910 182.440 81.230 182.500 ;
        RECT 82.380 182.440 82.520 182.935 ;
        RECT 80.910 182.300 82.520 182.440 ;
        RECT 80.910 182.240 81.230 182.300 ;
        RECT 18.280 181.620 93.120 182.100 ;
        RECT 43.190 181.420 43.510 181.480 ;
        RECT 48.250 181.420 48.570 181.480 ;
        RECT 43.190 181.280 48.570 181.420 ;
        RECT 43.190 181.220 43.510 181.280 ;
        RECT 48.250 181.220 48.570 181.280 ;
        RECT 50.550 181.420 50.870 181.480 ;
        RECT 52.390 181.420 52.710 181.480 ;
        RECT 50.550 181.280 52.710 181.420 ;
        RECT 50.550 181.220 50.870 181.280 ;
        RECT 52.390 181.220 52.710 181.280 ;
        RECT 53.770 181.220 54.090 181.480 ;
        RECT 58.370 181.220 58.690 181.480 ;
        RECT 58.830 181.420 59.150 181.480 ;
        RECT 64.825 181.420 65.115 181.465 ;
        RECT 58.830 181.280 65.115 181.420 ;
        RECT 58.830 181.220 59.150 181.280 ;
        RECT 64.825 181.235 65.115 181.280 ;
        RECT 69.870 181.420 70.190 181.480 ;
        RECT 72.645 181.420 72.935 181.465 ;
        RECT 85.970 181.420 86.290 181.480 ;
        RECT 69.870 181.280 72.935 181.420 ;
        RECT 69.870 181.220 70.190 181.280 ;
        RECT 72.645 181.235 72.935 181.280 ;
        RECT 77.320 181.280 86.290 181.420 ;
        RECT 43.650 181.080 43.970 181.140 ;
        RECT 45.045 181.080 45.335 181.125 ;
        RECT 47.805 181.080 48.095 181.125 ;
        RECT 43.650 180.940 48.095 181.080 ;
        RECT 43.650 180.880 43.970 180.940 ;
        RECT 45.045 180.895 45.335 180.940 ;
        RECT 47.805 180.895 48.095 180.940 ;
        RECT 41.365 180.555 41.655 180.785 ;
        RECT 42.285 180.740 42.575 180.785 ;
        RECT 44.570 180.740 44.890 180.800 ;
        RECT 42.285 180.600 44.890 180.740 ;
        RECT 42.285 180.555 42.575 180.600 ;
        RECT 41.440 180.400 41.580 180.555 ;
        RECT 44.570 180.540 44.890 180.600 ;
        RECT 46.870 180.540 47.190 180.800 ;
        RECT 48.340 180.785 48.480 181.220 ;
        RECT 53.310 181.080 53.630 181.140 ;
        RECT 66.190 181.080 66.510 181.140 ;
        RECT 53.310 180.940 66.510 181.080 ;
        RECT 53.310 180.880 53.630 180.940 ;
        RECT 48.265 180.555 48.555 180.785 ;
        RECT 52.865 180.555 53.155 180.785 ;
        RECT 42.730 180.400 43.050 180.460 ;
        RECT 41.440 180.260 43.050 180.400 ;
        RECT 46.960 180.400 47.100 180.540 ;
        RECT 50.090 180.400 50.410 180.460 ;
        RECT 52.940 180.400 53.080 180.555 ;
        RECT 54.230 180.540 54.550 180.800 ;
        RECT 57.910 180.540 58.230 180.800 ;
        RECT 58.830 180.740 59.150 180.800 ;
        RECT 59.305 180.740 59.595 180.785 ;
        RECT 60.685 180.740 60.975 180.785 ;
        RECT 58.830 180.600 59.595 180.740 ;
        RECT 58.830 180.540 59.150 180.600 ;
        RECT 59.305 180.555 59.595 180.600 ;
        RECT 59.840 180.600 60.975 180.740 ;
        RECT 46.960 180.260 53.080 180.400 ;
        RECT 42.730 180.200 43.050 180.260 ;
        RECT 50.090 180.200 50.410 180.260 ;
        RECT 59.840 180.060 59.980 180.600 ;
        RECT 60.685 180.555 60.975 180.600 ;
        RECT 61.605 180.555 61.895 180.785 ;
        RECT 62.065 180.555 62.355 180.785 ;
        RECT 60.225 180.400 60.515 180.445 ;
        RECT 61.680 180.400 61.820 180.555 ;
        RECT 60.225 180.260 61.820 180.400 ;
        RECT 62.140 180.400 62.280 180.555 ;
        RECT 62.510 180.540 62.830 180.800 ;
        RECT 64.440 180.785 64.580 180.940 ;
        RECT 66.190 180.880 66.510 180.940 ;
        RECT 66.650 181.080 66.970 181.140 ;
        RECT 71.250 181.080 71.570 181.140 ;
        RECT 72.185 181.080 72.475 181.125 ;
        RECT 76.310 181.080 76.630 181.140 ;
        RECT 66.650 180.940 76.630 181.080 ;
        RECT 66.650 180.880 66.970 180.940 ;
        RECT 71.250 180.880 71.570 180.940 ;
        RECT 72.185 180.895 72.475 180.940 ;
        RECT 76.310 180.880 76.630 180.940 ;
        RECT 64.365 180.555 64.655 180.785 ;
        RECT 65.745 180.555 66.035 180.785 ;
        RECT 67.110 180.740 67.430 180.800 ;
        RECT 76.785 180.740 77.075 180.785 ;
        RECT 77.320 180.740 77.460 181.280 ;
        RECT 85.970 181.220 86.290 181.280 ;
        RECT 83.230 181.080 83.520 181.125 ;
        RECT 84.630 181.080 84.920 181.125 ;
        RECT 86.470 181.080 86.760 181.125 ;
        RECT 78.240 180.940 80.220 181.080 ;
        RECT 67.110 180.600 77.460 180.740 ;
        RECT 65.820 180.400 65.960 180.555 ;
        RECT 67.110 180.540 67.430 180.600 ;
        RECT 76.785 180.555 77.075 180.600 ;
        RECT 77.690 180.540 78.010 180.800 ;
        RECT 70.790 180.400 71.110 180.460 ;
        RECT 78.240 180.445 78.380 180.940 ;
        RECT 79.530 180.540 79.850 180.800 ;
        RECT 80.080 180.730 80.220 180.940 ;
        RECT 83.230 180.940 86.760 181.080 ;
        RECT 83.230 180.895 83.520 180.940 ;
        RECT 84.630 180.895 84.920 180.940 ;
        RECT 86.470 180.895 86.760 180.940 ;
        RECT 80.865 180.770 81.155 180.785 ;
        RECT 80.540 180.730 81.155 180.770 ;
        RECT 80.080 180.630 81.155 180.730 ;
        RECT 80.080 180.590 80.680 180.630 ;
        RECT 80.865 180.555 81.155 180.630 ;
        RECT 81.385 180.555 81.675 180.785 ;
        RECT 81.845 180.555 82.135 180.785 ;
        RECT 78.165 180.400 78.455 180.445 ;
        RECT 62.140 180.260 62.740 180.400 ;
        RECT 65.820 180.260 71.110 180.400 ;
        RECT 60.225 180.215 60.515 180.260 ;
        RECT 62.050 180.060 62.370 180.120 ;
        RECT 59.840 179.920 62.370 180.060 ;
        RECT 62.050 179.860 62.370 179.920 ;
        RECT 41.350 179.720 41.670 179.780 ;
        RECT 42.285 179.720 42.575 179.765 ;
        RECT 41.350 179.580 42.575 179.720 ;
        RECT 41.350 179.520 41.670 179.580 ;
        RECT 42.285 179.535 42.575 179.580 ;
        RECT 46.425 179.720 46.715 179.765 ;
        RECT 48.710 179.720 49.030 179.780 ;
        RECT 46.425 179.580 49.030 179.720 ;
        RECT 62.600 179.720 62.740 180.260 ;
        RECT 70.790 180.200 71.110 180.260 ;
        RECT 77.780 180.260 78.455 180.400 ;
        RECT 63.905 180.060 64.195 180.105 ;
        RECT 66.190 180.060 66.510 180.120 ;
        RECT 63.905 179.920 66.510 180.060 ;
        RECT 63.905 179.875 64.195 179.920 ;
        RECT 66.190 179.860 66.510 179.920 ;
        RECT 77.780 179.780 77.920 180.260 ;
        RECT 78.165 180.215 78.455 180.260 ;
        RECT 78.625 180.400 78.915 180.445 ;
        RECT 81.460 180.400 81.600 180.555 ;
        RECT 78.625 180.260 81.600 180.400 ;
        RECT 78.625 180.215 78.915 180.260 ;
        RECT 79.530 180.060 79.850 180.120 ;
        RECT 79.530 179.920 80.220 180.060 ;
        RECT 79.530 179.860 79.850 179.920 ;
        RECT 65.730 179.720 66.050 179.780 ;
        RECT 62.600 179.580 66.050 179.720 ;
        RECT 46.425 179.535 46.715 179.580 ;
        RECT 48.710 179.520 49.030 179.580 ;
        RECT 65.730 179.520 66.050 179.580 ;
        RECT 77.690 179.520 78.010 179.780 ;
        RECT 80.080 179.720 80.220 179.920 ;
        RECT 80.465 179.875 80.755 180.105 ;
        RECT 81.370 180.060 81.690 180.120 ;
        RECT 81.920 180.060 82.060 180.555 ;
        RECT 82.750 180.540 83.070 180.800 ;
        RECT 82.290 180.200 82.610 180.460 ;
        RECT 82.840 180.400 82.980 180.540 ;
        RECT 83.685 180.400 83.975 180.445 ;
        RECT 82.840 180.260 83.975 180.400 ;
        RECT 83.685 180.215 83.975 180.260 ;
        RECT 81.370 179.920 82.060 180.060 ;
        RECT 82.770 180.060 83.060 180.105 ;
        RECT 85.090 180.060 85.380 180.105 ;
        RECT 86.470 180.060 86.760 180.105 ;
        RECT 82.770 179.920 86.760 180.060 ;
        RECT 80.540 179.720 80.680 179.875 ;
        RECT 81.370 179.860 81.690 179.920 ;
        RECT 82.770 179.875 83.060 179.920 ;
        RECT 85.090 179.875 85.380 179.920 ;
        RECT 86.470 179.875 86.760 179.920 ;
        RECT 80.080 179.580 80.680 179.720 ;
        RECT 90.125 179.720 90.415 179.765 ;
        RECT 91.030 179.720 91.350 179.780 ;
        RECT 90.125 179.580 91.350 179.720 ;
        RECT 90.125 179.535 90.415 179.580 ;
        RECT 91.030 179.520 91.350 179.580 ;
        RECT 18.280 178.900 92.340 179.380 ;
        RECT 41.810 178.700 42.130 178.760 ;
        RECT 40.060 178.560 42.130 178.700 ;
        RECT 40.060 178.065 40.200 178.560 ;
        RECT 41.810 178.500 42.130 178.560 ;
        RECT 44.570 178.700 44.890 178.760 ;
        RECT 49.185 178.700 49.475 178.745 ;
        RECT 44.570 178.560 49.475 178.700 ;
        RECT 44.570 178.500 44.890 178.560 ;
        RECT 49.185 178.515 49.475 178.560 ;
        RECT 53.310 178.500 53.630 178.760 ;
        RECT 54.230 178.500 54.550 178.760 ;
        RECT 57.910 178.500 58.230 178.760 ;
        RECT 58.370 178.500 58.690 178.760 ;
        RECT 58.830 178.700 59.150 178.760 ;
        RECT 62.065 178.700 62.355 178.745 ;
        RECT 58.830 178.560 62.355 178.700 ;
        RECT 58.830 178.500 59.150 178.560 ;
        RECT 62.065 178.515 62.355 178.560 ;
        RECT 71.710 178.700 72.030 178.760 ;
        RECT 72.185 178.700 72.475 178.745 ;
        RECT 81.370 178.700 81.690 178.760 ;
        RECT 82.305 178.700 82.595 178.745 ;
        RECT 71.710 178.560 72.475 178.700 ;
        RECT 71.710 178.500 72.030 178.560 ;
        RECT 72.185 178.515 72.475 178.560 ;
        RECT 79.160 178.560 82.595 178.700 ;
        RECT 40.470 178.360 40.760 178.405 ;
        RECT 42.570 178.360 42.860 178.405 ;
        RECT 44.140 178.360 44.430 178.405 ;
        RECT 40.470 178.220 44.430 178.360 ;
        RECT 40.470 178.175 40.760 178.220 ;
        RECT 42.570 178.175 42.860 178.220 ;
        RECT 44.140 178.175 44.430 178.220 ;
        RECT 46.870 178.160 47.190 178.420 ;
        RECT 39.985 177.835 40.275 178.065 ;
        RECT 40.865 178.020 41.155 178.065 ;
        RECT 42.055 178.020 42.345 178.065 ;
        RECT 44.575 178.020 44.865 178.065 ;
        RECT 40.865 177.880 44.865 178.020 ;
        RECT 40.865 177.835 41.155 177.880 ;
        RECT 42.055 177.835 42.345 177.880 ;
        RECT 44.575 177.835 44.865 177.880 ;
        RECT 51.025 178.020 51.315 178.065 ;
        RECT 53.400 178.020 53.540 178.500 ;
        RECT 51.025 177.880 53.540 178.020 ;
        RECT 54.320 178.020 54.460 178.500 ;
        RECT 58.000 178.360 58.140 178.500 ;
        RECT 59.305 178.360 59.595 178.405 ;
        RECT 58.000 178.220 59.595 178.360 ;
        RECT 59.305 178.175 59.595 178.220 ;
        RECT 64.810 178.360 65.100 178.405 ;
        RECT 66.380 178.360 66.670 178.405 ;
        RECT 68.480 178.360 68.770 178.405 ;
        RECT 64.810 178.220 68.770 178.360 ;
        RECT 64.810 178.175 65.100 178.220 ;
        RECT 66.380 178.175 66.670 178.220 ;
        RECT 68.480 178.175 68.770 178.220 ;
        RECT 69.870 178.360 70.190 178.420 ;
        RECT 78.610 178.360 78.930 178.420 ;
        RECT 69.870 178.220 78.930 178.360 ;
        RECT 69.870 178.160 70.190 178.220 ;
        RECT 78.610 178.160 78.930 178.220 ;
        RECT 58.370 178.020 58.690 178.080 ;
        RECT 54.320 177.880 58.690 178.020 ;
        RECT 51.025 177.835 51.315 177.880 ;
        RECT 58.370 177.820 58.690 177.880 ;
        RECT 64.375 178.020 64.665 178.065 ;
        RECT 66.895 178.020 67.185 178.065 ;
        RECT 68.085 178.020 68.375 178.065 ;
        RECT 64.375 177.880 68.375 178.020 ;
        RECT 64.375 177.835 64.665 177.880 ;
        RECT 66.895 177.835 67.185 177.880 ;
        RECT 68.085 177.835 68.375 177.880 ;
        RECT 68.965 178.020 69.255 178.065 ;
        RECT 75.850 178.020 76.170 178.080 ;
        RECT 68.965 177.880 76.170 178.020 ;
        RECT 68.965 177.835 69.255 177.880 ;
        RECT 75.850 177.820 76.170 177.880 ;
        RECT 41.350 177.725 41.670 177.740 ;
        RECT 41.320 177.680 41.670 177.725 ;
        RECT 50.105 177.680 50.395 177.725 ;
        RECT 41.155 177.540 41.670 177.680 ;
        RECT 41.320 177.495 41.670 177.540 ;
        RECT 41.350 177.480 41.670 177.495 ;
        RECT 47.880 177.540 50.395 177.680 ;
        RECT 47.880 177.060 48.020 177.540 ;
        RECT 50.105 177.495 50.395 177.540 ;
        RECT 50.550 177.480 50.870 177.740 ;
        RECT 51.485 177.680 51.775 177.725 ;
        RECT 51.930 177.680 52.250 177.740 ;
        RECT 51.485 177.540 52.250 177.680 ;
        RECT 51.485 177.495 51.775 177.540 ;
        RECT 51.930 177.480 52.250 177.540 ;
        RECT 52.390 177.480 52.710 177.740 ;
        RECT 66.190 177.680 66.510 177.740 ;
        RECT 67.630 177.680 67.920 177.725 ;
        RECT 66.190 177.540 67.920 177.680 ;
        RECT 66.190 177.480 66.510 177.540 ;
        RECT 67.630 177.495 67.920 177.540 ;
        RECT 69.410 177.480 69.730 177.740 ;
        RECT 69.870 177.680 70.190 177.740 ;
        RECT 70.345 177.680 70.635 177.725 ;
        RECT 69.870 177.540 70.635 177.680 ;
        RECT 69.870 177.480 70.190 177.540 ;
        RECT 70.345 177.495 70.635 177.540 ;
        RECT 71.250 177.480 71.570 177.740 ;
        RECT 77.690 177.480 78.010 177.740 ;
        RECT 78.610 177.725 78.930 177.740 ;
        RECT 79.160 177.725 79.300 178.560 ;
        RECT 81.370 178.500 81.690 178.560 ;
        RECT 82.305 178.515 82.595 178.560 ;
        RECT 80.925 178.360 81.215 178.405 ;
        RECT 80.925 178.220 85.740 178.360 ;
        RECT 80.925 178.175 81.215 178.220 ;
        RECT 78.445 177.495 78.930 177.725 ;
        RECT 79.085 177.495 79.375 177.725 ;
        RECT 78.610 177.480 78.930 177.495 ;
        RECT 79.530 177.480 79.850 177.740 ;
        RECT 80.030 177.495 80.320 177.725 ;
        RECT 55.165 177.340 55.455 177.385 ;
        RECT 56.990 177.340 57.310 177.400 ;
        RECT 57.465 177.340 57.755 177.385 ;
        RECT 50.180 177.200 57.755 177.340 ;
        RECT 50.180 177.060 50.320 177.200 ;
        RECT 55.165 177.155 55.455 177.200 ;
        RECT 56.990 177.140 57.310 177.200 ;
        RECT 57.465 177.155 57.755 177.200 ;
        RECT 60.670 177.340 60.990 177.400 ;
        RECT 60.670 177.200 78.840 177.340 ;
        RECT 60.670 177.140 60.990 177.200 ;
        RECT 47.790 176.800 48.110 177.060 ;
        RECT 50.090 176.800 50.410 177.060 ;
        RECT 52.850 177.000 53.170 177.060 ;
        RECT 54.115 177.000 54.405 177.045 ;
        RECT 52.850 176.860 54.405 177.000 ;
        RECT 52.850 176.800 53.170 176.860 ;
        RECT 54.115 176.815 54.405 176.860 ;
        RECT 58.515 177.000 58.805 177.045 ;
        RECT 61.130 177.000 61.450 177.060 ;
        RECT 58.515 176.860 61.450 177.000 ;
        RECT 58.515 176.815 58.805 176.860 ;
        RECT 61.130 176.800 61.450 176.860 ;
        RECT 62.510 177.000 62.830 177.060 ;
        RECT 69.870 177.000 70.190 177.060 ;
        RECT 62.510 176.860 70.190 177.000 ;
        RECT 62.510 176.800 62.830 176.860 ;
        RECT 69.870 176.800 70.190 176.860 ;
        RECT 70.330 176.800 70.650 177.060 ;
        RECT 78.700 177.000 78.840 177.200 ;
        RECT 80.080 177.000 80.220 177.495 ;
        RECT 81.370 177.480 81.690 177.740 ;
        RECT 82.305 177.495 82.595 177.725 ;
        RECT 84.605 177.495 84.895 177.725 ;
        RECT 82.380 177.340 82.520 177.495 ;
        RECT 81.460 177.200 82.520 177.340 ;
        RECT 84.680 177.340 84.820 177.495 ;
        RECT 85.050 177.480 85.370 177.740 ;
        RECT 85.600 177.725 85.740 178.220 ;
        RECT 85.525 177.495 85.815 177.725 ;
        RECT 85.970 177.680 86.290 177.740 ;
        RECT 86.445 177.680 86.735 177.725 ;
        RECT 85.970 177.540 86.735 177.680 ;
        RECT 85.970 177.480 86.290 177.540 ;
        RECT 86.445 177.495 86.735 177.540 ;
        RECT 90.110 177.480 90.430 177.740 ;
        RECT 90.200 177.340 90.340 177.480 ;
        RECT 84.680 177.200 90.340 177.340 ;
        RECT 81.460 177.060 81.600 177.200 ;
        RECT 78.700 176.860 80.220 177.000 ;
        RECT 81.370 176.800 81.690 177.060 ;
        RECT 83.225 177.000 83.515 177.045 ;
        RECT 83.670 177.000 83.990 177.060 ;
        RECT 83.225 176.860 83.990 177.000 ;
        RECT 83.225 176.815 83.515 176.860 ;
        RECT 83.670 176.800 83.990 176.860 ;
        RECT 18.280 176.180 93.120 176.660 ;
        RECT 41.810 175.780 42.130 176.040 ;
        RECT 42.730 175.780 43.050 176.040 ;
        RECT 49.645 175.980 49.935 176.025 ;
        RECT 51.010 175.980 51.330 176.040 ;
        RECT 49.645 175.840 51.330 175.980 ;
        RECT 49.645 175.795 49.935 175.840 ;
        RECT 41.900 175.640 42.040 175.780 ;
        RECT 42.820 175.640 42.960 175.780 ;
        RECT 47.790 175.640 48.110 175.700 ;
        RECT 49.720 175.640 49.860 175.795 ;
        RECT 51.010 175.780 51.330 175.840 ;
        RECT 53.785 175.980 54.075 176.025 ;
        RECT 56.530 175.980 56.850 176.040 ;
        RECT 73.090 175.980 73.410 176.040 ;
        RECT 53.785 175.840 56.850 175.980 ;
        RECT 53.785 175.795 54.075 175.840 ;
        RECT 56.530 175.780 56.850 175.840 ;
        RECT 66.740 175.840 73.410 175.980 ;
        RECT 41.440 175.500 42.040 175.640 ;
        RECT 42.360 175.500 42.960 175.640 ;
        RECT 46.500 175.500 48.110 175.640 ;
        RECT 41.440 175.345 41.580 175.500 ;
        RECT 40.085 175.300 40.375 175.345 ;
        RECT 40.085 175.160 41.120 175.300 ;
        RECT 40.085 175.115 40.375 175.160 ;
        RECT 36.775 174.960 37.065 175.005 ;
        RECT 39.295 174.960 39.585 175.005 ;
        RECT 40.485 174.960 40.775 175.005 ;
        RECT 36.775 174.820 40.775 174.960 ;
        RECT 40.980 174.960 41.120 175.160 ;
        RECT 41.365 175.115 41.655 175.345 ;
        RECT 41.825 175.300 42.115 175.345 ;
        RECT 42.360 175.300 42.500 175.500 ;
        RECT 46.500 175.345 46.640 175.500 ;
        RECT 47.790 175.440 48.110 175.500 ;
        RECT 48.800 175.500 49.860 175.640 ;
        RECT 41.825 175.160 42.500 175.300 ;
        RECT 42.745 175.300 43.035 175.345 ;
        RECT 42.745 175.160 43.420 175.300 ;
        RECT 41.825 175.115 42.115 175.160 ;
        RECT 42.745 175.115 43.035 175.160 ;
        RECT 42.285 174.960 42.575 175.005 ;
        RECT 40.980 174.820 42.575 174.960 ;
        RECT 43.280 174.960 43.420 175.160 ;
        RECT 46.425 175.115 46.715 175.345 ;
        RECT 47.345 175.300 47.635 175.345 ;
        RECT 48.250 175.300 48.570 175.360 ;
        RECT 48.800 175.345 48.940 175.500 ;
        RECT 50.090 175.440 50.410 175.700 ;
        RECT 66.740 175.685 66.880 175.840 ;
        RECT 73.090 175.780 73.410 175.840 ;
        RECT 73.565 175.795 73.855 176.025 ;
        RECT 74.010 175.980 74.330 176.040 ;
        RECT 90.570 175.980 90.890 176.040 ;
        RECT 74.010 175.840 90.890 175.980 ;
        RECT 51.945 175.640 52.235 175.685 ;
        RECT 51.945 175.500 58.600 175.640 ;
        RECT 51.945 175.455 52.235 175.500 ;
        RECT 47.345 175.160 48.570 175.300 ;
        RECT 47.345 175.115 47.635 175.160 ;
        RECT 48.250 175.100 48.570 175.160 ;
        RECT 48.725 175.115 49.015 175.345 ;
        RECT 49.185 175.115 49.475 175.345 ;
        RECT 50.180 175.300 50.320 175.440 ;
        RECT 58.460 175.360 58.600 175.500 ;
        RECT 66.665 175.455 66.955 175.685 ;
        RECT 51.025 175.300 51.315 175.345 ;
        RECT 50.180 175.160 51.315 175.300 ;
        RECT 51.025 175.115 51.315 175.160 ;
        RECT 52.405 175.300 52.695 175.345 ;
        RECT 52.850 175.300 53.170 175.360 ;
        RECT 52.405 175.160 53.170 175.300 ;
        RECT 52.405 175.115 52.695 175.160 ;
        RECT 45.505 174.960 45.795 175.005 ;
        RECT 43.280 174.820 45.795 174.960 ;
        RECT 36.775 174.775 37.065 174.820 ;
        RECT 39.295 174.775 39.585 174.820 ;
        RECT 40.485 174.775 40.775 174.820 ;
        RECT 42.285 174.775 42.575 174.820 ;
        RECT 45.505 174.775 45.795 174.820 ;
        RECT 47.805 174.775 48.095 175.005 ;
        RECT 37.210 174.620 37.500 174.665 ;
        RECT 38.780 174.620 39.070 174.665 ;
        RECT 40.880 174.620 41.170 174.665 ;
        RECT 37.210 174.480 41.170 174.620 ;
        RECT 37.210 174.435 37.500 174.480 ;
        RECT 38.780 174.435 39.070 174.480 ;
        RECT 40.880 174.435 41.170 174.480 ;
        RECT 46.870 174.420 47.190 174.680 ;
        RECT 47.880 174.620 48.020 174.775 ;
        RECT 48.710 174.620 49.030 174.680 ;
        RECT 47.880 174.480 49.030 174.620 ;
        RECT 48.710 174.420 49.030 174.480 ;
        RECT 49.260 174.340 49.400 175.115 ;
        RECT 52.850 175.100 53.170 175.160 ;
        RECT 53.310 175.100 53.630 175.360 ;
        RECT 58.370 175.100 58.690 175.360 ;
        RECT 70.330 175.300 70.650 175.360 ;
        RECT 71.720 175.300 72.010 175.345 ;
        RECT 70.330 175.160 72.010 175.300 ;
        RECT 70.330 175.100 70.650 175.160 ;
        RECT 71.720 175.115 72.010 175.160 ;
        RECT 72.185 175.300 72.475 175.345 ;
        RECT 73.640 175.300 73.780 175.795 ;
        RECT 74.010 175.780 74.330 175.840 ;
        RECT 90.570 175.780 90.890 175.840 ;
        RECT 76.310 175.640 76.630 175.700 ;
        RECT 75.020 175.500 76.630 175.640 ;
        RECT 75.020 175.345 75.160 175.500 ;
        RECT 76.310 175.440 76.630 175.500 ;
        RECT 78.610 175.640 78.930 175.700 ;
        RECT 79.085 175.640 79.375 175.685 ;
        RECT 78.610 175.500 79.375 175.640 ;
        RECT 78.610 175.440 78.930 175.500 ;
        RECT 79.085 175.455 79.375 175.500 ;
        RECT 81.830 175.640 82.150 175.700 ;
        RECT 83.230 175.640 83.520 175.685 ;
        RECT 84.630 175.640 84.920 175.685 ;
        RECT 86.470 175.640 86.760 175.685 ;
        RECT 81.830 175.500 82.520 175.640 ;
        RECT 81.830 175.440 82.150 175.500 ;
        RECT 72.185 175.160 73.780 175.300 ;
        RECT 72.185 175.115 72.475 175.160 ;
        RECT 74.945 175.115 75.235 175.345 ;
        RECT 75.390 175.300 75.710 175.360 ;
        RECT 77.245 175.300 77.535 175.345 ;
        RECT 75.390 175.160 77.535 175.300 ;
        RECT 75.390 175.100 75.710 175.160 ;
        RECT 77.245 175.115 77.535 175.160 ;
        RECT 78.150 175.100 78.470 175.360 ;
        RECT 82.380 175.345 82.520 175.500 ;
        RECT 83.230 175.500 86.760 175.640 ;
        RECT 83.230 175.455 83.520 175.500 ;
        RECT 84.630 175.455 84.920 175.500 ;
        RECT 86.470 175.455 86.760 175.500 ;
        RECT 82.305 175.115 82.595 175.345 ;
        RECT 83.670 175.100 83.990 175.360 ;
        RECT 85.050 175.100 85.370 175.360 ;
        RECT 50.550 174.760 50.870 175.020 ;
        RECT 68.950 174.960 69.270 175.020 ;
        RECT 70.805 174.960 71.095 175.005 ;
        RECT 68.950 174.820 71.095 174.960 ;
        RECT 68.950 174.760 69.270 174.820 ;
        RECT 70.805 174.775 71.095 174.820 ;
        RECT 71.250 174.760 71.570 175.020 ;
        RECT 73.090 174.760 73.410 175.020 ;
        RECT 74.010 174.960 74.330 175.020 ;
        RECT 85.140 174.960 85.280 175.100 ;
        RECT 74.010 174.820 85.280 174.960 ;
        RECT 74.010 174.760 74.330 174.820 ;
        RECT 50.640 174.620 50.780 174.760 ;
        RECT 51.025 174.620 51.315 174.665 ;
        RECT 50.640 174.480 51.315 174.620 ;
        RECT 71.340 174.620 71.480 174.760 ;
        RECT 73.180 174.620 73.320 174.760 ;
        RECT 71.340 174.480 73.320 174.620 ;
        RECT 82.770 174.620 83.060 174.665 ;
        RECT 85.090 174.620 85.380 174.665 ;
        RECT 86.470 174.620 86.760 174.665 ;
        RECT 82.770 174.480 86.760 174.620 ;
        RECT 51.025 174.435 51.315 174.480 ;
        RECT 82.770 174.435 83.060 174.480 ;
        RECT 85.090 174.435 85.380 174.480 ;
        RECT 86.470 174.435 86.760 174.480 ;
        RECT 34.465 174.280 34.755 174.325 ;
        RECT 44.570 174.280 44.890 174.340 ;
        RECT 49.170 174.280 49.490 174.340 ;
        RECT 34.465 174.140 49.490 174.280 ;
        RECT 34.465 174.095 34.755 174.140 ;
        RECT 44.570 174.080 44.890 174.140 ;
        RECT 49.170 174.080 49.490 174.140 ;
        RECT 60.210 174.080 60.530 174.340 ;
        RECT 73.105 174.280 73.395 174.325 ;
        RECT 74.010 174.280 74.330 174.340 ;
        RECT 73.105 174.140 74.330 174.280 ;
        RECT 73.105 174.095 73.395 174.140 ;
        RECT 74.010 174.080 74.330 174.140 ;
        RECT 74.470 174.080 74.790 174.340 ;
        RECT 90.125 174.280 90.415 174.325 ;
        RECT 90.570 174.280 90.890 174.340 ;
        RECT 90.125 174.140 90.890 174.280 ;
        RECT 90.125 174.095 90.415 174.140 ;
        RECT 90.570 174.080 90.890 174.140 ;
        RECT 18.280 173.460 92.340 173.940 ;
        RECT 46.425 173.260 46.715 173.305 ;
        RECT 46.870 173.260 47.190 173.320 ;
        RECT 46.425 173.120 47.190 173.260 ;
        RECT 46.425 173.075 46.715 173.120 ;
        RECT 46.870 173.060 47.190 173.120 ;
        RECT 48.250 173.260 48.570 173.320 ;
        RECT 52.850 173.260 53.170 173.320 ;
        RECT 48.250 173.120 53.170 173.260 ;
        RECT 48.250 173.060 48.570 173.120 ;
        RECT 52.850 173.060 53.170 173.120 ;
        RECT 53.400 173.120 70.100 173.260 ;
        RECT 48.710 172.920 49.030 172.980 ;
        RECT 51.930 172.920 52.250 172.980 ;
        RECT 53.400 172.920 53.540 173.120 ;
        RECT 69.960 172.980 70.100 173.120 ;
        RECT 74.470 173.060 74.790 173.320 ;
        RECT 75.390 173.060 75.710 173.320 ;
        RECT 76.325 173.260 76.615 173.305 ;
        RECT 79.530 173.260 79.850 173.320 ;
        RECT 76.325 173.120 79.850 173.260 ;
        RECT 76.325 173.075 76.615 173.120 ;
        RECT 48.710 172.780 53.540 172.920 ;
        RECT 48.710 172.720 49.030 172.780 ;
        RECT 51.930 172.720 52.250 172.780 ;
        RECT 62.525 172.735 62.815 172.965 ;
        RECT 65.270 172.920 65.560 172.965 ;
        RECT 66.840 172.920 67.130 172.965 ;
        RECT 68.940 172.920 69.230 172.965 ;
        RECT 65.270 172.780 69.230 172.920 ;
        RECT 65.270 172.735 65.560 172.780 ;
        RECT 66.840 172.735 67.130 172.780 ;
        RECT 68.940 172.735 69.230 172.780 ;
        RECT 69.870 172.920 70.190 172.980 ;
        RECT 72.630 172.920 72.950 172.980 ;
        RECT 69.870 172.780 72.950 172.920 ;
        RECT 54.245 172.580 54.535 172.625 ;
        RECT 58.830 172.580 59.150 172.640 ;
        RECT 62.600 172.580 62.740 172.735 ;
        RECT 69.870 172.720 70.190 172.780 ;
        RECT 72.630 172.720 72.950 172.780 ;
        RECT 44.660 172.440 46.640 172.580 ;
        RECT 44.660 172.300 44.800 172.440 ;
        RECT 38.130 172.040 38.450 172.300 ;
        RECT 44.570 172.040 44.890 172.300 ;
        RECT 46.500 172.285 46.640 172.440 ;
        RECT 54.245 172.440 59.150 172.580 ;
        RECT 54.245 172.395 54.535 172.440 ;
        RECT 58.830 172.380 59.150 172.440 ;
        RECT 59.380 172.440 62.740 172.580 ;
        RECT 45.045 172.055 45.335 172.285 ;
        RECT 46.425 172.055 46.715 172.285 ;
        RECT 47.330 172.240 47.650 172.300 ;
        RECT 51.025 172.240 51.315 172.285 ;
        RECT 47.330 172.100 51.315 172.240 ;
        RECT 45.120 171.620 45.260 172.055 ;
        RECT 47.330 172.040 47.650 172.100 ;
        RECT 51.025 172.055 51.315 172.100 ;
        RECT 51.470 172.240 51.790 172.300 ;
        RECT 51.945 172.240 52.235 172.285 ;
        RECT 52.405 172.240 52.695 172.285 ;
        RECT 51.470 172.100 52.695 172.240 ;
        RECT 51.100 171.900 51.240 172.055 ;
        RECT 51.470 172.040 51.790 172.100 ;
        RECT 51.945 172.055 52.235 172.100 ;
        RECT 52.405 172.055 52.695 172.100 ;
        RECT 53.325 172.055 53.615 172.285 ;
        RECT 56.990 172.240 57.310 172.300 ;
        RECT 58.370 172.285 58.690 172.300 ;
        RECT 57.465 172.240 57.755 172.285 ;
        RECT 56.990 172.100 57.755 172.240 ;
        RECT 53.400 171.900 53.540 172.055 ;
        RECT 56.990 172.040 57.310 172.100 ;
        RECT 57.465 172.055 57.755 172.100 ;
        RECT 58.255 172.240 58.690 172.285 ;
        RECT 59.380 172.240 59.520 172.440 ;
        RECT 58.255 172.100 59.520 172.240 ;
        RECT 58.255 172.055 58.690 172.100 ;
        RECT 59.765 172.055 60.055 172.285 ;
        RECT 58.370 172.040 58.690 172.055 ;
        RECT 51.100 171.760 53.540 171.900 ;
        RECT 54.705 171.715 54.995 171.945 ;
        RECT 55.625 171.900 55.915 171.945 ;
        RECT 58.460 171.900 58.600 172.040 ;
        RECT 55.625 171.760 58.600 171.900 ;
        RECT 55.625 171.715 55.915 171.760 ;
        RECT 41.365 171.560 41.655 171.605 ;
        RECT 42.270 171.560 42.590 171.620 ;
        RECT 41.365 171.420 42.590 171.560 ;
        RECT 41.365 171.375 41.655 171.420 ;
        RECT 42.270 171.360 42.590 171.420 ;
        RECT 45.030 171.360 45.350 171.620 ;
        RECT 45.505 171.560 45.795 171.605 ;
        RECT 45.950 171.560 46.270 171.620 ;
        RECT 45.505 171.420 46.270 171.560 ;
        RECT 45.505 171.375 45.795 171.420 ;
        RECT 45.950 171.360 46.270 171.420 ;
        RECT 51.945 171.560 52.235 171.605 ;
        RECT 52.390 171.560 52.710 171.620 ;
        RECT 51.945 171.420 52.710 171.560 ;
        RECT 51.945 171.375 52.235 171.420 ;
        RECT 52.390 171.360 52.710 171.420 ;
        RECT 52.850 171.560 53.170 171.620 ;
        RECT 54.780 171.560 54.920 171.715 ;
        RECT 58.830 171.700 59.150 171.960 ;
        RECT 59.305 171.715 59.595 171.945 ;
        RECT 59.840 171.900 59.980 172.055 ;
        RECT 61.130 172.040 61.450 172.300 ;
        RECT 62.065 172.240 62.355 172.285 ;
        RECT 62.600 172.240 62.740 172.440 ;
        RECT 64.835 172.580 65.125 172.625 ;
        RECT 67.355 172.580 67.645 172.625 ;
        RECT 68.545 172.580 68.835 172.625 ;
        RECT 76.400 172.580 76.540 173.075 ;
        RECT 79.530 173.060 79.850 173.120 ;
        RECT 81.370 173.260 81.690 173.320 ;
        RECT 81.845 173.260 82.135 173.305 ;
        RECT 81.370 173.120 82.135 173.260 ;
        RECT 81.370 173.060 81.690 173.120 ;
        RECT 81.845 173.075 82.135 173.120 ;
        RECT 64.835 172.440 68.835 172.580 ;
        RECT 64.835 172.395 65.125 172.440 ;
        RECT 67.355 172.395 67.645 172.440 ;
        RECT 68.545 172.395 68.835 172.440 ;
        RECT 73.640 172.440 76.540 172.580 ;
        RECT 78.150 172.580 78.470 172.640 ;
        RECT 79.085 172.580 79.375 172.625 ;
        RECT 90.570 172.580 90.890 172.640 ;
        RECT 78.150 172.440 90.890 172.580 ;
        RECT 62.065 172.100 62.740 172.240 ;
        RECT 62.065 172.055 62.355 172.100 ;
        RECT 69.410 172.040 69.730 172.300 ;
        RECT 73.640 172.285 73.780 172.440 ;
        RECT 78.150 172.380 78.470 172.440 ;
        RECT 79.085 172.395 79.375 172.440 ;
        RECT 90.570 172.380 90.890 172.440 ;
        RECT 73.105 172.055 73.395 172.285 ;
        RECT 73.565 172.055 73.855 172.285 ;
        RECT 74.010 172.240 74.330 172.300 ;
        RECT 84.145 172.240 84.435 172.285 ;
        RECT 74.010 172.100 84.435 172.240 ;
        RECT 61.605 171.900 61.895 171.945 ;
        RECT 59.840 171.760 61.895 171.900 ;
        RECT 61.605 171.715 61.895 171.760 ;
        RECT 63.890 171.900 64.210 171.960 ;
        RECT 68.090 171.900 68.380 171.945 ;
        RECT 63.890 171.760 68.380 171.900 ;
        RECT 52.850 171.420 54.920 171.560 ;
        RECT 56.545 171.560 56.835 171.605 ;
        RECT 59.380 171.560 59.520 171.715 ;
        RECT 63.890 171.700 64.210 171.760 ;
        RECT 68.090 171.715 68.380 171.760 ;
        RECT 56.545 171.420 59.520 171.560 ;
        RECT 52.850 171.360 53.170 171.420 ;
        RECT 56.545 171.375 56.835 171.420 ;
        RECT 60.670 171.360 60.990 171.620 ;
        RECT 72.630 171.560 72.950 171.620 ;
        RECT 73.180 171.560 73.320 172.055 ;
        RECT 74.010 172.040 74.330 172.100 ;
        RECT 84.145 172.055 84.435 172.100 ;
        RECT 85.050 172.240 85.370 172.300 ;
        RECT 85.525 172.240 85.815 172.285 ;
        RECT 85.050 172.100 85.815 172.240 ;
        RECT 85.050 172.040 85.370 172.100 ;
        RECT 85.525 172.055 85.815 172.100 ;
        RECT 86.445 172.240 86.735 172.285 ;
        RECT 87.365 172.240 87.655 172.285 ;
        RECT 86.445 172.100 87.655 172.240 ;
        RECT 86.445 172.055 86.735 172.100 ;
        RECT 87.365 172.055 87.655 172.100 ;
        RECT 90.125 172.240 90.415 172.285 ;
        RECT 91.030 172.240 91.350 172.300 ;
        RECT 90.125 172.100 91.350 172.240 ;
        RECT 90.125 172.055 90.415 172.100 ;
        RECT 74.485 171.900 74.775 171.945 ;
        RECT 77.245 171.900 77.535 171.945 ;
        RECT 80.005 171.900 80.295 171.945 ;
        RECT 90.200 171.900 90.340 172.055 ;
        RECT 91.030 172.040 91.350 172.100 ;
        RECT 74.485 171.760 90.340 171.900 ;
        RECT 74.485 171.715 74.775 171.760 ;
        RECT 77.245 171.715 77.535 171.760 ;
        RECT 80.005 171.715 80.295 171.760 ;
        RECT 76.245 171.560 76.535 171.605 ;
        RECT 78.610 171.560 78.930 171.620 ;
        RECT 72.630 171.420 78.930 171.560 ;
        RECT 72.630 171.360 72.950 171.420 ;
        RECT 76.245 171.375 76.535 171.420 ;
        RECT 78.610 171.360 78.930 171.420 ;
        RECT 79.530 171.560 79.850 171.620 ;
        RECT 80.465 171.560 80.755 171.605 ;
        RECT 79.530 171.420 80.755 171.560 ;
        RECT 79.530 171.360 79.850 171.420 ;
        RECT 80.465 171.375 80.755 171.420 ;
        RECT 80.925 171.560 81.215 171.605 ;
        RECT 81.370 171.560 81.690 171.620 ;
        RECT 80.925 171.420 81.690 171.560 ;
        RECT 80.925 171.375 81.215 171.420 ;
        RECT 81.370 171.360 81.690 171.420 ;
        RECT 83.225 171.560 83.515 171.605 ;
        RECT 83.670 171.560 83.990 171.620 ;
        RECT 83.225 171.420 83.990 171.560 ;
        RECT 83.225 171.375 83.515 171.420 ;
        RECT 83.670 171.360 83.990 171.420 ;
        RECT 18.280 170.740 93.120 171.220 ;
        RECT 33.085 170.540 33.375 170.585 ;
        RECT 38.130 170.540 38.450 170.600 ;
        RECT 50.105 170.540 50.395 170.585 ;
        RECT 53.310 170.540 53.630 170.600 ;
        RECT 33.085 170.400 44.800 170.540 ;
        RECT 33.085 170.355 33.375 170.400 ;
        RECT 38.130 170.340 38.450 170.400 ;
        RECT 38.760 170.200 39.050 170.245 ;
        RECT 41.365 170.200 41.655 170.245 ;
        RECT 42.745 170.200 43.035 170.245 ;
        RECT 38.760 170.060 41.120 170.200 ;
        RECT 38.760 170.015 39.050 170.060 ;
        RECT 40.430 169.660 40.750 169.920 ;
        RECT 35.395 169.520 35.685 169.565 ;
        RECT 37.915 169.520 38.205 169.565 ;
        RECT 39.105 169.520 39.395 169.565 ;
        RECT 35.395 169.380 39.395 169.520 ;
        RECT 35.395 169.335 35.685 169.380 ;
        RECT 37.915 169.335 38.205 169.380 ;
        RECT 39.105 169.335 39.395 169.380 ;
        RECT 39.985 169.335 40.275 169.565 ;
        RECT 40.980 169.520 41.120 170.060 ;
        RECT 41.365 170.060 43.035 170.200 ;
        RECT 41.365 170.015 41.655 170.060 ;
        RECT 42.745 170.015 43.035 170.060 ;
        RECT 41.825 169.675 42.115 169.905 ;
        RECT 40.520 169.380 41.120 169.520 ;
        RECT 41.900 169.520 42.040 169.675 ;
        RECT 42.270 169.660 42.590 169.920 ;
        RECT 43.205 169.860 43.495 169.905 ;
        RECT 44.110 169.860 44.430 169.920 ;
        RECT 43.205 169.720 44.430 169.860 ;
        RECT 44.660 169.860 44.800 170.400 ;
        RECT 50.105 170.400 53.630 170.540 ;
        RECT 50.105 170.355 50.395 170.400 ;
        RECT 45.030 170.200 45.350 170.260 ;
        RECT 45.030 170.060 48.020 170.200 ;
        RECT 45.030 170.000 45.350 170.060 ;
        RECT 45.580 169.905 45.720 170.060 ;
        RECT 47.880 169.920 48.020 170.060 ;
        RECT 49.170 170.000 49.490 170.260 ;
        RECT 44.660 169.720 45.260 169.860 ;
        RECT 43.205 169.675 43.495 169.720 ;
        RECT 44.110 169.660 44.430 169.720 ;
        RECT 44.585 169.520 44.875 169.565 ;
        RECT 41.900 169.380 44.875 169.520 ;
        RECT 45.120 169.520 45.260 169.720 ;
        RECT 45.505 169.675 45.795 169.905 ;
        RECT 45.950 169.860 46.270 169.920 ;
        RECT 45.950 169.720 46.640 169.860 ;
        RECT 45.950 169.660 46.270 169.720 ;
        RECT 46.500 169.520 46.640 169.720 ;
        RECT 46.885 169.675 47.175 169.905 ;
        RECT 45.120 169.380 46.640 169.520 ;
        RECT 46.960 169.520 47.100 169.675 ;
        RECT 47.330 169.660 47.650 169.920 ;
        RECT 47.790 169.660 48.110 169.920 ;
        RECT 48.725 169.860 49.015 169.905 ;
        RECT 50.180 169.860 50.320 170.355 ;
        RECT 53.310 170.340 53.630 170.400 ;
        RECT 57.450 170.340 57.770 170.600 ;
        RECT 60.670 170.340 60.990 170.600 ;
        RECT 63.890 170.340 64.210 170.600 ;
        RECT 73.180 170.400 77.000 170.540 ;
        RECT 50.550 170.200 50.870 170.260 ;
        RECT 57.540 170.200 57.680 170.340 ;
        RECT 50.550 170.060 57.680 170.200 ;
        RECT 50.550 170.000 50.870 170.060 ;
        RECT 48.725 169.720 50.320 169.860 ;
        RECT 51.025 169.860 51.315 169.905 ;
        RECT 59.750 169.860 60.070 169.920 ;
        RECT 51.025 169.720 60.070 169.860 ;
        RECT 60.760 169.860 60.900 170.340 ;
        RECT 71.710 170.200 72.030 170.260 ;
        RECT 73.180 170.200 73.320 170.400 ;
        RECT 67.660 170.060 73.320 170.200 ;
        RECT 67.660 169.920 67.800 170.060 ;
        RECT 71.710 170.000 72.030 170.060 ;
        RECT 61.605 169.860 61.895 169.905 ;
        RECT 60.760 169.720 61.895 169.860 ;
        RECT 48.725 169.675 49.015 169.720 ;
        RECT 51.025 169.675 51.315 169.720 ;
        RECT 48.265 169.520 48.555 169.565 ;
        RECT 46.960 169.380 48.555 169.520 ;
        RECT 35.830 169.180 36.120 169.225 ;
        RECT 37.400 169.180 37.690 169.225 ;
        RECT 39.500 169.180 39.790 169.225 ;
        RECT 35.830 169.040 39.790 169.180 ;
        RECT 35.830 168.995 36.120 169.040 ;
        RECT 37.400 168.995 37.690 169.040 ;
        RECT 39.500 168.995 39.790 169.040 ;
        RECT 38.130 168.840 38.450 168.900 ;
        RECT 40.060 168.840 40.200 169.335 ;
        RECT 40.520 169.225 40.660 169.380 ;
        RECT 44.585 169.335 44.875 169.380 ;
        RECT 40.445 168.995 40.735 169.225 ;
        RECT 44.110 168.980 44.430 169.240 ;
        RECT 46.500 169.180 46.640 169.380 ;
        RECT 48.265 169.335 48.555 169.380 ;
        RECT 48.800 169.180 48.940 169.675 ;
        RECT 59.750 169.660 60.070 169.720 ;
        RECT 61.605 169.675 61.895 169.720 ;
        RECT 62.525 169.860 62.815 169.905 ;
        RECT 62.985 169.860 63.275 169.905 ;
        RECT 62.525 169.720 63.275 169.860 ;
        RECT 62.525 169.675 62.815 169.720 ;
        RECT 62.985 169.675 63.275 169.720 ;
        RECT 67.570 169.660 67.890 169.920 ;
        RECT 72.630 169.660 72.950 169.920 ;
        RECT 73.180 169.860 73.320 170.060 ;
        RECT 73.565 170.200 73.855 170.245 ;
        RECT 76.325 170.200 76.615 170.245 ;
        RECT 73.565 170.060 76.615 170.200 ;
        RECT 73.565 170.015 73.855 170.060 ;
        RECT 76.325 170.015 76.615 170.060 ;
        RECT 76.860 169.920 77.000 170.400 ;
        RECT 83.230 170.200 83.520 170.245 ;
        RECT 84.630 170.200 84.920 170.245 ;
        RECT 86.470 170.200 86.760 170.245 ;
        RECT 83.230 170.060 86.760 170.200 ;
        RECT 83.230 170.015 83.520 170.060 ;
        RECT 84.630 170.015 84.920 170.060 ;
        RECT 86.470 170.015 86.760 170.060 ;
        RECT 74.025 169.860 74.315 169.905 ;
        RECT 73.180 169.720 74.315 169.860 ;
        RECT 74.025 169.675 74.315 169.720 ;
        RECT 74.485 169.675 74.775 169.905 ;
        RECT 75.865 169.675 76.155 169.905 ;
        RECT 60.670 169.520 60.990 169.580 ;
        RECT 62.050 169.520 62.370 169.580 ;
        RECT 60.670 169.380 62.370 169.520 ;
        RECT 60.670 169.320 60.990 169.380 ;
        RECT 62.050 169.320 62.370 169.380 ;
        RECT 72.170 169.520 72.490 169.580 ;
        RECT 74.560 169.520 74.700 169.675 ;
        RECT 72.170 169.380 74.700 169.520 ;
        RECT 75.940 169.520 76.080 169.675 ;
        RECT 76.770 169.660 77.090 169.920 ;
        RECT 79.530 169.660 79.850 169.920 ;
        RECT 83.670 169.660 83.990 169.920 ;
        RECT 79.620 169.520 79.760 169.660 ;
        RECT 75.940 169.380 79.760 169.520 ;
        RECT 81.830 169.520 82.150 169.580 ;
        RECT 82.305 169.520 82.595 169.565 ;
        RECT 81.830 169.380 82.595 169.520 ;
        RECT 72.170 169.320 72.490 169.380 ;
        RECT 81.830 169.320 82.150 169.380 ;
        RECT 82.305 169.335 82.595 169.380 ;
        RECT 62.510 169.180 62.830 169.240 ;
        RECT 46.500 169.040 48.940 169.180 ;
        RECT 51.560 169.040 62.830 169.180 ;
        RECT 38.130 168.700 40.200 168.840 ;
        RECT 44.200 168.840 44.340 168.980 ;
        RECT 51.560 168.840 51.700 169.040 ;
        RECT 62.510 168.980 62.830 169.040 ;
        RECT 82.770 169.180 83.060 169.225 ;
        RECT 85.090 169.180 85.380 169.225 ;
        RECT 86.470 169.180 86.760 169.225 ;
        RECT 82.770 169.040 86.760 169.180 ;
        RECT 82.770 168.995 83.060 169.040 ;
        RECT 85.090 168.995 85.380 169.040 ;
        RECT 86.470 168.995 86.760 169.040 ;
        RECT 44.200 168.700 51.700 168.840 ;
        RECT 38.130 168.640 38.450 168.700 ;
        RECT 51.930 168.640 52.250 168.900 ;
        RECT 75.405 168.840 75.695 168.885 ;
        RECT 76.310 168.840 76.630 168.900 ;
        RECT 75.405 168.700 76.630 168.840 ;
        RECT 75.405 168.655 75.695 168.700 ;
        RECT 76.310 168.640 76.630 168.700 ;
        RECT 90.125 168.840 90.415 168.885 ;
        RECT 91.030 168.840 91.350 168.900 ;
        RECT 90.125 168.700 91.350 168.840 ;
        RECT 90.125 168.655 90.415 168.700 ;
        RECT 91.030 168.640 91.350 168.700 ;
        RECT 18.280 168.020 92.340 168.500 ;
        RECT 55.165 167.820 55.455 167.865 ;
        RECT 61.130 167.820 61.450 167.880 ;
        RECT 55.165 167.680 61.450 167.820 ;
        RECT 55.165 167.635 55.455 167.680 ;
        RECT 61.130 167.620 61.450 167.680 ;
        RECT 77.705 167.480 77.995 167.525 ;
        RECT 80.910 167.480 81.230 167.540 ;
        RECT 77.705 167.340 81.230 167.480 ;
        RECT 77.705 167.295 77.995 167.340 ;
        RECT 80.910 167.280 81.230 167.340 ;
        RECT 51.930 167.140 52.250 167.200 ;
        RECT 56.990 167.140 57.310 167.200 ;
        RECT 60.685 167.140 60.975 167.185 ;
        RECT 67.570 167.140 67.890 167.200 ;
        RECT 51.930 167.000 54.460 167.140 ;
        RECT 51.930 166.940 52.250 167.000 ;
        RECT 53.770 166.600 54.090 166.860 ;
        RECT 54.320 166.845 54.460 167.000 ;
        RECT 56.990 167.000 67.890 167.140 ;
        RECT 56.990 166.940 57.310 167.000 ;
        RECT 60.685 166.955 60.975 167.000 ;
        RECT 67.570 166.940 67.890 167.000 ;
        RECT 68.030 167.140 68.350 167.200 ;
        RECT 78.610 167.140 78.930 167.200 ;
        RECT 68.030 167.000 76.540 167.140 ;
        RECT 68.030 166.940 68.350 167.000 ;
        RECT 54.245 166.615 54.535 166.845 ;
        RECT 56.530 166.800 56.850 166.860 ;
        RECT 59.750 166.845 60.070 166.860 ;
        RECT 58.385 166.800 58.675 166.845 ;
        RECT 56.530 166.660 58.675 166.800 ;
        RECT 56.530 166.600 56.850 166.660 ;
        RECT 58.385 166.615 58.675 166.660 ;
        RECT 59.750 166.615 60.185 166.845 ;
        RECT 75.405 166.800 75.695 166.845 ;
        RECT 75.850 166.800 76.170 166.860 ;
        RECT 76.400 166.845 76.540 167.000 ;
        RECT 78.610 167.000 81.600 167.140 ;
        RECT 78.610 166.940 78.930 167.000 ;
        RECT 75.405 166.660 76.170 166.800 ;
        RECT 75.405 166.615 75.695 166.660 ;
        RECT 59.750 166.600 60.070 166.615 ;
        RECT 75.850 166.600 76.170 166.660 ;
        RECT 76.325 166.615 76.615 166.845 ;
        RECT 76.770 166.600 77.090 166.860 ;
        RECT 78.195 166.800 78.485 166.845 ;
        RECT 78.700 166.800 78.840 166.940 ;
        RECT 81.460 166.860 81.600 167.000 ;
        RECT 78.195 166.660 78.840 166.800 ;
        RECT 78.195 166.615 78.485 166.660 ;
        RECT 79.085 166.615 79.375 166.845 ;
        RECT 81.370 166.800 81.690 166.860 ;
        RECT 90.110 166.800 90.430 166.860 ;
        RECT 81.370 166.660 90.430 166.800 ;
        RECT 56.990 166.460 57.310 166.520 ;
        RECT 58.845 166.460 59.135 166.505 ;
        RECT 56.990 166.320 59.135 166.460 ;
        RECT 56.990 166.260 57.310 166.320 ;
        RECT 58.845 166.275 59.135 166.320 ;
        RECT 59.290 166.460 59.610 166.520 ;
        RECT 61.605 166.460 61.895 166.505 ;
        RECT 59.290 166.320 61.895 166.460 ;
        RECT 59.290 166.260 59.610 166.320 ;
        RECT 61.605 166.275 61.895 166.320 ;
        RECT 63.445 166.460 63.735 166.505 ;
        RECT 66.650 166.460 66.970 166.520 ;
        RECT 63.445 166.320 66.970 166.460 ;
        RECT 63.445 166.275 63.735 166.320 ;
        RECT 66.650 166.260 66.970 166.320 ;
        RECT 46.870 166.120 47.190 166.180 ;
        RECT 48.710 166.120 49.030 166.180 ;
        RECT 46.870 165.980 49.030 166.120 ;
        RECT 46.870 165.920 47.190 165.980 ;
        RECT 48.710 165.920 49.030 165.980 ;
        RECT 57.450 165.920 57.770 166.180 ;
        RECT 68.030 166.120 68.350 166.180 ;
        RECT 72.185 166.120 72.475 166.165 ;
        RECT 68.030 165.980 72.475 166.120 ;
        RECT 76.860 166.120 77.000 166.600 ;
        RECT 77.705 166.460 77.995 166.505 ;
        RECT 78.610 166.460 78.930 166.520 ;
        RECT 77.705 166.320 78.930 166.460 ;
        RECT 77.705 166.275 77.995 166.320 ;
        RECT 78.610 166.260 78.930 166.320 ;
        RECT 79.160 166.120 79.300 166.615 ;
        RECT 81.370 166.600 81.690 166.660 ;
        RECT 90.110 166.600 90.430 166.660 ;
        RECT 76.860 165.980 79.300 166.120 ;
        RECT 68.030 165.920 68.350 165.980 ;
        RECT 72.185 165.935 72.475 165.980 ;
        RECT 18.280 165.300 93.120 165.780 ;
        RECT 47.790 165.100 48.110 165.160 ;
        RECT 48.265 165.100 48.555 165.145 ;
        RECT 47.790 164.960 48.555 165.100 ;
        RECT 47.790 164.900 48.110 164.960 ;
        RECT 48.265 164.915 48.555 164.960 ;
        RECT 49.105 165.100 49.395 165.145 ;
        RECT 53.770 165.100 54.090 165.160 ;
        RECT 49.105 164.960 54.090 165.100 ;
        RECT 49.105 164.915 49.395 164.960 ;
        RECT 48.340 164.760 48.480 164.915 ;
        RECT 53.770 164.900 54.090 164.960 ;
        RECT 56.085 165.100 56.375 165.145 ;
        RECT 56.990 165.100 57.310 165.160 ;
        RECT 56.085 164.960 57.310 165.100 ;
        RECT 56.085 164.915 56.375 164.960 ;
        RECT 56.990 164.900 57.310 164.960 ;
        RECT 57.450 164.900 57.770 165.160 ;
        RECT 58.845 165.100 59.135 165.145 ;
        RECT 59.750 165.100 60.070 165.160 ;
        RECT 58.845 164.960 60.070 165.100 ;
        RECT 58.845 164.915 59.135 164.960 ;
        RECT 46.500 164.620 48.480 164.760 ;
        RECT 50.105 164.760 50.395 164.805 ;
        RECT 50.550 164.760 50.870 164.820 ;
        RECT 53.325 164.760 53.615 164.805 ;
        RECT 56.530 164.760 56.850 164.820 ;
        RECT 50.105 164.620 50.870 164.760 ;
        RECT 38.605 164.235 38.895 164.465 ;
        RECT 39.525 164.420 39.815 164.465 ;
        RECT 42.730 164.420 43.050 164.480 ;
        RECT 46.500 164.465 46.640 164.620 ;
        RECT 50.105 164.575 50.395 164.620 ;
        RECT 50.550 164.560 50.870 164.620 ;
        RECT 51.560 164.620 56.850 164.760 ;
        RECT 39.525 164.280 43.050 164.420 ;
        RECT 39.525 164.235 39.815 164.280 ;
        RECT 38.680 164.080 38.820 164.235 ;
        RECT 42.730 164.220 43.050 164.280 ;
        RECT 45.505 164.235 45.795 164.465 ;
        RECT 46.425 164.235 46.715 164.465 ;
        RECT 44.585 164.080 44.875 164.125 ;
        RECT 38.680 163.940 44.875 164.080 ;
        RECT 45.580 164.080 45.720 164.235 ;
        RECT 46.870 164.220 47.190 164.480 ;
        RECT 47.790 164.420 48.110 164.480 ;
        RECT 51.560 164.465 51.700 164.620 ;
        RECT 53.325 164.575 53.615 164.620 ;
        RECT 56.530 164.560 56.850 164.620 ;
        RECT 47.790 164.410 48.480 164.420 ;
        RECT 47.790 164.280 48.940 164.410 ;
        RECT 47.790 164.220 48.110 164.280 ;
        RECT 48.340 164.270 48.940 164.280 ;
        RECT 47.330 164.080 47.650 164.140 ;
        RECT 45.580 163.940 47.650 164.080 ;
        RECT 48.800 164.080 48.940 164.270 ;
        RECT 51.485 164.235 51.775 164.465 ;
        RECT 52.865 164.235 53.155 164.465 ;
        RECT 53.770 164.420 54.090 164.480 ;
        RECT 57.540 164.465 57.680 164.900 ;
        RECT 54.245 164.420 54.535 164.465 ;
        RECT 53.770 164.280 54.535 164.420 ;
        RECT 52.405 164.080 52.695 164.125 ;
        RECT 48.800 163.940 52.695 164.080 ;
        RECT 44.585 163.895 44.875 163.940 ;
        RECT 47.330 163.880 47.650 163.940 ;
        RECT 52.405 163.895 52.695 163.940 ;
        RECT 52.940 164.080 53.080 164.235 ;
        RECT 53.770 164.220 54.090 164.280 ;
        RECT 54.245 164.235 54.535 164.280 ;
        RECT 55.165 164.420 55.455 164.465 ;
        RECT 55.165 164.280 57.220 164.420 ;
        RECT 55.165 164.235 55.455 164.280 ;
        RECT 55.240 164.080 55.380 164.235 ;
        RECT 52.940 163.940 55.380 164.080 ;
        RECT 45.965 163.740 46.255 163.785 ;
        RECT 50.565 163.740 50.855 163.785 ;
        RECT 45.965 163.600 47.560 163.740 ;
        RECT 45.965 163.555 46.255 163.600 ;
        RECT 37.670 163.400 37.990 163.460 ;
        RECT 38.605 163.400 38.895 163.445 ;
        RECT 37.670 163.260 38.895 163.400 ;
        RECT 47.420 163.400 47.560 163.600 ;
        RECT 48.340 163.600 50.855 163.740 ;
        RECT 48.340 163.400 48.480 163.600 ;
        RECT 50.565 163.555 50.855 163.600 ;
        RECT 47.420 163.260 48.480 163.400 ;
        RECT 49.185 163.400 49.475 163.445 ;
        RECT 52.940 163.400 53.080 163.940 ;
        RECT 56.545 163.895 56.835 164.125 ;
        RECT 57.080 164.080 57.220 164.280 ;
        RECT 57.465 164.235 57.755 164.465 ;
        RECT 58.920 164.080 59.060 164.915 ;
        RECT 59.750 164.900 60.070 164.960 ;
        RECT 69.425 165.100 69.715 165.145 ;
        RECT 74.010 165.100 74.330 165.160 ;
        RECT 75.850 165.100 76.170 165.160 ;
        RECT 77.245 165.100 77.535 165.145 ;
        RECT 85.050 165.100 85.370 165.160 ;
        RECT 69.425 164.960 70.560 165.100 ;
        RECT 69.425 164.915 69.715 164.960 ;
        RECT 70.420 164.760 70.560 164.960 ;
        RECT 74.010 164.960 77.535 165.100 ;
        RECT 74.010 164.900 74.330 164.960 ;
        RECT 75.850 164.900 76.170 164.960 ;
        RECT 77.245 164.915 77.535 164.960 ;
        RECT 80.540 164.960 85.370 165.100 ;
        RECT 71.570 164.760 71.860 164.805 ;
        RECT 65.820 164.620 69.640 164.760 ;
        RECT 70.420 164.620 71.860 164.760 ;
        RECT 62.970 164.420 63.290 164.480 ;
        RECT 65.820 164.465 65.960 164.620 ;
        RECT 69.500 164.480 69.640 164.620 ;
        RECT 71.570 164.575 71.860 164.620 ;
        RECT 77.690 164.760 78.010 164.820 ;
        RECT 77.690 164.620 79.300 164.760 ;
        RECT 77.690 164.560 78.010 164.620 ;
        RECT 64.410 164.420 64.700 164.465 ;
        RECT 62.970 164.280 64.700 164.420 ;
        RECT 62.970 164.220 63.290 164.280 ;
        RECT 64.410 164.235 64.700 164.280 ;
        RECT 65.745 164.235 66.035 164.465 ;
        RECT 66.650 164.220 66.970 164.480 ;
        RECT 67.125 164.420 67.415 164.465 ;
        RECT 68.030 164.420 68.350 164.480 ;
        RECT 67.125 164.280 68.350 164.420 ;
        RECT 67.125 164.235 67.415 164.280 ;
        RECT 68.030 164.220 68.350 164.280 ;
        RECT 68.490 164.220 68.810 164.480 ;
        RECT 69.410 164.420 69.730 164.480 ;
        RECT 70.345 164.420 70.635 164.465 ;
        RECT 78.240 164.420 78.380 164.620 ;
        RECT 69.410 164.280 70.635 164.420 ;
        RECT 69.410 164.220 69.730 164.280 ;
        RECT 70.345 164.235 70.635 164.280 ;
        RECT 70.880 164.280 78.380 164.420 ;
        RECT 57.080 163.940 59.060 164.080 ;
        RECT 61.155 164.080 61.445 164.125 ;
        RECT 63.675 164.080 63.965 164.125 ;
        RECT 64.865 164.080 65.155 164.125 ;
        RECT 61.155 163.940 65.155 164.080 ;
        RECT 66.740 164.080 66.880 164.220 ;
        RECT 67.585 164.080 67.875 164.125 ;
        RECT 70.880 164.080 71.020 164.280 ;
        RECT 78.610 164.220 78.930 164.480 ;
        RECT 79.160 164.465 79.300 164.620 ;
        RECT 80.540 164.465 80.680 164.960 ;
        RECT 85.050 164.900 85.370 164.960 ;
        RECT 81.830 164.560 82.150 164.820 ;
        RECT 83.230 164.760 83.520 164.805 ;
        RECT 84.630 164.760 84.920 164.805 ;
        RECT 86.470 164.760 86.760 164.805 ;
        RECT 83.230 164.620 86.760 164.760 ;
        RECT 83.230 164.575 83.520 164.620 ;
        RECT 84.630 164.575 84.920 164.620 ;
        RECT 86.470 164.575 86.760 164.620 ;
        RECT 79.085 164.235 79.375 164.465 ;
        RECT 80.465 164.235 80.755 164.465 ;
        RECT 80.910 164.220 81.230 164.480 ;
        RECT 81.920 164.420 82.060 164.560 ;
        RECT 82.305 164.420 82.595 164.465 ;
        RECT 85.970 164.420 86.290 164.480 ;
        RECT 81.920 164.280 82.595 164.420 ;
        RECT 82.305 164.235 82.595 164.280 ;
        RECT 83.300 164.280 86.290 164.420 ;
        RECT 66.740 163.940 71.020 164.080 ;
        RECT 71.225 164.080 71.515 164.125 ;
        RECT 72.415 164.080 72.705 164.125 ;
        RECT 74.935 164.080 75.225 164.125 ;
        RECT 71.225 163.940 75.225 164.080 ;
        RECT 61.155 163.895 61.445 163.940 ;
        RECT 63.675 163.895 63.965 163.940 ;
        RECT 64.865 163.895 65.155 163.940 ;
        RECT 67.585 163.895 67.875 163.940 ;
        RECT 71.225 163.895 71.515 163.940 ;
        RECT 72.415 163.895 72.705 163.940 ;
        RECT 74.935 163.895 75.225 163.940 ;
        RECT 77.705 163.895 77.995 164.125 ;
        RECT 81.845 164.080 82.135 164.125 ;
        RECT 83.300 164.080 83.440 164.280 ;
        RECT 85.970 164.220 86.290 164.280 ;
        RECT 81.845 163.940 83.440 164.080 ;
        RECT 83.685 164.080 83.975 164.125 ;
        RECT 84.130 164.080 84.450 164.140 ;
        RECT 83.685 163.940 84.450 164.080 ;
        RECT 81.845 163.895 82.135 163.940 ;
        RECT 83.685 163.895 83.975 163.940 ;
        RECT 56.620 163.740 56.760 163.895 ;
        RECT 60.670 163.740 60.990 163.800 ;
        RECT 56.620 163.600 60.990 163.740 ;
        RECT 60.670 163.540 60.990 163.600 ;
        RECT 61.590 163.740 61.880 163.785 ;
        RECT 63.160 163.740 63.450 163.785 ;
        RECT 65.260 163.740 65.550 163.785 ;
        RECT 61.590 163.600 65.550 163.740 ;
        RECT 61.590 163.555 61.880 163.600 ;
        RECT 63.160 163.555 63.450 163.600 ;
        RECT 65.260 163.555 65.550 163.600 ;
        RECT 70.830 163.740 71.120 163.785 ;
        RECT 72.930 163.740 73.220 163.785 ;
        RECT 74.500 163.740 74.790 163.785 ;
        RECT 70.830 163.600 74.790 163.740 ;
        RECT 77.780 163.740 77.920 163.895 ;
        RECT 84.130 163.880 84.450 163.940 ;
        RECT 79.530 163.740 79.850 163.800 ;
        RECT 82.770 163.740 83.060 163.785 ;
        RECT 85.090 163.740 85.380 163.785 ;
        RECT 86.470 163.740 86.760 163.785 ;
        RECT 77.780 163.600 82.060 163.740 ;
        RECT 70.830 163.555 71.120 163.600 ;
        RECT 72.930 163.555 73.220 163.600 ;
        RECT 74.500 163.555 74.790 163.600 ;
        RECT 79.530 163.540 79.850 163.600 ;
        RECT 49.185 163.260 53.080 163.400 ;
        RECT 37.670 163.200 37.990 163.260 ;
        RECT 38.605 163.215 38.895 163.260 ;
        RECT 49.185 163.215 49.475 163.260 ;
        RECT 58.370 163.200 58.690 163.460 ;
        RECT 78.150 163.200 78.470 163.460 ;
        RECT 81.370 163.200 81.690 163.460 ;
        RECT 81.920 163.400 82.060 163.600 ;
        RECT 82.770 163.600 86.760 163.740 ;
        RECT 82.770 163.555 83.060 163.600 ;
        RECT 85.090 163.555 85.380 163.600 ;
        RECT 86.470 163.555 86.760 163.600 ;
        RECT 87.810 163.540 88.130 163.800 ;
        RECT 87.900 163.400 88.040 163.540 ;
        RECT 81.920 163.260 88.040 163.400 ;
        RECT 90.125 163.400 90.415 163.445 ;
        RECT 90.570 163.400 90.890 163.460 ;
        RECT 90.125 163.260 90.890 163.400 ;
        RECT 90.125 163.215 90.415 163.260 ;
        RECT 90.570 163.200 90.890 163.260 ;
        RECT 18.280 162.580 92.340 163.060 ;
        RECT 47.345 162.380 47.635 162.425 ;
        RECT 47.790 162.380 48.110 162.440 ;
        RECT 47.345 162.240 48.110 162.380 ;
        RECT 47.345 162.195 47.635 162.240 ;
        RECT 47.790 162.180 48.110 162.240 ;
        RECT 52.405 162.380 52.695 162.425 ;
        RECT 61.145 162.380 61.435 162.425 ;
        RECT 62.970 162.380 63.290 162.440 ;
        RECT 52.405 162.240 53.540 162.380 ;
        RECT 52.405 162.195 52.695 162.240 ;
        RECT 53.400 162.100 53.540 162.240 ;
        RECT 61.145 162.240 63.290 162.380 ;
        RECT 61.145 162.195 61.435 162.240 ;
        RECT 62.970 162.180 63.290 162.240 ;
        RECT 68.490 162.180 68.810 162.440 ;
        RECT 76.785 162.195 77.075 162.425 ;
        RECT 83.225 162.380 83.515 162.425 ;
        RECT 84.130 162.380 84.450 162.440 ;
        RECT 83.225 162.240 84.450 162.380 ;
        RECT 83.225 162.195 83.515 162.240 ;
        RECT 36.790 162.040 37.080 162.085 ;
        RECT 38.890 162.040 39.180 162.085 ;
        RECT 40.460 162.040 40.750 162.085 ;
        RECT 36.790 161.900 40.750 162.040 ;
        RECT 36.790 161.855 37.080 161.900 ;
        RECT 38.890 161.855 39.180 161.900 ;
        RECT 40.460 161.855 40.750 161.900 ;
        RECT 43.205 162.040 43.495 162.085 ;
        RECT 51.485 162.040 51.775 162.085 ;
        RECT 52.850 162.040 53.170 162.100 ;
        RECT 43.205 161.900 47.100 162.040 ;
        RECT 43.205 161.855 43.495 161.900 ;
        RECT 37.185 161.700 37.475 161.745 ;
        RECT 38.375 161.700 38.665 161.745 ;
        RECT 40.895 161.700 41.185 161.745 ;
        RECT 37.185 161.560 41.185 161.700 ;
        RECT 37.185 161.515 37.475 161.560 ;
        RECT 38.375 161.515 38.665 161.560 ;
        RECT 40.895 161.515 41.185 161.560 ;
        RECT 46.960 161.405 47.100 161.900 ;
        RECT 51.485 161.900 53.170 162.040 ;
        RECT 51.485 161.855 51.775 161.900 ;
        RECT 52.850 161.840 53.170 161.900 ;
        RECT 53.310 162.040 53.630 162.100 ;
        RECT 76.860 162.040 77.000 162.195 ;
        RECT 84.130 162.180 84.450 162.240 ;
        RECT 79.085 162.040 79.375 162.085 ;
        RECT 80.450 162.040 80.770 162.100 ;
        RECT 53.310 161.900 54.460 162.040 ;
        RECT 76.860 161.900 77.920 162.040 ;
        RECT 53.310 161.840 53.630 161.900 ;
        RECT 51.560 161.560 53.080 161.700 ;
        RECT 36.305 161.360 36.595 161.405 ;
        RECT 46.885 161.360 47.175 161.405 ;
        RECT 50.550 161.360 50.870 161.420 ;
        RECT 36.305 161.220 38.360 161.360 ;
        RECT 36.305 161.175 36.595 161.220 ;
        RECT 37.670 161.065 37.990 161.080 ;
        RECT 37.640 161.020 37.990 161.065 ;
        RECT 37.475 160.880 37.990 161.020 ;
        RECT 37.640 160.835 37.990 160.880 ;
        RECT 37.670 160.820 37.990 160.835 ;
        RECT 38.220 160.740 38.360 161.220 ;
        RECT 46.885 161.220 50.870 161.360 ;
        RECT 46.885 161.175 47.175 161.220 ;
        RECT 50.550 161.160 50.870 161.220 ;
        RECT 50.090 161.020 50.410 161.080 ;
        RECT 51.560 161.020 51.700 161.560 ;
        RECT 50.090 160.880 51.700 161.020 ;
        RECT 52.175 161.020 52.465 161.235 ;
        RECT 52.940 161.020 53.080 161.560 ;
        RECT 53.785 161.370 54.075 161.405 ;
        RECT 54.320 161.370 54.460 161.900 ;
        RECT 59.305 161.700 59.595 161.745 ;
        RECT 74.930 161.700 75.250 161.760 ;
        RECT 59.305 161.560 75.250 161.700 ;
        RECT 59.305 161.515 59.595 161.560 ;
        RECT 74.930 161.500 75.250 161.560 ;
        RECT 53.785 161.230 54.460 161.370 ;
        RECT 53.785 161.175 54.075 161.230 ;
        RECT 54.705 161.175 54.995 161.405 ;
        RECT 58.370 161.360 58.690 161.420 ;
        RECT 76.310 161.405 76.630 161.420 ;
        RECT 77.780 161.405 77.920 161.900 ;
        RECT 79.085 161.900 80.770 162.040 ;
        RECT 79.085 161.855 79.375 161.900 ;
        RECT 80.450 161.840 80.770 161.900 ;
        RECT 60.225 161.360 60.515 161.405 ;
        RECT 58.370 161.220 60.515 161.360 ;
        RECT 53.325 161.020 53.615 161.065 ;
        RECT 54.780 161.020 54.920 161.175 ;
        RECT 58.370 161.160 58.690 161.220 ;
        RECT 60.225 161.175 60.515 161.220 ;
        RECT 69.885 161.175 70.175 161.405 ;
        RECT 76.275 161.360 76.630 161.405 ;
        RECT 76.115 161.220 76.630 161.360 ;
        RECT 76.275 161.175 76.630 161.220 ;
        RECT 77.245 161.175 77.535 161.405 ;
        RECT 77.705 161.175 77.995 161.405 ;
        RECT 52.175 161.005 52.620 161.020 ;
        RECT 52.320 160.880 52.620 161.005 ;
        RECT 52.940 160.880 54.920 161.020 ;
        RECT 56.530 161.020 56.850 161.080 ;
        RECT 57.925 161.020 58.215 161.065 ;
        RECT 56.530 160.880 58.215 161.020 ;
        RECT 50.090 160.820 50.410 160.880 ;
        RECT 38.130 160.480 38.450 160.740 ;
        RECT 51.930 160.680 52.250 160.740 ;
        RECT 52.480 160.680 52.620 160.880 ;
        RECT 53.325 160.835 53.615 160.880 ;
        RECT 56.530 160.820 56.850 160.880 ;
        RECT 57.925 160.835 58.215 160.880 ;
        RECT 68.030 161.020 68.350 161.080 ;
        RECT 68.505 161.020 68.795 161.065 ;
        RECT 68.950 161.020 69.270 161.080 ;
        RECT 68.030 160.880 69.270 161.020 ;
        RECT 69.960 161.020 70.100 161.175 ;
        RECT 76.310 161.160 76.630 161.175 ;
        RECT 72.170 161.020 72.490 161.080 ;
        RECT 74.010 161.020 74.330 161.080 ;
        RECT 69.960 160.880 74.330 161.020 ;
        RECT 68.030 160.820 68.350 160.880 ;
        RECT 68.505 160.835 68.795 160.880 ;
        RECT 68.950 160.820 69.270 160.880 ;
        RECT 72.170 160.820 72.490 160.880 ;
        RECT 74.010 160.820 74.330 160.880 ;
        RECT 51.930 160.540 52.620 160.680 ;
        RECT 51.930 160.480 52.250 160.540 ;
        RECT 54.230 160.480 54.550 160.740 ;
        RECT 69.425 160.680 69.715 160.725 ;
        RECT 69.870 160.680 70.190 160.740 ;
        RECT 69.425 160.540 70.190 160.680 ;
        RECT 69.425 160.495 69.715 160.540 ;
        RECT 69.870 160.480 70.190 160.540 ;
        RECT 74.930 160.680 75.250 160.740 ;
        RECT 77.320 160.680 77.460 161.175 ;
        RECT 78.150 161.160 78.470 161.420 ;
        RECT 79.085 161.360 79.375 161.405 ;
        RECT 79.990 161.360 80.310 161.420 ;
        RECT 79.085 161.220 80.310 161.360 ;
        RECT 79.085 161.175 79.375 161.220 ;
        RECT 79.990 161.160 80.310 161.220 ;
        RECT 80.910 161.160 81.230 161.420 ;
        RECT 81.370 161.360 81.690 161.420 ;
        RECT 83.225 161.360 83.515 161.405 ;
        RECT 81.370 161.220 83.515 161.360 ;
        RECT 81.370 161.160 81.690 161.220 ;
        RECT 83.225 161.175 83.515 161.220 ;
        RECT 84.605 161.175 84.895 161.405 ;
        RECT 81.000 161.020 81.140 161.160 ;
        RECT 84.680 161.020 84.820 161.175 ;
        RECT 85.050 161.160 85.370 161.420 ;
        RECT 81.000 160.880 84.820 161.020 ;
        RECT 84.145 160.680 84.435 160.725 ;
        RECT 85.140 160.680 85.280 161.160 ;
        RECT 74.930 160.540 85.280 160.680 ;
        RECT 74.930 160.480 75.250 160.540 ;
        RECT 84.145 160.495 84.435 160.540 ;
        RECT 18.280 159.860 93.120 160.340 ;
        RECT 69.410 159.660 69.730 159.720 ;
        RECT 75.390 159.660 75.710 159.720 ;
        RECT 69.410 159.520 79.300 159.660 ;
        RECT 69.410 159.460 69.730 159.520 ;
        RECT 75.390 159.460 75.710 159.520 ;
        RECT 53.325 159.320 53.615 159.365 ;
        RECT 60.210 159.320 60.530 159.380 ;
        RECT 70.345 159.320 70.635 159.365 ;
        RECT 53.325 159.180 70.635 159.320 ;
        RECT 53.325 159.135 53.615 159.180 ;
        RECT 60.210 159.120 60.530 159.180 ;
        RECT 70.345 159.135 70.635 159.180 ;
        RECT 38.100 158.980 38.390 159.025 ;
        RECT 43.190 158.980 43.510 159.040 ;
        RECT 38.100 158.840 43.510 158.980 ;
        RECT 38.100 158.795 38.390 158.840 ;
        RECT 43.190 158.780 43.510 158.840 ;
        RECT 52.390 158.980 52.710 159.040 ;
        RECT 54.705 158.980 54.995 159.025 ;
        RECT 56.530 158.980 56.850 159.040 ;
        RECT 79.160 159.025 79.300 159.520 ;
        RECT 80.470 159.320 80.760 159.365 ;
        RECT 81.870 159.320 82.160 159.365 ;
        RECT 83.710 159.320 84.000 159.365 ;
        RECT 80.470 159.180 84.000 159.320 ;
        RECT 80.470 159.135 80.760 159.180 ;
        RECT 81.870 159.135 82.160 159.180 ;
        RECT 83.710 159.135 84.000 159.180 ;
        RECT 52.390 158.840 56.850 158.980 ;
        RECT 52.390 158.780 52.710 158.840 ;
        RECT 54.705 158.795 54.995 158.840 ;
        RECT 56.530 158.780 56.850 158.840 ;
        RECT 79.085 158.980 79.375 159.025 ;
        RECT 79.545 158.980 79.835 159.025 ;
        RECT 79.085 158.840 82.060 158.980 ;
        RECT 79.085 158.795 79.375 158.840 ;
        RECT 79.545 158.795 79.835 158.840 ;
        RECT 81.920 158.700 82.060 158.840 ;
        RECT 36.765 158.455 37.055 158.685 ;
        RECT 37.645 158.640 37.935 158.685 ;
        RECT 38.835 158.640 39.125 158.685 ;
        RECT 41.355 158.640 41.645 158.685 ;
        RECT 55.610 158.640 55.930 158.700 ;
        RECT 37.645 158.500 41.645 158.640 ;
        RECT 37.645 158.455 37.935 158.500 ;
        RECT 38.835 158.455 39.125 158.500 ;
        RECT 41.355 158.455 41.645 158.500 ;
        RECT 46.960 158.500 55.930 158.640 ;
        RECT 36.840 157.960 36.980 158.455 ;
        RECT 46.960 158.345 47.100 158.500 ;
        RECT 55.610 158.440 55.930 158.500 ;
        RECT 80.450 158.640 80.770 158.700 ;
        RECT 80.925 158.640 81.215 158.685 ;
        RECT 80.450 158.500 81.215 158.640 ;
        RECT 80.450 158.440 80.770 158.500 ;
        RECT 80.925 158.455 81.215 158.500 ;
        RECT 81.830 158.440 82.150 158.700 ;
        RECT 37.250 158.300 37.540 158.345 ;
        RECT 39.350 158.300 39.640 158.345 ;
        RECT 40.920 158.300 41.210 158.345 ;
        RECT 46.885 158.300 47.175 158.345 ;
        RECT 37.250 158.160 41.210 158.300 ;
        RECT 37.250 158.115 37.540 158.160 ;
        RECT 39.350 158.115 39.640 158.160 ;
        RECT 40.920 158.115 41.210 158.160 ;
        RECT 43.050 158.160 47.175 158.300 ;
        RECT 38.130 157.960 38.450 158.020 ;
        RECT 43.050 157.960 43.190 158.160 ;
        RECT 46.885 158.115 47.175 158.160 ;
        RECT 47.330 158.300 47.650 158.360 ;
        RECT 80.010 158.300 80.300 158.345 ;
        RECT 82.330 158.300 82.620 158.345 ;
        RECT 83.710 158.300 84.000 158.345 ;
        RECT 47.330 158.160 55.840 158.300 ;
        RECT 47.330 158.100 47.650 158.160 ;
        RECT 36.840 157.820 43.190 157.960 ;
        RECT 43.665 157.960 43.955 158.005 ;
        RECT 50.090 157.960 50.410 158.020 ;
        RECT 55.700 158.005 55.840 158.160 ;
        RECT 80.010 158.160 84.000 158.300 ;
        RECT 80.010 158.115 80.300 158.160 ;
        RECT 82.330 158.115 82.620 158.160 ;
        RECT 83.710 158.115 84.000 158.160 ;
        RECT 43.665 157.820 50.410 157.960 ;
        RECT 38.130 157.760 38.450 157.820 ;
        RECT 43.665 157.775 43.955 157.820 ;
        RECT 50.090 157.760 50.410 157.820 ;
        RECT 55.625 157.960 55.915 158.005 ;
        RECT 56.530 157.960 56.850 158.020 ;
        RECT 55.625 157.820 56.850 157.960 ;
        RECT 55.625 157.775 55.915 157.820 ;
        RECT 56.530 157.760 56.850 157.820 ;
        RECT 69.870 157.960 70.190 158.020 ;
        RECT 75.850 157.960 76.170 158.020 ;
        RECT 69.870 157.820 76.170 157.960 ;
        RECT 69.870 157.760 70.190 157.820 ;
        RECT 75.850 157.760 76.170 157.820 ;
        RECT 87.365 157.960 87.655 158.005 ;
        RECT 87.810 157.960 88.130 158.020 ;
        RECT 87.365 157.820 88.130 157.960 ;
        RECT 87.365 157.775 87.655 157.820 ;
        RECT 87.810 157.760 88.130 157.820 ;
        RECT 18.280 157.140 92.340 157.620 ;
        RECT 43.190 156.940 43.510 157.000 ;
        RECT 45.505 156.940 45.795 156.985 ;
        RECT 72.170 156.940 72.490 157.000 ;
        RECT 77.690 156.940 78.010 157.000 ;
        RECT 43.190 156.800 45.795 156.940 ;
        RECT 43.190 156.740 43.510 156.800 ;
        RECT 45.505 156.755 45.795 156.800 ;
        RECT 56.620 156.800 67.340 156.940 ;
        RECT 56.620 156.660 56.760 156.800 ;
        RECT 56.530 156.400 56.850 156.660 ;
        RECT 59.330 156.600 59.620 156.645 ;
        RECT 61.430 156.600 61.720 156.645 ;
        RECT 63.000 156.600 63.290 156.645 ;
        RECT 59.330 156.460 63.290 156.600 ;
        RECT 59.330 156.415 59.620 156.460 ;
        RECT 61.430 156.415 61.720 156.460 ;
        RECT 63.000 156.415 63.290 156.460 ;
        RECT 67.200 156.600 67.340 156.800 ;
        RECT 72.170 156.800 78.010 156.940 ;
        RECT 72.170 156.740 72.490 156.800 ;
        RECT 77.690 156.740 78.010 156.800 ;
        RECT 82.305 156.600 82.595 156.645 ;
        RECT 67.200 156.460 70.560 156.600 ;
        RECT 50.090 156.260 50.410 156.320 ;
        RECT 51.945 156.260 52.235 156.305 ;
        RECT 50.090 156.120 52.235 156.260 ;
        RECT 50.090 156.060 50.410 156.120 ;
        RECT 51.945 156.075 52.235 156.120 ;
        RECT 55.610 156.260 55.930 156.320 ;
        RECT 58.845 156.260 59.135 156.305 ;
        RECT 55.610 156.120 59.135 156.260 ;
        RECT 55.610 156.060 55.930 156.120 ;
        RECT 58.845 156.075 59.135 156.120 ;
        RECT 59.725 156.260 60.015 156.305 ;
        RECT 60.915 156.260 61.205 156.305 ;
        RECT 63.435 156.260 63.725 156.305 ;
        RECT 59.725 156.120 63.725 156.260 ;
        RECT 59.725 156.075 60.015 156.120 ;
        RECT 60.915 156.075 61.205 156.120 ;
        RECT 63.435 156.075 63.725 156.120 ;
        RECT 66.205 156.075 66.495 156.305 ;
        RECT 43.650 155.920 43.970 155.980 ;
        RECT 44.570 155.920 44.890 155.980 ;
        RECT 43.650 155.780 44.890 155.920 ;
        RECT 43.650 155.720 43.970 155.780 ;
        RECT 44.570 155.720 44.890 155.780 ;
        RECT 45.490 155.720 45.810 155.980 ;
        RECT 46.885 155.920 47.175 155.965 ;
        RECT 47.345 155.920 47.635 155.965 ;
        RECT 46.885 155.780 47.635 155.920 ;
        RECT 46.885 155.735 47.175 155.780 ;
        RECT 47.345 155.735 47.635 155.780 ;
        RECT 52.865 155.920 53.155 155.965 ;
        RECT 56.990 155.920 57.310 155.980 ;
        RECT 52.865 155.780 57.310 155.920 ;
        RECT 52.865 155.735 53.155 155.780 ;
        RECT 56.990 155.720 57.310 155.780 ;
        RECT 57.465 155.735 57.755 155.965 ;
        RECT 58.385 155.920 58.675 155.965 ;
        RECT 66.280 155.920 66.420 156.075 ;
        RECT 67.200 155.965 67.340 156.460 ;
        RECT 68.045 156.075 68.335 156.305 ;
        RECT 58.385 155.780 66.420 155.920 ;
        RECT 58.385 155.735 58.675 155.780 ;
        RECT 67.125 155.735 67.415 155.965 ;
        RECT 54.230 155.580 54.550 155.640 ;
        RECT 54.705 155.580 54.995 155.625 ;
        RECT 52.020 155.440 54.995 155.580 ;
        RECT 52.020 155.300 52.160 155.440 ;
        RECT 54.230 155.380 54.550 155.440 ;
        RECT 54.705 155.395 54.995 155.440 ;
        RECT 46.425 155.240 46.715 155.285 ;
        RECT 48.250 155.240 48.570 155.300 ;
        RECT 46.425 155.100 48.570 155.240 ;
        RECT 46.425 155.055 46.715 155.100 ;
        RECT 48.250 155.040 48.570 155.100 ;
        RECT 51.930 155.040 52.250 155.300 ;
        RECT 52.850 155.240 53.170 155.300 ;
        RECT 53.325 155.240 53.615 155.285 ;
        RECT 52.850 155.100 53.615 155.240 ;
        RECT 52.850 155.040 53.170 155.100 ;
        RECT 53.325 155.055 53.615 155.100 ;
        RECT 53.770 155.040 54.090 155.300 ;
        RECT 57.540 155.240 57.680 155.735 ;
        RECT 67.570 155.720 67.890 155.980 ;
        RECT 68.120 155.920 68.260 156.075 ;
        RECT 68.490 156.060 68.810 156.320 ;
        RECT 68.950 155.920 69.270 155.980 ;
        RECT 68.120 155.780 69.270 155.920 ;
        RECT 68.950 155.720 69.270 155.780 ;
        RECT 69.410 155.720 69.730 155.980 ;
        RECT 69.885 155.735 70.175 155.965 ;
        RECT 70.420 155.920 70.560 156.460 ;
        RECT 75.480 156.460 82.595 156.600 ;
        RECT 75.480 156.305 75.620 156.460 ;
        RECT 82.305 156.415 82.595 156.460 ;
        RECT 75.405 156.075 75.695 156.305 ;
        RECT 75.850 156.060 76.170 156.320 ;
        RECT 80.465 156.260 80.755 156.305 ;
        RECT 80.465 156.120 83.440 156.260 ;
        RECT 80.465 156.075 80.755 156.120 ;
        RECT 74.485 155.920 74.775 155.965 ;
        RECT 70.420 155.780 74.775 155.920 ;
        RECT 74.485 155.735 74.775 155.780 ;
        RECT 57.925 155.580 58.215 155.625 ;
        RECT 60.070 155.580 60.360 155.625 ;
        RECT 69.960 155.580 70.100 155.735 ;
        RECT 74.930 155.720 75.250 155.980 ;
        RECT 76.785 155.735 77.075 155.965 ;
        RECT 57.925 155.440 60.360 155.580 ;
        RECT 57.925 155.395 58.215 155.440 ;
        RECT 60.070 155.395 60.360 155.440 ;
        RECT 65.820 155.440 70.100 155.580 ;
        RECT 71.710 155.580 72.030 155.640 ;
        RECT 76.860 155.580 77.000 155.735 ;
        RECT 77.230 155.720 77.550 155.980 ;
        RECT 77.690 155.920 78.010 155.980 ;
        RECT 83.300 155.965 83.440 156.120 ;
        RECT 80.925 155.920 81.215 155.965 ;
        RECT 77.690 155.780 81.215 155.920 ;
        RECT 77.690 155.720 78.010 155.780 ;
        RECT 80.925 155.735 81.215 155.780 ;
        RECT 83.225 155.735 83.515 155.965 ;
        RECT 71.710 155.440 75.620 155.580 ;
        RECT 76.860 155.440 82.060 155.580 ;
        RECT 65.820 155.300 65.960 155.440 ;
        RECT 71.710 155.380 72.030 155.440 ;
        RECT 65.270 155.240 65.590 155.300 ;
        RECT 57.540 155.100 65.590 155.240 ;
        RECT 65.270 155.040 65.590 155.100 ;
        RECT 65.730 155.040 66.050 155.300 ;
        RECT 72.630 155.240 72.950 155.300 ;
        RECT 73.105 155.240 73.395 155.285 ;
        RECT 72.630 155.100 73.395 155.240 ;
        RECT 72.630 155.040 72.950 155.100 ;
        RECT 73.105 155.055 73.395 155.100 ;
        RECT 73.565 155.240 73.855 155.285 ;
        RECT 74.930 155.240 75.250 155.300 ;
        RECT 73.565 155.100 75.250 155.240 ;
        RECT 75.480 155.240 75.620 155.440 ;
        RECT 81.385 155.240 81.675 155.285 ;
        RECT 75.480 155.100 81.675 155.240 ;
        RECT 81.920 155.240 82.060 155.440 ;
        RECT 82.290 155.380 82.610 155.640 ;
        RECT 83.685 155.240 83.975 155.285 ;
        RECT 81.920 155.100 83.975 155.240 ;
        RECT 73.565 155.055 73.855 155.100 ;
        RECT 74.930 155.040 75.250 155.100 ;
        RECT 81.385 155.055 81.675 155.100 ;
        RECT 83.685 155.055 83.975 155.100 ;
        RECT 18.280 154.420 93.120 154.900 ;
        RECT 45.490 154.220 45.810 154.280 ;
        RECT 46.425 154.220 46.715 154.265 ;
        RECT 45.490 154.080 46.715 154.220 ;
        RECT 45.490 154.020 45.810 154.080 ;
        RECT 46.425 154.035 46.715 154.080 ;
        RECT 48.250 154.020 48.570 154.280 ;
        RECT 53.310 154.020 53.630 154.280 ;
        RECT 53.770 154.220 54.090 154.280 ;
        RECT 56.545 154.220 56.835 154.265 ;
        RECT 53.770 154.080 56.835 154.220 ;
        RECT 53.770 154.020 54.090 154.080 ;
        RECT 56.545 154.035 56.835 154.080 ;
        RECT 56.990 154.020 57.310 154.280 ;
        RECT 67.585 154.220 67.875 154.265 ;
        RECT 69.870 154.220 70.190 154.280 ;
        RECT 67.585 154.080 70.190 154.220 ;
        RECT 67.585 154.035 67.875 154.080 ;
        RECT 42.745 153.880 43.035 153.925 ;
        RECT 46.870 153.880 47.190 153.940 ;
        RECT 42.745 153.740 47.190 153.880 ;
        RECT 48.340 153.880 48.480 154.020 ;
        RECT 53.400 153.880 53.540 154.020 ;
        RECT 48.340 153.740 49.860 153.880 ;
        RECT 42.745 153.695 43.035 153.740 ;
        RECT 46.870 153.680 47.190 153.740 ;
        RECT 40.430 153.540 40.750 153.600 ;
        RECT 41.825 153.540 42.115 153.585 ;
        RECT 42.270 153.540 42.590 153.600 ;
        RECT 40.430 153.400 42.590 153.540 ;
        RECT 40.430 153.340 40.750 153.400 ;
        RECT 41.825 153.355 42.115 153.400 ;
        RECT 42.270 153.340 42.590 153.400 ;
        RECT 43.205 153.355 43.495 153.585 ;
        RECT 41.810 152.320 42.130 152.580 ;
        RECT 43.280 152.520 43.420 153.355 ;
        RECT 47.330 153.340 47.650 153.600 ;
        RECT 48.710 153.340 49.030 153.600 ;
        RECT 49.720 153.585 49.860 153.740 ;
        RECT 51.560 153.740 53.540 153.880 ;
        RECT 54.690 153.880 55.010 153.940 ;
        RECT 57.080 153.880 57.220 154.020 ;
        RECT 54.690 153.740 57.220 153.880 ;
        RECT 51.560 153.585 51.700 153.740 ;
        RECT 54.690 153.680 55.010 153.740 ;
        RECT 49.645 153.355 49.935 153.585 ;
        RECT 51.485 153.355 51.775 153.585 ;
        RECT 52.390 153.340 52.710 153.600 ;
        RECT 52.865 153.355 53.155 153.585 ;
        RECT 53.310 153.540 53.630 153.600 ;
        RECT 54.245 153.540 54.535 153.585 ;
        RECT 53.310 153.400 54.535 153.540 ;
        RECT 48.265 153.200 48.555 153.245 ;
        RECT 51.930 153.200 52.250 153.260 ;
        RECT 48.265 153.060 52.250 153.200 ;
        RECT 48.265 153.015 48.555 153.060 ;
        RECT 51.930 153.000 52.250 153.060 ;
        RECT 47.805 152.860 48.095 152.905 ;
        RECT 52.480 152.860 52.620 153.340 ;
        RECT 52.940 152.920 53.080 153.355 ;
        RECT 53.310 153.340 53.630 153.400 ;
        RECT 54.245 153.355 54.535 153.400 ;
        RECT 55.150 153.540 55.470 153.600 ;
        RECT 57.465 153.540 57.755 153.585 ;
        RECT 55.150 153.400 57.755 153.540 ;
        RECT 47.805 152.720 52.620 152.860 ;
        RECT 47.805 152.675 48.095 152.720 ;
        RECT 52.850 152.660 53.170 152.920 ;
        RECT 50.105 152.520 50.395 152.565 ;
        RECT 43.280 152.380 50.395 152.520 ;
        RECT 50.105 152.335 50.395 152.380 ;
        RECT 51.470 152.320 51.790 152.580 ;
        RECT 54.320 152.520 54.460 153.355 ;
        RECT 55.150 153.340 55.470 153.400 ;
        RECT 57.465 153.355 57.755 153.400 ;
        RECT 65.730 153.540 66.050 153.600 ;
        RECT 66.205 153.540 66.495 153.585 ;
        RECT 65.730 153.400 66.495 153.540 ;
        RECT 65.730 153.340 66.050 153.400 ;
        RECT 66.205 153.355 66.495 153.400 ;
        RECT 67.125 153.540 67.415 153.585 ;
        RECT 67.660 153.540 67.800 154.035 ;
        RECT 69.870 154.020 70.190 154.080 ;
        RECT 71.710 154.020 72.030 154.280 ;
        RECT 72.170 154.020 72.490 154.280 ;
        RECT 77.230 154.220 77.550 154.280 ;
        RECT 82.290 154.220 82.610 154.280 ;
        RECT 74.100 154.080 82.610 154.220 ;
        RECT 68.425 153.880 68.715 153.925 ;
        RECT 69.425 153.880 69.715 153.925 ;
        RECT 71.265 153.880 71.555 153.925 ;
        RECT 74.100 153.880 74.240 154.080 ;
        RECT 77.230 154.020 77.550 154.080 ;
        RECT 82.290 154.020 82.610 154.080 ;
        RECT 68.425 153.740 69.180 153.880 ;
        RECT 68.425 153.695 68.715 153.740 ;
        RECT 67.125 153.400 67.800 153.540 ;
        RECT 69.040 153.540 69.180 153.740 ;
        RECT 69.425 153.740 74.240 153.880 ;
        RECT 74.470 153.880 74.790 153.940 ;
        RECT 76.630 153.880 76.920 153.925 ;
        RECT 74.470 153.740 76.920 153.880 ;
        RECT 69.425 153.695 69.715 153.740 ;
        RECT 71.265 153.695 71.555 153.740 ;
        RECT 74.470 153.680 74.790 153.740 ;
        RECT 76.630 153.695 76.920 153.740 ;
        RECT 72.170 153.540 72.490 153.600 ;
        RECT 69.040 153.400 72.490 153.540 ;
        RECT 67.125 153.355 67.415 153.400 ;
        RECT 56.070 153.200 56.390 153.260 ;
        RECT 58.385 153.200 58.675 153.245 ;
        RECT 56.070 153.060 58.675 153.200 ;
        RECT 66.280 153.200 66.420 153.355 ;
        RECT 72.170 153.340 72.490 153.400 ;
        RECT 72.630 153.540 72.950 153.600 ;
        RECT 74.025 153.540 74.315 153.585 ;
        RECT 72.630 153.400 74.315 153.540 ;
        RECT 72.630 153.340 72.950 153.400 ;
        RECT 74.025 153.355 74.315 153.400 ;
        RECT 75.390 153.340 75.710 153.600 ;
        RECT 70.345 153.200 70.635 153.245 ;
        RECT 76.285 153.200 76.575 153.245 ;
        RECT 77.475 153.200 77.765 153.245 ;
        RECT 79.995 153.200 80.285 153.245 ;
        RECT 66.280 153.060 70.635 153.200 ;
        RECT 56.070 153.000 56.390 153.060 ;
        RECT 58.385 153.015 58.675 153.060 ;
        RECT 70.345 153.015 70.635 153.060 ;
        RECT 72.720 153.060 74.700 153.200 ;
        RECT 67.125 152.860 67.415 152.905 ;
        RECT 68.950 152.860 69.270 152.920 ;
        RECT 67.125 152.720 69.270 152.860 ;
        RECT 67.125 152.675 67.415 152.720 ;
        RECT 68.950 152.660 69.270 152.720 ;
        RECT 69.410 152.860 69.730 152.920 ;
        RECT 72.720 152.860 72.860 153.060 ;
        RECT 69.410 152.720 72.860 152.860 ;
        RECT 69.410 152.660 69.730 152.720 ;
        RECT 73.090 152.660 73.410 152.920 ;
        RECT 74.560 152.905 74.700 153.060 ;
        RECT 76.285 153.060 80.285 153.200 ;
        RECT 76.285 153.015 76.575 153.060 ;
        RECT 77.475 153.015 77.765 153.060 ;
        RECT 79.995 153.015 80.285 153.060 ;
        RECT 74.485 152.675 74.775 152.905 ;
        RECT 75.890 152.860 76.180 152.905 ;
        RECT 77.990 152.860 78.280 152.905 ;
        RECT 79.560 152.860 79.850 152.905 ;
        RECT 75.890 152.720 79.850 152.860 ;
        RECT 75.890 152.675 76.180 152.720 ;
        RECT 77.990 152.675 78.280 152.720 ;
        RECT 79.560 152.675 79.850 152.720 ;
        RECT 62.970 152.520 63.290 152.580 ;
        RECT 54.320 152.380 63.290 152.520 ;
        RECT 62.970 152.320 63.290 152.380 ;
        RECT 68.505 152.520 68.795 152.565 ;
        RECT 71.710 152.520 72.030 152.580 ;
        RECT 68.505 152.380 72.030 152.520 ;
        RECT 68.505 152.335 68.795 152.380 ;
        RECT 71.710 152.320 72.030 152.380 ;
        RECT 18.280 151.700 92.340 152.180 ;
        RECT 42.270 151.500 42.590 151.560 ;
        RECT 46.870 151.500 47.190 151.560 ;
        RECT 48.725 151.500 49.015 151.545 ;
        RECT 42.270 151.360 46.640 151.500 ;
        RECT 42.270 151.300 42.590 151.360 ;
        RECT 37.250 151.160 37.540 151.205 ;
        RECT 39.350 151.160 39.640 151.205 ;
        RECT 40.920 151.160 41.210 151.205 ;
        RECT 37.250 151.020 41.210 151.160 ;
        RECT 37.250 150.975 37.540 151.020 ;
        RECT 39.350 150.975 39.640 151.020 ;
        RECT 40.920 150.975 41.210 151.020 ;
        RECT 43.665 150.975 43.955 151.205 ;
        RECT 46.500 151.160 46.640 151.360 ;
        RECT 46.870 151.360 49.015 151.500 ;
        RECT 46.870 151.300 47.190 151.360 ;
        RECT 48.725 151.315 49.015 151.360 ;
        RECT 50.105 151.500 50.395 151.545 ;
        RECT 52.850 151.500 53.170 151.560 ;
        RECT 50.105 151.360 53.170 151.500 ;
        RECT 50.105 151.315 50.395 151.360 ;
        RECT 52.850 151.300 53.170 151.360 ;
        RECT 72.170 151.300 72.490 151.560 ;
        RECT 74.025 151.500 74.315 151.545 ;
        RECT 74.470 151.500 74.790 151.560 ;
        RECT 74.025 151.360 74.790 151.500 ;
        RECT 74.025 151.315 74.315 151.360 ;
        RECT 74.470 151.300 74.790 151.360 ;
        RECT 74.930 151.300 75.250 151.560 ;
        RECT 59.290 151.160 59.610 151.220 ;
        RECT 46.500 151.020 59.610 151.160 ;
        RECT 37.645 150.820 37.935 150.865 ;
        RECT 38.835 150.820 39.125 150.865 ;
        RECT 41.355 150.820 41.645 150.865 ;
        RECT 37.645 150.680 41.645 150.820 ;
        RECT 43.740 150.820 43.880 150.975 ;
        RECT 59.290 150.960 59.610 151.020 ;
        RECT 60.210 150.960 60.530 151.220 ;
        RECT 45.045 150.820 45.335 150.865 ;
        RECT 52.405 150.820 52.695 150.865 ;
        RECT 56.070 150.820 56.390 150.880 ;
        RECT 70.805 150.820 71.095 150.865 ;
        RECT 72.260 150.820 72.400 151.300 ;
        RECT 75.020 150.820 75.160 151.300 ;
        RECT 43.740 150.680 56.390 150.820 ;
        RECT 37.645 150.635 37.935 150.680 ;
        RECT 38.835 150.635 39.125 150.680 ;
        RECT 41.355 150.635 41.645 150.680 ;
        RECT 45.045 150.635 45.335 150.680 ;
        RECT 52.405 150.635 52.695 150.680 ;
        RECT 56.070 150.620 56.390 150.680 ;
        RECT 57.080 150.680 62.280 150.820 ;
        RECT 36.765 150.295 37.055 150.525 ;
        RECT 38.100 150.480 38.390 150.525 ;
        RECT 41.810 150.480 42.130 150.540 ;
        RECT 38.100 150.340 42.130 150.480 ;
        RECT 38.100 150.295 38.390 150.340 ;
        RECT 36.840 150.140 36.980 150.295 ;
        RECT 41.810 150.280 42.130 150.340 ;
        RECT 44.110 150.280 44.430 150.540 ;
        RECT 47.805 150.480 48.095 150.525 ;
        RECT 48.265 150.480 48.555 150.525 ;
        RECT 49.140 150.480 49.430 150.525 ;
        RECT 47.805 150.340 48.555 150.480 ;
        RECT 47.805 150.295 48.095 150.340 ;
        RECT 48.265 150.295 48.555 150.340 ;
        RECT 48.800 150.340 49.430 150.480 ;
        RECT 44.200 150.140 44.340 150.280 ;
        RECT 48.800 150.200 48.940 150.340 ;
        RECT 49.140 150.295 49.430 150.340 ;
        RECT 51.025 150.295 51.315 150.525 ;
        RECT 51.485 150.295 51.775 150.525 ;
        RECT 51.945 150.480 52.235 150.525 ;
        RECT 55.150 150.480 55.470 150.540 ;
        RECT 56.530 150.480 56.850 150.540 ;
        RECT 51.945 150.340 56.850 150.480 ;
        RECT 51.945 150.295 52.235 150.340 ;
        RECT 48.710 150.140 49.030 150.200 ;
        RECT 36.840 150.000 38.360 150.140 ;
        RECT 44.200 150.000 49.030 150.140 ;
        RECT 38.220 149.860 38.360 150.000 ;
        RECT 48.710 149.940 49.030 150.000 ;
        RECT 38.130 149.600 38.450 149.860 ;
        RECT 51.100 149.800 51.240 150.295 ;
        RECT 51.560 150.140 51.700 150.295 ;
        RECT 55.150 150.280 55.470 150.340 ;
        RECT 56.530 150.280 56.850 150.340 ;
        RECT 53.770 150.140 54.090 150.200 ;
        RECT 54.690 150.140 55.010 150.200 ;
        RECT 57.080 150.140 57.220 150.680 ;
        RECT 61.590 150.280 61.910 150.540 ;
        RECT 62.140 150.525 62.280 150.680 ;
        RECT 70.805 150.680 72.400 150.820 ;
        RECT 74.100 150.680 75.160 150.820 ;
        RECT 70.805 150.635 71.095 150.680 ;
        RECT 62.065 150.295 62.355 150.525 ;
        RECT 62.970 150.480 63.290 150.540 ;
        RECT 67.570 150.480 67.890 150.540 ;
        RECT 62.970 150.340 67.890 150.480 ;
        RECT 62.970 150.280 63.290 150.340 ;
        RECT 67.570 150.280 67.890 150.340 ;
        RECT 68.030 150.280 68.350 150.540 ;
        RECT 70.345 150.480 70.635 150.525 ;
        RECT 71.710 150.480 72.030 150.540 ;
        RECT 74.100 150.525 74.240 150.680 ;
        RECT 70.345 150.340 72.030 150.480 ;
        RECT 70.345 150.295 70.635 150.340 ;
        RECT 71.710 150.280 72.030 150.340 ;
        RECT 74.025 150.295 74.315 150.525 ;
        RECT 74.930 150.480 75.250 150.540 ;
        RECT 79.990 150.480 80.310 150.540 ;
        RECT 74.930 150.340 80.310 150.480 ;
        RECT 74.930 150.280 75.250 150.340 ;
        RECT 79.990 150.280 80.310 150.340 ;
        RECT 51.560 150.000 57.220 150.140 ;
        RECT 59.290 150.140 59.610 150.200 ;
        RECT 60.225 150.140 60.515 150.185 ;
        RECT 68.120 150.140 68.260 150.280 ;
        RECT 59.290 150.000 68.260 150.140 ;
        RECT 53.770 149.940 54.090 150.000 ;
        RECT 54.690 149.940 55.010 150.000 ;
        RECT 59.290 149.940 59.610 150.000 ;
        RECT 60.225 149.955 60.515 150.000 ;
        RECT 53.310 149.800 53.630 149.860 ;
        RECT 51.100 149.660 53.630 149.800 ;
        RECT 53.310 149.600 53.630 149.660 ;
        RECT 61.130 149.600 61.450 149.860 ;
        RECT 62.510 149.600 62.830 149.860 ;
        RECT 72.170 149.600 72.490 149.860 ;
        RECT 18.280 148.980 93.120 149.460 ;
        RECT 53.310 148.580 53.630 148.840 ;
        RECT 56.085 148.780 56.375 148.825 ;
        RECT 61.130 148.780 61.450 148.840 ;
        RECT 56.085 148.640 61.450 148.780 ;
        RECT 56.085 148.595 56.375 148.640 ;
        RECT 61.130 148.580 61.450 148.640 ;
        RECT 61.590 148.780 61.910 148.840 ;
        RECT 63.445 148.780 63.735 148.825 ;
        RECT 61.590 148.640 63.735 148.780 ;
        RECT 61.590 148.580 61.910 148.640 ;
        RECT 63.445 148.595 63.735 148.640 ;
        RECT 65.285 148.780 65.575 148.825 ;
        RECT 66.650 148.780 66.970 148.840 ;
        RECT 71.265 148.780 71.555 148.825 ;
        RECT 71.710 148.780 72.030 148.840 ;
        RECT 65.285 148.640 68.720 148.780 ;
        RECT 65.285 148.595 65.575 148.640 ;
        RECT 66.650 148.580 66.970 148.640 ;
        RECT 53.400 148.100 53.540 148.580 ;
        RECT 54.245 148.440 54.535 148.485 ;
        RECT 55.150 148.440 55.470 148.500 ;
        RECT 65.745 148.440 66.035 148.485 ;
        RECT 68.030 148.440 68.350 148.500 ;
        RECT 54.245 148.300 60.900 148.440 ;
        RECT 54.245 148.255 54.535 148.300 ;
        RECT 55.150 148.240 55.470 148.300 ;
        RECT 60.760 148.145 60.900 148.300 ;
        RECT 61.220 148.300 63.200 148.440 ;
        RECT 61.220 148.160 61.360 148.300 ;
        RECT 53.785 148.100 54.075 148.145 ;
        RECT 54.745 148.100 55.035 148.145 ;
        RECT 55.625 148.100 55.915 148.145 ;
        RECT 53.400 147.960 54.075 148.100 ;
        RECT 53.785 147.915 54.075 147.960 ;
        RECT 54.320 147.960 55.035 148.100 ;
        RECT 54.320 147.820 54.460 147.960 ;
        RECT 54.745 147.915 55.035 147.960 ;
        RECT 55.240 147.960 55.915 148.100 ;
        RECT 54.230 147.560 54.550 147.820 ;
        RECT 48.710 147.420 49.030 147.480 ;
        RECT 55.240 147.420 55.380 147.960 ;
        RECT 55.625 147.915 55.915 147.960 ;
        RECT 56.545 148.100 56.835 148.145 ;
        RECT 57.005 148.100 57.295 148.145 ;
        RECT 56.545 147.960 57.295 148.100 ;
        RECT 56.545 147.915 56.835 147.960 ;
        RECT 57.005 147.915 57.295 147.960 ;
        RECT 60.685 147.915 60.975 148.145 ;
        RECT 61.130 147.900 61.450 148.160 ;
        RECT 62.510 147.900 62.830 148.160 ;
        RECT 63.060 148.100 63.200 148.300 ;
        RECT 65.745 148.300 68.350 148.440 ;
        RECT 68.580 148.440 68.720 148.640 ;
        RECT 71.265 148.640 72.030 148.780 ;
        RECT 71.265 148.595 71.555 148.640 ;
        RECT 71.710 148.580 72.030 148.640 ;
        RECT 74.930 148.580 75.250 148.840 ;
        RECT 75.020 148.440 75.160 148.580 ;
        RECT 68.580 148.300 75.160 148.440 ;
        RECT 65.745 148.255 66.035 148.300 ;
        RECT 68.030 148.240 68.350 148.300 ;
        RECT 70.970 148.100 71.260 148.145 ;
        RECT 63.060 147.960 71.260 148.100 ;
        RECT 70.970 147.915 71.260 147.960 ;
        RECT 72.170 148.100 72.490 148.160 ;
        RECT 73.105 148.100 73.395 148.145 ;
        RECT 72.170 147.960 73.395 148.100 ;
        RECT 72.170 147.900 72.490 147.960 ;
        RECT 73.105 147.915 73.395 147.960 ;
        RECT 59.290 147.760 59.610 147.820 ;
        RECT 59.765 147.760 60.055 147.805 ;
        RECT 59.290 147.620 60.055 147.760 ;
        RECT 59.290 147.560 59.610 147.620 ;
        RECT 59.765 147.575 60.055 147.620 ;
        RECT 73.565 147.575 73.855 147.805 ;
        RECT 60.670 147.420 60.990 147.480 ;
        RECT 73.640 147.420 73.780 147.575 ;
        RECT 48.710 147.280 60.990 147.420 ;
        RECT 48.710 147.220 49.030 147.280 ;
        RECT 60.670 147.220 60.990 147.280 ;
        RECT 61.220 147.280 73.780 147.420 ;
        RECT 53.310 147.080 53.630 147.140 ;
        RECT 56.990 147.080 57.310 147.140 ;
        RECT 61.220 147.125 61.360 147.280 ;
        RECT 61.145 147.080 61.435 147.125 ;
        RECT 53.310 146.940 61.435 147.080 ;
        RECT 53.310 146.880 53.630 146.940 ;
        RECT 56.990 146.880 57.310 146.940 ;
        RECT 61.145 146.895 61.435 146.940 ;
        RECT 70.330 146.880 70.650 147.140 ;
        RECT 131.170 147.000 131.835 147.605 ;
        RECT 18.280 146.260 92.340 146.740 ;
        RECT 53.770 146.060 54.090 146.120 ;
        RECT 57.465 146.060 57.755 146.105 ;
        RECT 59.290 146.060 59.610 146.120 ;
        RECT 53.770 145.920 59.610 146.060 ;
        RECT 53.770 145.860 54.090 145.920 ;
        RECT 57.465 145.875 57.755 145.920 ;
        RECT 59.290 145.860 59.610 145.920 ;
        RECT 71.710 146.060 72.030 146.120 ;
        RECT 72.185 146.060 72.475 146.105 ;
        RECT 71.710 145.920 72.475 146.060 ;
        RECT 71.710 145.860 72.030 145.920 ;
        RECT 72.185 145.875 72.475 145.920 ;
        RECT 108.700 145.830 109.300 145.860 ;
        RECT 43.230 145.720 43.520 145.765 ;
        RECT 45.330 145.720 45.620 145.765 ;
        RECT 46.900 145.720 47.190 145.765 ;
        RECT 43.230 145.580 47.190 145.720 ;
        RECT 43.230 145.535 43.520 145.580 ;
        RECT 45.330 145.535 45.620 145.580 ;
        RECT 46.900 145.535 47.190 145.580 ;
        RECT 60.210 145.720 60.500 145.765 ;
        RECT 61.780 145.720 62.070 145.765 ;
        RECT 63.880 145.720 64.170 145.765 ;
        RECT 60.210 145.580 64.170 145.720 ;
        RECT 60.210 145.535 60.500 145.580 ;
        RECT 61.780 145.535 62.070 145.580 ;
        RECT 63.880 145.535 64.170 145.580 ;
        RECT 65.770 145.720 66.060 145.765 ;
        RECT 67.870 145.720 68.160 145.765 ;
        RECT 69.440 145.720 69.730 145.765 ;
        RECT 65.770 145.580 69.730 145.720 ;
        RECT 65.770 145.535 66.060 145.580 ;
        RECT 67.870 145.535 68.160 145.580 ;
        RECT 69.440 145.535 69.730 145.580 ;
        RECT 38.130 145.380 38.450 145.440 ;
        RECT 42.745 145.380 43.035 145.425 ;
        RECT 38.130 145.240 43.035 145.380 ;
        RECT 38.130 145.180 38.450 145.240 ;
        RECT 42.745 145.195 43.035 145.240 ;
        RECT 43.625 145.380 43.915 145.425 ;
        RECT 44.815 145.380 45.105 145.425 ;
        RECT 47.335 145.380 47.625 145.425 ;
        RECT 43.625 145.240 47.625 145.380 ;
        RECT 43.625 145.195 43.915 145.240 ;
        RECT 44.815 145.195 45.105 145.240 ;
        RECT 47.335 145.195 47.625 145.240 ;
        RECT 52.865 145.380 53.155 145.425 ;
        RECT 53.785 145.380 54.075 145.425 ;
        RECT 52.865 145.240 54.075 145.380 ;
        RECT 52.865 145.195 53.155 145.240 ;
        RECT 53.785 145.195 54.075 145.240 ;
        RECT 55.150 145.180 55.470 145.440 ;
        RECT 59.775 145.380 60.065 145.425 ;
        RECT 62.295 145.380 62.585 145.425 ;
        RECT 63.485 145.380 63.775 145.425 ;
        RECT 59.775 145.240 63.775 145.380 ;
        RECT 59.775 145.195 60.065 145.240 ;
        RECT 62.295 145.195 62.585 145.240 ;
        RECT 63.485 145.195 63.775 145.240 ;
        RECT 66.165 145.380 66.455 145.425 ;
        RECT 67.355 145.380 67.645 145.425 ;
        RECT 69.875 145.380 70.165 145.425 ;
        RECT 66.165 145.240 70.165 145.380 ;
        RECT 66.165 145.195 66.455 145.240 ;
        RECT 67.355 145.195 67.645 145.240 ;
        RECT 69.875 145.195 70.165 145.240 ;
        RECT 75.390 145.180 75.710 145.440 ;
        RECT 108.700 145.230 110.800 145.830 ;
        RECT 113.170 145.800 113.830 146.400 ;
        RECT 116.370 145.900 117.030 146.500 ;
        RECT 119.270 146.000 119.930 146.600 ;
        RECT 108.700 145.200 109.300 145.230 ;
        RECT 48.710 145.040 49.030 145.100 ;
        RECT 50.730 145.040 51.020 145.085 ;
        RECT 48.710 144.900 51.020 145.040 ;
        RECT 48.710 144.840 49.030 144.900 ;
        RECT 50.730 144.855 51.020 144.900 ;
        RECT 53.310 144.840 53.630 145.100 ;
        RECT 55.625 145.040 55.915 145.085 ;
        RECT 56.530 145.040 56.850 145.100 ;
        RECT 55.625 144.900 56.850 145.040 ;
        RECT 55.625 144.855 55.915 144.900 ;
        RECT 44.080 144.700 44.370 144.745 ;
        RECT 45.030 144.700 45.350 144.760 ;
        RECT 44.080 144.560 45.350 144.700 ;
        RECT 44.080 144.515 44.370 144.560 ;
        RECT 45.030 144.500 45.350 144.560 ;
        RECT 49.720 144.560 51.240 144.700 ;
        RECT 49.720 144.405 49.860 144.560 ;
        RECT 49.645 144.175 49.935 144.405 ;
        RECT 50.090 144.160 50.410 144.420 ;
        RECT 51.100 144.405 51.240 144.560 ;
        RECT 51.025 144.360 51.315 144.405 ;
        RECT 55.700 144.360 55.840 144.855 ;
        RECT 56.530 144.840 56.850 144.900 ;
        RECT 60.210 145.040 60.530 145.100 ;
        RECT 63.030 145.040 63.320 145.085 ;
        RECT 60.210 144.900 63.320 145.040 ;
        RECT 60.210 144.840 60.530 144.900 ;
        RECT 63.030 144.855 63.320 144.900 ;
        RECT 64.365 145.040 64.655 145.085 ;
        RECT 65.285 145.040 65.575 145.085 ;
        RECT 75.480 145.040 75.620 145.180 ;
        RECT 64.365 144.900 75.620 145.040 ;
        RECT 110.200 145.000 110.800 145.230 ;
        RECT 113.200 145.000 113.800 145.800 ;
        RECT 116.400 145.000 117.000 145.900 ;
        RECT 119.300 145.000 119.900 146.000 ;
        RECT 122.270 145.900 122.930 146.500 ;
        RECT 125.270 145.900 125.930 146.500 ;
        RECT 128.270 145.900 128.930 146.500 ;
        RECT 122.300 145.000 122.900 145.900 ;
        RECT 125.300 145.000 125.900 145.900 ;
        RECT 128.300 145.000 128.900 145.900 ;
        RECT 131.200 145.000 131.805 147.000 ;
        RECT 64.365 144.855 64.655 144.900 ;
        RECT 65.285 144.855 65.575 144.900 ;
        RECT 66.620 144.700 66.910 144.745 ;
        RECT 67.110 144.700 67.430 144.760 ;
        RECT 66.620 144.560 67.430 144.700 ;
        RECT 66.620 144.515 66.910 144.560 ;
        RECT 67.110 144.500 67.430 144.560 ;
        RECT 51.025 144.220 55.840 144.360 ;
        RECT 51.025 144.175 51.315 144.220 ;
        RECT 18.280 143.540 93.120 144.020 ;
        RECT 110.000 144.000 111.200 145.000 ;
        RECT 113.000 144.000 114.200 145.000 ;
        RECT 116.000 144.000 117.200 145.000 ;
        RECT 119.000 144.000 120.200 145.000 ;
        RECT 122.000 144.000 123.200 145.000 ;
        RECT 125.000 144.000 126.200 145.000 ;
        RECT 128.000 144.000 129.200 145.000 ;
        RECT 131.000 144.000 132.200 145.000 ;
        RECT 45.030 143.140 45.350 143.400 ;
        RECT 67.110 143.140 67.430 143.400 ;
        RECT 44.570 142.460 44.890 142.720 ;
        RECT 45.505 142.660 45.795 142.705 ;
        RECT 50.090 142.660 50.410 142.720 ;
        RECT 45.505 142.520 50.410 142.660 ;
        RECT 45.505 142.475 45.795 142.520 ;
        RECT 50.090 142.460 50.410 142.520 ;
        RECT 66.650 142.460 66.970 142.720 ;
        RECT 67.585 142.660 67.875 142.705 ;
        RECT 70.330 142.660 70.650 142.720 ;
        RECT 67.585 142.520 70.650 142.660 ;
        RECT 67.585 142.475 67.875 142.520 ;
        RECT 70.330 142.460 70.650 142.520 ;
        RECT 44.660 142.320 44.800 142.460 ;
        RECT 66.740 142.320 66.880 142.460 ;
        RECT 44.660 142.180 66.880 142.320 ;
        RECT 18.280 140.820 92.340 141.300 ;
        RECT 110.800 139.300 111.200 144.000 ;
        RECT 113.800 139.300 114.200 144.000 ;
        RECT 116.800 139.300 117.200 144.000 ;
        RECT 119.800 139.300 120.200 144.000 ;
        RECT 122.800 139.300 123.200 144.000 ;
        RECT 125.800 139.300 126.200 144.000 ;
        RECT 128.800 139.300 129.200 144.000 ;
        RECT 131.800 139.300 132.200 144.000 ;
        RECT 110.880 139.015 111.130 139.300 ;
        RECT 113.880 139.015 114.130 139.300 ;
        RECT 116.880 139.015 117.130 139.300 ;
        RECT 119.880 139.015 120.130 139.300 ;
        RECT 122.880 139.015 123.130 139.300 ;
        RECT 125.880 139.015 126.130 139.300 ;
        RECT 128.880 139.015 129.130 139.300 ;
        RECT 131.880 139.015 132.130 139.300 ;
        RECT 18.280 138.100 93.120 138.580 ;
        RECT 18.280 135.380 92.340 135.860 ;
        RECT 18.280 132.660 93.120 133.140 ;
        RECT 106.800 115.100 109.100 115.500 ;
        RECT 106.800 112.300 107.200 115.100 ;
        RECT 106.880 112.015 107.130 112.300 ;
        RECT 108.700 98.000 109.100 115.100 ;
        RECT 110.880 98.000 111.130 98.965 ;
        RECT 113.880 98.000 114.130 98.965 ;
        RECT 116.880 98.000 117.130 98.965 ;
        RECT 119.880 98.000 120.130 98.965 ;
        RECT 122.880 98.000 123.130 98.965 ;
        RECT 125.880 98.000 126.130 98.965 ;
        RECT 128.880 98.100 129.130 98.965 ;
        RECT 131.880 98.100 132.130 98.965 ;
        RECT 108.700 97.600 111.200 98.000 ;
        RECT 110.800 92.200 111.200 97.600 ;
        RECT 112.300 97.600 114.200 98.000 ;
        RECT 110.880 92.015 111.130 92.200 ;
        RECT 102.970 77.700 104.030 78.700 ;
        RECT 103.000 70.700 104.000 77.700 ;
        RECT 106.880 71.600 107.130 71.965 ;
        RECT 106.800 70.700 107.200 71.600 ;
        RECT 110.880 70.700 111.130 71.965 ;
        RECT 112.300 70.700 112.700 97.600 ;
        RECT 113.880 96.860 114.130 97.600 ;
        RECT 113.880 93.300 114.130 94.120 ;
        RECT 116.800 93.300 117.200 98.000 ;
        RECT 113.800 92.900 117.200 93.300 ;
        RECT 113.880 92.015 114.130 92.900 ;
        RECT 116.800 92.200 117.200 92.900 ;
        RECT 118.300 97.600 120.200 98.000 ;
        RECT 116.880 92.015 117.130 92.200 ;
        RECT 113.880 70.700 114.130 71.965 ;
        RECT 116.880 70.700 117.130 71.965 ;
        RECT 118.300 70.700 118.700 97.600 ;
        RECT 119.880 96.860 120.130 97.600 ;
        RECT 119.880 93.300 120.130 94.120 ;
        RECT 122.800 93.300 123.200 98.000 ;
        RECT 119.800 92.900 123.200 93.300 ;
        RECT 119.880 92.015 120.130 92.900 ;
        RECT 122.800 92.200 123.200 92.900 ;
        RECT 124.300 97.600 126.200 98.000 ;
        RECT 122.880 92.015 123.130 92.200 ;
        RECT 119.880 70.700 120.130 71.965 ;
        RECT 122.880 70.700 123.130 71.965 ;
        RECT 124.300 70.700 124.700 97.600 ;
        RECT 125.880 96.860 126.130 97.600 ;
        RECT 125.880 93.300 126.130 94.120 ;
        RECT 128.800 93.300 129.200 98.100 ;
        RECT 125.800 92.900 129.200 93.300 ;
        RECT 125.880 92.015 126.130 92.900 ;
        RECT 128.800 92.300 129.200 92.900 ;
        RECT 131.800 94.700 132.200 98.100 ;
        RECT 136.000 97.800 137.000 98.000 ;
        RECT 136.000 97.200 138.500 97.800 ;
        RECT 136.000 97.000 137.000 97.200 ;
        RECT 136.000 94.700 136.400 97.000 ;
        RECT 131.800 94.300 136.400 94.700 ;
        RECT 128.880 92.015 129.130 92.300 ;
        RECT 125.880 70.700 126.130 71.965 ;
        RECT 128.880 71.500 129.130 71.965 ;
        RECT 128.800 70.800 129.200 71.500 ;
        RECT 131.800 70.800 132.200 94.300 ;
        RECT 103.000 70.300 107.200 70.700 ;
        RECT 110.800 70.300 114.200 70.700 ;
        RECT 116.800 70.300 120.200 70.700 ;
        RECT 122.800 70.300 126.200 70.700 ;
        RECT 128.800 70.400 132.200 70.800 ;
        RECT 103.000 69.900 104.000 70.300 ;
        RECT 106.880 69.860 107.130 70.300 ;
        RECT 110.880 69.860 111.130 70.300 ;
        RECT 113.880 69.860 114.130 70.300 ;
        RECT 116.880 69.860 117.130 70.300 ;
        RECT 119.880 69.860 120.130 70.300 ;
        RECT 122.880 69.860 123.130 70.300 ;
        RECT 125.880 69.860 126.130 70.300 ;
        RECT 128.880 69.860 129.130 70.400 ;
        RECT 137.900 35.670 138.500 97.200 ;
      LAYER via ;
        RECT 26.765 206.210 27.025 206.470 ;
        RECT 27.085 206.210 27.345 206.470 ;
        RECT 27.405 206.210 27.665 206.470 ;
        RECT 27.725 206.210 27.985 206.470 ;
        RECT 28.045 206.210 28.305 206.470 ;
        RECT 45.275 206.210 45.535 206.470 ;
        RECT 45.595 206.210 45.855 206.470 ;
        RECT 45.915 206.210 46.175 206.470 ;
        RECT 46.235 206.210 46.495 206.470 ;
        RECT 46.555 206.210 46.815 206.470 ;
        RECT 63.785 206.210 64.045 206.470 ;
        RECT 64.105 206.210 64.365 206.470 ;
        RECT 64.425 206.210 64.685 206.470 ;
        RECT 64.745 206.210 65.005 206.470 ;
        RECT 65.065 206.210 65.325 206.470 ;
        RECT 82.295 206.210 82.555 206.470 ;
        RECT 82.615 206.210 82.875 206.470 ;
        RECT 82.935 206.210 83.195 206.470 ;
        RECT 83.255 206.210 83.515 206.470 ;
        RECT 83.575 206.210 83.835 206.470 ;
        RECT 40.000 205.700 40.260 205.960 ;
        RECT 69.900 205.700 70.160 205.960 ;
        RECT 43.220 205.360 43.480 205.620 ;
        RECT 19.760 204.680 20.020 204.940 ;
        RECT 26.200 204.680 26.460 204.940 ;
        RECT 32.640 204.680 32.900 204.940 ;
        RECT 39.540 205.020 39.800 205.280 ;
        RECT 40.920 204.680 41.180 204.940 ;
        RECT 58.400 205.020 58.660 205.280 ;
        RECT 39.080 204.340 39.340 204.600 ;
        RECT 44.600 204.680 44.860 204.940 ;
        RECT 51.960 204.680 52.220 204.940 ;
        RECT 53.340 204.680 53.600 204.940 ;
        RECT 60.240 204.680 60.500 204.940 ;
        RECT 65.760 204.680 66.020 204.940 ;
        RECT 71.280 204.680 71.540 204.940 ;
        RECT 77.720 204.680 77.980 204.940 ;
        RECT 84.160 204.680 84.420 204.940 ;
        RECT 68.060 204.340 68.320 204.600 ;
        RECT 37.700 204.000 37.960 204.260 ;
        RECT 38.620 204.000 38.880 204.260 ;
        RECT 42.760 204.000 43.020 204.260 ;
        RECT 46.900 204.000 47.160 204.260 ;
        RECT 53.800 204.000 54.060 204.260 ;
        RECT 57.480 204.000 57.740 204.260 ;
        RECT 60.700 204.000 60.960 204.260 ;
        RECT 69.440 204.000 69.700 204.260 ;
        RECT 72.200 204.000 72.460 204.260 ;
        RECT 79.560 204.000 79.820 204.260 ;
        RECT 85.540 204.000 85.800 204.260 ;
        RECT 36.020 203.490 36.280 203.750 ;
        RECT 36.340 203.490 36.600 203.750 ;
        RECT 36.660 203.490 36.920 203.750 ;
        RECT 36.980 203.490 37.240 203.750 ;
        RECT 37.300 203.490 37.560 203.750 ;
        RECT 54.530 203.490 54.790 203.750 ;
        RECT 54.850 203.490 55.110 203.750 ;
        RECT 55.170 203.490 55.430 203.750 ;
        RECT 55.490 203.490 55.750 203.750 ;
        RECT 55.810 203.490 56.070 203.750 ;
        RECT 73.040 203.490 73.300 203.750 ;
        RECT 73.360 203.490 73.620 203.750 ;
        RECT 73.680 203.490 73.940 203.750 ;
        RECT 74.000 203.490 74.260 203.750 ;
        RECT 74.320 203.490 74.580 203.750 ;
        RECT 91.550 203.490 91.810 203.750 ;
        RECT 91.870 203.490 92.130 203.750 ;
        RECT 92.190 203.490 92.450 203.750 ;
        RECT 92.510 203.490 92.770 203.750 ;
        RECT 92.830 203.490 93.090 203.750 ;
        RECT 52.880 202.980 53.140 203.240 ;
        RECT 40.460 202.300 40.720 202.560 ;
        RECT 41.840 202.640 42.100 202.900 ;
        RECT 41.380 202.300 41.640 202.560 ;
        RECT 39.540 201.280 39.800 201.540 ;
        RECT 41.380 201.280 41.640 201.540 ;
        RECT 42.300 201.280 42.560 201.540 ;
        RECT 50.120 202.300 50.380 202.560 ;
        RECT 53.340 202.300 53.600 202.560 ;
        RECT 56.560 202.980 56.820 203.240 ;
        RECT 60.240 202.980 60.500 203.240 ;
        RECT 85.540 202.980 85.800 203.240 ;
        RECT 61.620 202.300 61.880 202.560 ;
        RECT 79.560 202.640 79.820 202.900 ;
        RECT 77.720 202.300 77.980 202.560 ;
        RECT 57.940 201.960 58.200 202.220 ;
        RECT 63.000 201.960 63.260 202.220 ;
        RECT 66.220 201.960 66.480 202.220 ;
        RECT 66.680 201.960 66.940 202.220 ;
        RECT 72.200 201.960 72.460 202.220 ;
        RECT 51.960 201.280 52.220 201.540 ;
        RECT 52.420 201.280 52.680 201.540 ;
        RECT 61.160 201.280 61.420 201.540 ;
        RECT 70.360 201.280 70.620 201.540 ;
        RECT 86.460 201.280 86.720 201.540 ;
        RECT 26.765 200.770 27.025 201.030 ;
        RECT 27.085 200.770 27.345 201.030 ;
        RECT 27.405 200.770 27.665 201.030 ;
        RECT 27.725 200.770 27.985 201.030 ;
        RECT 28.045 200.770 28.305 201.030 ;
        RECT 45.275 200.770 45.535 201.030 ;
        RECT 45.595 200.770 45.855 201.030 ;
        RECT 45.915 200.770 46.175 201.030 ;
        RECT 46.235 200.770 46.495 201.030 ;
        RECT 46.555 200.770 46.815 201.030 ;
        RECT 63.785 200.770 64.045 201.030 ;
        RECT 64.105 200.770 64.365 201.030 ;
        RECT 64.425 200.770 64.685 201.030 ;
        RECT 64.745 200.770 65.005 201.030 ;
        RECT 65.065 200.770 65.325 201.030 ;
        RECT 82.295 200.770 82.555 201.030 ;
        RECT 82.615 200.770 82.875 201.030 ;
        RECT 82.935 200.770 83.195 201.030 ;
        RECT 83.255 200.770 83.515 201.030 ;
        RECT 83.575 200.770 83.835 201.030 ;
        RECT 40.000 200.260 40.260 200.520 ;
        RECT 40.460 200.260 40.720 200.520 ;
        RECT 50.120 200.260 50.380 200.520 ;
        RECT 61.620 200.260 61.880 200.520 ;
        RECT 66.220 200.260 66.480 200.520 ;
        RECT 69.900 200.260 70.160 200.520 ;
        RECT 70.820 200.260 71.080 200.520 ;
        RECT 75.880 200.260 76.140 200.520 ;
        RECT 85.080 200.260 85.340 200.520 ;
        RECT 46.440 199.920 46.700 200.180 ;
        RECT 38.620 199.580 38.880 199.840 ;
        RECT 38.160 199.240 38.420 199.500 ;
        RECT 41.380 199.580 41.640 199.840 ;
        RECT 59.320 199.920 59.580 200.180 ;
        RECT 51.960 199.580 52.220 199.840 ;
        RECT 57.480 199.580 57.740 199.840 ;
        RECT 53.800 199.240 54.060 199.500 ;
        RECT 59.780 199.240 60.040 199.500 ;
        RECT 69.440 199.920 69.700 200.180 ;
        RECT 80.020 199.920 80.280 200.180 ;
        RECT 66.680 199.240 66.940 199.500 ;
        RECT 70.360 199.240 70.620 199.500 ;
        RECT 42.760 198.900 43.020 199.160 ;
        RECT 72.660 198.900 72.920 199.160 ;
        RECT 86.460 199.580 86.720 199.840 ;
        RECT 74.960 199.240 75.220 199.500 ;
        RECT 75.880 199.240 76.140 199.500 ;
        RECT 76.340 199.240 76.600 199.500 ;
        RECT 77.260 199.240 77.520 199.500 ;
        RECT 78.640 199.240 78.900 199.500 ;
        RECT 87.840 199.240 88.100 199.500 ;
        RECT 91.060 199.240 91.320 199.500 ;
        RECT 46.440 198.560 46.700 198.820 ;
        RECT 52.420 198.560 52.680 198.820 ;
        RECT 53.800 198.560 54.060 198.820 ;
        RECT 80.480 198.900 80.740 199.160 ;
        RECT 76.800 198.560 77.060 198.820 ;
        RECT 79.560 198.560 79.820 198.820 ;
        RECT 88.760 198.560 89.020 198.820 ;
        RECT 36.020 198.050 36.280 198.310 ;
        RECT 36.340 198.050 36.600 198.310 ;
        RECT 36.660 198.050 36.920 198.310 ;
        RECT 36.980 198.050 37.240 198.310 ;
        RECT 37.300 198.050 37.560 198.310 ;
        RECT 54.530 198.050 54.790 198.310 ;
        RECT 54.850 198.050 55.110 198.310 ;
        RECT 55.170 198.050 55.430 198.310 ;
        RECT 55.490 198.050 55.750 198.310 ;
        RECT 55.810 198.050 56.070 198.310 ;
        RECT 73.040 198.050 73.300 198.310 ;
        RECT 73.360 198.050 73.620 198.310 ;
        RECT 73.680 198.050 73.940 198.310 ;
        RECT 74.000 198.050 74.260 198.310 ;
        RECT 74.320 198.050 74.580 198.310 ;
        RECT 91.550 198.050 91.810 198.310 ;
        RECT 91.870 198.050 92.130 198.310 ;
        RECT 92.190 198.050 92.450 198.310 ;
        RECT 92.510 198.050 92.770 198.310 ;
        RECT 92.830 198.050 93.090 198.310 ;
        RECT 74.960 197.540 75.220 197.800 ;
        RECT 76.800 197.540 77.060 197.800 ;
        RECT 77.720 197.540 77.980 197.800 ;
        RECT 78.640 197.540 78.900 197.800 ;
        RECT 91.060 197.540 91.320 197.800 ;
        RECT 38.160 196.860 38.420 197.120 ;
        RECT 75.880 197.200 76.140 197.460 ;
        RECT 36.320 196.520 36.580 196.780 ;
        RECT 46.900 196.520 47.160 196.780 ;
        RECT 58.860 196.860 59.120 197.120 ;
        RECT 62.080 196.860 62.340 197.120 ;
        RECT 47.820 196.520 48.080 196.780 ;
        RECT 58.400 196.520 58.660 196.780 ;
        RECT 37.240 196.180 37.500 196.440 ;
        RECT 38.160 195.840 38.420 196.100 ;
        RECT 44.600 195.840 44.860 196.100 ;
        RECT 52.420 195.840 52.680 196.100 ;
        RECT 74.500 196.860 74.760 197.120 ;
        RECT 74.960 196.860 75.220 197.120 ;
        RECT 81.860 197.200 82.120 197.460 ;
        RECT 77.260 196.860 77.520 197.120 ;
        RECT 79.560 196.860 79.820 197.120 ;
        RECT 80.020 196.860 80.280 197.120 ;
        RECT 71.740 196.520 72.000 196.780 ;
        RECT 67.600 195.840 67.860 196.100 ;
        RECT 78.180 195.840 78.440 196.100 ;
        RECT 26.765 195.330 27.025 195.590 ;
        RECT 27.085 195.330 27.345 195.590 ;
        RECT 27.405 195.330 27.665 195.590 ;
        RECT 27.725 195.330 27.985 195.590 ;
        RECT 28.045 195.330 28.305 195.590 ;
        RECT 45.275 195.330 45.535 195.590 ;
        RECT 45.595 195.330 45.855 195.590 ;
        RECT 45.915 195.330 46.175 195.590 ;
        RECT 46.235 195.330 46.495 195.590 ;
        RECT 46.555 195.330 46.815 195.590 ;
        RECT 63.785 195.330 64.045 195.590 ;
        RECT 64.105 195.330 64.365 195.590 ;
        RECT 64.425 195.330 64.685 195.590 ;
        RECT 64.745 195.330 65.005 195.590 ;
        RECT 65.065 195.330 65.325 195.590 ;
        RECT 82.295 195.330 82.555 195.590 ;
        RECT 82.615 195.330 82.875 195.590 ;
        RECT 82.935 195.330 83.195 195.590 ;
        RECT 83.255 195.330 83.515 195.590 ;
        RECT 83.575 195.330 83.835 195.590 ;
        RECT 47.820 194.820 48.080 195.080 ;
        RECT 51.960 194.820 52.220 195.080 ;
        RECT 53.340 194.820 53.600 195.080 ;
        RECT 53.800 194.820 54.060 195.080 ;
        RECT 58.860 194.820 59.120 195.080 ;
        RECT 62.080 194.820 62.340 195.080 ;
        RECT 68.980 194.820 69.240 195.080 ;
        RECT 70.820 194.820 71.080 195.080 ;
        RECT 74.500 194.820 74.760 195.080 ;
        RECT 41.840 194.140 42.100 194.400 ;
        RECT 38.160 193.800 38.420 194.060 ;
        RECT 44.600 193.800 44.860 194.060 ;
        RECT 52.420 194.140 52.680 194.400 ;
        RECT 59.320 194.140 59.580 194.400 ;
        RECT 66.680 194.140 66.940 194.400 ;
        RECT 60.700 193.800 60.960 194.060 ;
        RECT 31.720 193.120 31.980 193.380 ;
        RECT 50.120 193.120 50.380 193.380 ;
        RECT 51.960 193.120 52.220 193.380 ;
        RECT 67.600 193.800 67.860 194.060 ;
        RECT 68.060 193.120 68.320 193.380 ;
        RECT 71.740 193.120 72.000 193.380 ;
        RECT 72.660 193.800 72.920 194.060 ;
        RECT 74.960 194.140 75.220 194.400 ;
        RECT 78.640 194.480 78.900 194.740 ;
        RECT 77.260 194.140 77.520 194.400 ;
        RECT 80.020 194.480 80.280 194.740 ;
        RECT 76.800 193.460 77.060 193.720 ;
        RECT 75.420 193.120 75.680 193.380 ;
        RECT 78.640 193.460 78.900 193.720 ;
        RECT 80.020 193.460 80.280 193.720 ;
        RECT 85.080 193.800 85.340 194.060 ;
        RECT 86.460 193.800 86.720 194.060 ;
        RECT 88.760 193.800 89.020 194.060 ;
        RECT 91.060 193.800 91.320 194.060 ;
        RECT 83.700 193.120 83.960 193.380 ;
        RECT 36.020 192.610 36.280 192.870 ;
        RECT 36.340 192.610 36.600 192.870 ;
        RECT 36.660 192.610 36.920 192.870 ;
        RECT 36.980 192.610 37.240 192.870 ;
        RECT 37.300 192.610 37.560 192.870 ;
        RECT 54.530 192.610 54.790 192.870 ;
        RECT 54.850 192.610 55.110 192.870 ;
        RECT 55.170 192.610 55.430 192.870 ;
        RECT 55.490 192.610 55.750 192.870 ;
        RECT 55.810 192.610 56.070 192.870 ;
        RECT 73.040 192.610 73.300 192.870 ;
        RECT 73.360 192.610 73.620 192.870 ;
        RECT 73.680 192.610 73.940 192.870 ;
        RECT 74.000 192.610 74.260 192.870 ;
        RECT 74.320 192.610 74.580 192.870 ;
        RECT 91.550 192.610 91.810 192.870 ;
        RECT 91.870 192.610 92.130 192.870 ;
        RECT 92.190 192.610 92.450 192.870 ;
        RECT 92.510 192.610 92.770 192.870 ;
        RECT 92.830 192.610 93.090 192.870 ;
        RECT 37.700 192.100 37.960 192.360 ;
        RECT 59.780 192.100 60.040 192.360 ;
        RECT 74.960 192.100 75.220 192.360 ;
        RECT 75.420 192.100 75.680 192.360 ;
        RECT 78.180 192.100 78.440 192.360 ;
        RECT 42.300 191.760 42.560 192.020 ;
        RECT 50.580 191.420 50.840 191.680 ;
        RECT 56.100 191.420 56.360 191.680 ;
        RECT 56.560 191.420 56.820 191.680 ;
        RECT 91.060 191.760 91.320 192.020 ;
        RECT 81.860 191.420 82.120 191.680 ;
        RECT 83.700 191.420 83.960 191.680 ;
        RECT 52.420 191.080 52.680 191.340 ;
        RECT 58.400 191.080 58.660 191.340 ;
        RECT 59.780 191.080 60.040 191.340 ;
        RECT 72.660 191.080 72.920 191.340 ;
        RECT 76.800 191.080 77.060 191.340 ;
        RECT 58.860 190.740 59.120 191.000 ;
        RECT 59.320 190.740 59.580 191.000 ;
        RECT 61.160 190.740 61.420 191.000 ;
        RECT 67.600 190.740 67.860 191.000 ;
        RECT 34.940 190.400 35.200 190.660 ;
        RECT 35.400 190.400 35.660 190.660 ;
        RECT 40.000 190.400 40.260 190.660 ;
        RECT 57.480 190.400 57.740 190.660 ;
        RECT 61.620 190.400 61.880 190.660 ;
        RECT 62.540 190.400 62.800 190.660 ;
        RECT 26.765 189.890 27.025 190.150 ;
        RECT 27.085 189.890 27.345 190.150 ;
        RECT 27.405 189.890 27.665 190.150 ;
        RECT 27.725 189.890 27.985 190.150 ;
        RECT 28.045 189.890 28.305 190.150 ;
        RECT 45.275 189.890 45.535 190.150 ;
        RECT 45.595 189.890 45.855 190.150 ;
        RECT 45.915 189.890 46.175 190.150 ;
        RECT 46.235 189.890 46.495 190.150 ;
        RECT 46.555 189.890 46.815 190.150 ;
        RECT 63.785 189.890 64.045 190.150 ;
        RECT 64.105 189.890 64.365 190.150 ;
        RECT 64.425 189.890 64.685 190.150 ;
        RECT 64.745 189.890 65.005 190.150 ;
        RECT 65.065 189.890 65.325 190.150 ;
        RECT 82.295 189.890 82.555 190.150 ;
        RECT 82.615 189.890 82.875 190.150 ;
        RECT 82.935 189.890 83.195 190.150 ;
        RECT 83.255 189.890 83.515 190.150 ;
        RECT 83.575 189.890 83.835 190.150 ;
        RECT 50.120 189.040 50.380 189.300 ;
        RECT 31.720 188.700 31.980 188.960 ;
        RECT 34.940 188.700 35.200 188.960 ;
        RECT 40.460 188.700 40.720 188.960 ;
        RECT 35.400 188.360 35.660 188.620 ;
        RECT 38.620 188.360 38.880 188.620 ;
        RECT 42.300 188.360 42.560 188.620 ;
        RECT 43.680 188.020 43.940 188.280 ;
        RECT 46.900 188.020 47.160 188.280 ;
        RECT 44.140 187.680 44.400 187.940 ;
        RECT 45.520 187.680 45.780 187.940 ;
        RECT 50.580 188.360 50.840 188.620 ;
        RECT 52.420 189.380 52.680 189.640 ;
        RECT 56.560 189.380 56.820 189.640 ;
        RECT 58.860 189.380 59.120 189.640 ;
        RECT 62.080 189.380 62.340 189.640 ;
        RECT 51.960 189.040 52.220 189.300 ;
        RECT 57.020 188.700 57.280 188.960 ;
        RECT 52.880 188.360 53.140 188.620 ;
        RECT 56.100 188.020 56.360 188.280 ;
        RECT 63.000 188.700 63.260 188.960 ;
        RECT 78.640 189.380 78.900 189.640 ;
        RECT 80.020 189.380 80.280 189.640 ;
        RECT 61.620 188.360 61.880 188.620 ;
        RECT 62.540 188.360 62.800 188.620 ;
        RECT 52.880 187.680 53.140 187.940 ;
        RECT 53.340 187.680 53.600 187.940 ;
        RECT 53.800 187.680 54.060 187.940 ;
        RECT 60.240 188.020 60.500 188.280 ;
        RECT 63.920 188.020 64.180 188.280 ;
        RECT 71.740 188.360 72.000 188.620 ;
        RECT 58.400 187.680 58.660 187.940 ;
        RECT 80.940 188.020 81.200 188.280 ;
        RECT 85.080 188.360 85.340 188.620 ;
        RECT 85.540 188.360 85.800 188.620 ;
        RECT 86.460 188.360 86.720 188.620 ;
        RECT 71.280 187.680 71.540 187.940 ;
        RECT 77.720 187.680 77.980 187.940 ;
        RECT 80.020 187.680 80.280 187.940 ;
        RECT 83.700 187.680 83.960 187.940 ;
        RECT 36.020 187.170 36.280 187.430 ;
        RECT 36.340 187.170 36.600 187.430 ;
        RECT 36.660 187.170 36.920 187.430 ;
        RECT 36.980 187.170 37.240 187.430 ;
        RECT 37.300 187.170 37.560 187.430 ;
        RECT 54.530 187.170 54.790 187.430 ;
        RECT 54.850 187.170 55.110 187.430 ;
        RECT 55.170 187.170 55.430 187.430 ;
        RECT 55.490 187.170 55.750 187.430 ;
        RECT 55.810 187.170 56.070 187.430 ;
        RECT 73.040 187.170 73.300 187.430 ;
        RECT 73.360 187.170 73.620 187.430 ;
        RECT 73.680 187.170 73.940 187.430 ;
        RECT 74.000 187.170 74.260 187.430 ;
        RECT 74.320 187.170 74.580 187.430 ;
        RECT 91.550 187.170 91.810 187.430 ;
        RECT 91.870 187.170 92.130 187.430 ;
        RECT 92.190 187.170 92.450 187.430 ;
        RECT 92.510 187.170 92.770 187.430 ;
        RECT 92.830 187.170 93.090 187.430 ;
        RECT 35.400 186.660 35.660 186.920 ;
        RECT 38.620 186.660 38.880 186.920 ;
        RECT 37.240 185.980 37.500 186.240 ;
        RECT 42.300 186.660 42.560 186.920 ;
        RECT 44.140 185.980 44.400 186.240 ;
        RECT 45.520 185.980 45.780 186.240 ;
        RECT 52.420 186.660 52.680 186.920 ;
        RECT 58.400 186.660 58.660 186.920 ;
        RECT 60.240 186.660 60.500 186.920 ;
        RECT 63.920 186.660 64.180 186.920 ;
        RECT 74.960 186.660 75.220 186.920 ;
        RECT 85.540 186.660 85.800 186.920 ;
        RECT 58.860 186.320 59.120 186.580 ;
        RECT 41.380 185.640 41.640 185.900 ;
        RECT 50.580 185.980 50.840 186.240 ;
        RECT 52.880 185.980 53.140 186.240 ;
        RECT 53.340 185.980 53.600 186.240 ;
        RECT 53.800 185.980 54.060 186.240 ;
        RECT 57.480 185.980 57.740 186.240 ;
        RECT 50.120 185.300 50.380 185.560 ;
        RECT 34.940 184.960 35.200 185.220 ;
        RECT 39.540 184.960 39.800 185.220 ;
        RECT 40.460 184.960 40.720 185.220 ;
        RECT 47.360 184.960 47.620 185.220 ;
        RECT 51.500 184.960 51.760 185.220 ;
        RECT 57.480 185.300 57.740 185.560 ;
        RECT 66.220 185.980 66.480 186.240 ;
        RECT 63.000 185.300 63.260 185.560 ;
        RECT 65.760 185.300 66.020 185.560 ;
        RECT 71.280 185.980 71.540 186.240 ;
        RECT 75.880 185.980 76.140 186.240 ;
        RECT 77.260 185.980 77.520 186.240 ;
        RECT 77.720 185.980 77.980 186.240 ;
        RECT 78.640 185.980 78.900 186.240 ;
        RECT 79.100 185.980 79.360 186.240 ;
        RECT 81.860 185.980 82.120 186.240 ;
        RECT 83.700 185.980 83.960 186.240 ;
        RECT 72.660 185.640 72.920 185.900 ;
        RECT 81.400 185.640 81.660 185.900 ;
        RECT 80.940 185.300 81.200 185.560 ;
        RECT 91.060 185.640 91.320 185.900 ;
        RECT 59.320 184.960 59.580 185.220 ;
        RECT 62.540 184.960 62.800 185.220 ;
        RECT 67.140 184.960 67.400 185.220 ;
        RECT 77.720 184.960 77.980 185.220 ;
        RECT 91.060 184.960 91.320 185.220 ;
        RECT 26.765 184.450 27.025 184.710 ;
        RECT 27.085 184.450 27.345 184.710 ;
        RECT 27.405 184.450 27.665 184.710 ;
        RECT 27.725 184.450 27.985 184.710 ;
        RECT 28.045 184.450 28.305 184.710 ;
        RECT 45.275 184.450 45.535 184.710 ;
        RECT 45.595 184.450 45.855 184.710 ;
        RECT 45.915 184.450 46.175 184.710 ;
        RECT 46.235 184.450 46.495 184.710 ;
        RECT 46.555 184.450 46.815 184.710 ;
        RECT 63.785 184.450 64.045 184.710 ;
        RECT 64.105 184.450 64.365 184.710 ;
        RECT 64.425 184.450 64.685 184.710 ;
        RECT 64.745 184.450 65.005 184.710 ;
        RECT 65.065 184.450 65.325 184.710 ;
        RECT 82.295 184.450 82.555 184.710 ;
        RECT 82.615 184.450 82.875 184.710 ;
        RECT 82.935 184.450 83.195 184.710 ;
        RECT 83.255 184.450 83.515 184.710 ;
        RECT 83.575 184.450 83.835 184.710 ;
        RECT 41.380 183.940 41.640 184.200 ;
        RECT 41.840 183.940 42.100 184.200 ;
        RECT 66.220 183.940 66.480 184.200 ;
        RECT 78.640 183.940 78.900 184.200 ;
        RECT 39.540 183.600 39.800 183.860 ;
        RECT 58.400 183.600 58.660 183.860 ;
        RECT 37.240 183.260 37.500 183.520 ;
        RECT 58.860 183.260 59.120 183.520 ;
        RECT 77.260 183.260 77.520 183.520 ;
        RECT 62.080 182.920 62.340 183.180 ;
        RECT 66.220 182.920 66.480 183.180 ;
        RECT 80.940 183.940 81.200 184.200 ;
        RECT 81.400 183.940 81.660 184.200 ;
        RECT 79.560 183.600 79.820 183.860 ;
        RECT 80.020 182.920 80.280 183.180 ;
        RECT 80.940 182.920 81.200 183.180 ;
        RECT 60.240 182.580 60.500 182.840 ;
        RECT 75.880 182.580 76.140 182.840 ;
        RECT 81.860 182.580 82.120 182.840 ;
        RECT 48.280 182.240 48.540 182.500 ;
        RECT 66.680 182.240 66.940 182.500 ;
        RECT 80.020 182.240 80.280 182.500 ;
        RECT 80.940 182.240 81.200 182.500 ;
        RECT 36.020 181.730 36.280 181.990 ;
        RECT 36.340 181.730 36.600 181.990 ;
        RECT 36.660 181.730 36.920 181.990 ;
        RECT 36.980 181.730 37.240 181.990 ;
        RECT 37.300 181.730 37.560 181.990 ;
        RECT 54.530 181.730 54.790 181.990 ;
        RECT 54.850 181.730 55.110 181.990 ;
        RECT 55.170 181.730 55.430 181.990 ;
        RECT 55.490 181.730 55.750 181.990 ;
        RECT 55.810 181.730 56.070 181.990 ;
        RECT 73.040 181.730 73.300 181.990 ;
        RECT 73.360 181.730 73.620 181.990 ;
        RECT 73.680 181.730 73.940 181.990 ;
        RECT 74.000 181.730 74.260 181.990 ;
        RECT 74.320 181.730 74.580 181.990 ;
        RECT 91.550 181.730 91.810 181.990 ;
        RECT 91.870 181.730 92.130 181.990 ;
        RECT 92.190 181.730 92.450 181.990 ;
        RECT 92.510 181.730 92.770 181.990 ;
        RECT 92.830 181.730 93.090 181.990 ;
        RECT 43.220 181.220 43.480 181.480 ;
        RECT 48.280 181.220 48.540 181.480 ;
        RECT 50.580 181.220 50.840 181.480 ;
        RECT 52.420 181.220 52.680 181.480 ;
        RECT 53.800 181.220 54.060 181.480 ;
        RECT 58.400 181.220 58.660 181.480 ;
        RECT 58.860 181.220 59.120 181.480 ;
        RECT 69.900 181.220 70.160 181.480 ;
        RECT 43.680 180.880 43.940 181.140 ;
        RECT 44.600 180.540 44.860 180.800 ;
        RECT 46.900 180.540 47.160 180.800 ;
        RECT 53.340 180.880 53.600 181.140 ;
        RECT 42.760 180.200 43.020 180.460 ;
        RECT 50.120 180.200 50.380 180.460 ;
        RECT 54.260 180.540 54.520 180.800 ;
        RECT 57.940 180.540 58.200 180.800 ;
        RECT 58.860 180.540 59.120 180.800 ;
        RECT 62.540 180.540 62.800 180.800 ;
        RECT 66.220 180.880 66.480 181.140 ;
        RECT 66.680 180.880 66.940 181.140 ;
        RECT 71.280 180.880 71.540 181.140 ;
        RECT 76.340 180.880 76.600 181.140 ;
        RECT 67.140 180.540 67.400 180.800 ;
        RECT 86.000 181.220 86.260 181.480 ;
        RECT 77.720 180.540 77.980 180.800 ;
        RECT 62.080 179.860 62.340 180.120 ;
        RECT 41.380 179.520 41.640 179.780 ;
        RECT 48.740 179.520 49.000 179.780 ;
        RECT 70.820 180.200 71.080 180.460 ;
        RECT 79.560 180.540 79.820 180.800 ;
        RECT 66.220 179.860 66.480 180.120 ;
        RECT 79.560 179.860 79.820 180.120 ;
        RECT 65.760 179.520 66.020 179.780 ;
        RECT 77.720 179.520 77.980 179.780 ;
        RECT 81.400 179.860 81.660 180.120 ;
        RECT 82.780 180.540 83.040 180.800 ;
        RECT 82.320 180.200 82.580 180.460 ;
        RECT 91.060 179.520 91.320 179.780 ;
        RECT 26.765 179.010 27.025 179.270 ;
        RECT 27.085 179.010 27.345 179.270 ;
        RECT 27.405 179.010 27.665 179.270 ;
        RECT 27.725 179.010 27.985 179.270 ;
        RECT 28.045 179.010 28.305 179.270 ;
        RECT 45.275 179.010 45.535 179.270 ;
        RECT 45.595 179.010 45.855 179.270 ;
        RECT 45.915 179.010 46.175 179.270 ;
        RECT 46.235 179.010 46.495 179.270 ;
        RECT 46.555 179.010 46.815 179.270 ;
        RECT 63.785 179.010 64.045 179.270 ;
        RECT 64.105 179.010 64.365 179.270 ;
        RECT 64.425 179.010 64.685 179.270 ;
        RECT 64.745 179.010 65.005 179.270 ;
        RECT 65.065 179.010 65.325 179.270 ;
        RECT 82.295 179.010 82.555 179.270 ;
        RECT 82.615 179.010 82.875 179.270 ;
        RECT 82.935 179.010 83.195 179.270 ;
        RECT 83.255 179.010 83.515 179.270 ;
        RECT 83.575 179.010 83.835 179.270 ;
        RECT 41.840 178.500 42.100 178.760 ;
        RECT 44.600 178.500 44.860 178.760 ;
        RECT 53.340 178.500 53.600 178.760 ;
        RECT 54.260 178.500 54.520 178.760 ;
        RECT 57.940 178.500 58.200 178.760 ;
        RECT 58.400 178.500 58.660 178.760 ;
        RECT 58.860 178.500 59.120 178.760 ;
        RECT 71.740 178.500 72.000 178.760 ;
        RECT 46.900 178.160 47.160 178.420 ;
        RECT 69.900 178.160 70.160 178.420 ;
        RECT 78.640 178.160 78.900 178.420 ;
        RECT 58.400 177.820 58.660 178.080 ;
        RECT 75.880 177.820 76.140 178.080 ;
        RECT 41.380 177.480 41.640 177.740 ;
        RECT 50.580 177.480 50.840 177.740 ;
        RECT 51.960 177.480 52.220 177.740 ;
        RECT 52.420 177.480 52.680 177.740 ;
        RECT 66.220 177.480 66.480 177.740 ;
        RECT 69.440 177.480 69.700 177.740 ;
        RECT 69.900 177.480 70.160 177.740 ;
        RECT 71.280 177.480 71.540 177.740 ;
        RECT 77.720 177.480 77.980 177.740 ;
        RECT 78.640 177.480 78.900 177.740 ;
        RECT 81.400 178.500 81.660 178.760 ;
        RECT 79.560 177.480 79.820 177.740 ;
        RECT 57.020 177.140 57.280 177.400 ;
        RECT 60.700 177.140 60.960 177.400 ;
        RECT 47.820 176.800 48.080 177.060 ;
        RECT 50.120 176.800 50.380 177.060 ;
        RECT 52.880 176.800 53.140 177.060 ;
        RECT 61.160 176.800 61.420 177.060 ;
        RECT 62.540 176.800 62.800 177.060 ;
        RECT 69.900 176.800 70.160 177.060 ;
        RECT 70.360 176.800 70.620 177.060 ;
        RECT 81.400 177.480 81.660 177.740 ;
        RECT 85.080 177.480 85.340 177.740 ;
        RECT 86.000 177.480 86.260 177.740 ;
        RECT 90.140 177.480 90.400 177.740 ;
        RECT 81.400 176.800 81.660 177.060 ;
        RECT 83.700 176.800 83.960 177.060 ;
        RECT 36.020 176.290 36.280 176.550 ;
        RECT 36.340 176.290 36.600 176.550 ;
        RECT 36.660 176.290 36.920 176.550 ;
        RECT 36.980 176.290 37.240 176.550 ;
        RECT 37.300 176.290 37.560 176.550 ;
        RECT 54.530 176.290 54.790 176.550 ;
        RECT 54.850 176.290 55.110 176.550 ;
        RECT 55.170 176.290 55.430 176.550 ;
        RECT 55.490 176.290 55.750 176.550 ;
        RECT 55.810 176.290 56.070 176.550 ;
        RECT 73.040 176.290 73.300 176.550 ;
        RECT 73.360 176.290 73.620 176.550 ;
        RECT 73.680 176.290 73.940 176.550 ;
        RECT 74.000 176.290 74.260 176.550 ;
        RECT 74.320 176.290 74.580 176.550 ;
        RECT 91.550 176.290 91.810 176.550 ;
        RECT 91.870 176.290 92.130 176.550 ;
        RECT 92.190 176.290 92.450 176.550 ;
        RECT 92.510 176.290 92.770 176.550 ;
        RECT 92.830 176.290 93.090 176.550 ;
        RECT 41.840 175.780 42.100 176.040 ;
        RECT 42.760 175.780 43.020 176.040 ;
        RECT 47.820 175.440 48.080 175.700 ;
        RECT 51.040 175.780 51.300 176.040 ;
        RECT 56.560 175.780 56.820 176.040 ;
        RECT 48.280 175.100 48.540 175.360 ;
        RECT 50.120 175.440 50.380 175.700 ;
        RECT 73.120 175.780 73.380 176.040 ;
        RECT 46.900 174.420 47.160 174.680 ;
        RECT 48.740 174.420 49.000 174.680 ;
        RECT 52.880 175.100 53.140 175.360 ;
        RECT 53.340 175.100 53.600 175.360 ;
        RECT 58.400 175.100 58.660 175.360 ;
        RECT 70.360 175.100 70.620 175.360 ;
        RECT 74.040 175.780 74.300 176.040 ;
        RECT 90.600 175.780 90.860 176.040 ;
        RECT 76.340 175.440 76.600 175.700 ;
        RECT 78.640 175.440 78.900 175.700 ;
        RECT 81.860 175.440 82.120 175.700 ;
        RECT 75.420 175.100 75.680 175.360 ;
        RECT 78.180 175.100 78.440 175.360 ;
        RECT 83.700 175.100 83.960 175.360 ;
        RECT 85.080 175.100 85.340 175.360 ;
        RECT 50.580 174.760 50.840 175.020 ;
        RECT 68.980 174.760 69.240 175.020 ;
        RECT 71.280 174.760 71.540 175.020 ;
        RECT 73.120 174.760 73.380 175.020 ;
        RECT 74.040 174.760 74.300 175.020 ;
        RECT 44.600 174.080 44.860 174.340 ;
        RECT 49.200 174.080 49.460 174.340 ;
        RECT 60.240 174.080 60.500 174.340 ;
        RECT 74.040 174.080 74.300 174.340 ;
        RECT 74.500 174.080 74.760 174.340 ;
        RECT 90.600 174.080 90.860 174.340 ;
        RECT 26.765 173.570 27.025 173.830 ;
        RECT 27.085 173.570 27.345 173.830 ;
        RECT 27.405 173.570 27.665 173.830 ;
        RECT 27.725 173.570 27.985 173.830 ;
        RECT 28.045 173.570 28.305 173.830 ;
        RECT 45.275 173.570 45.535 173.830 ;
        RECT 45.595 173.570 45.855 173.830 ;
        RECT 45.915 173.570 46.175 173.830 ;
        RECT 46.235 173.570 46.495 173.830 ;
        RECT 46.555 173.570 46.815 173.830 ;
        RECT 63.785 173.570 64.045 173.830 ;
        RECT 64.105 173.570 64.365 173.830 ;
        RECT 64.425 173.570 64.685 173.830 ;
        RECT 64.745 173.570 65.005 173.830 ;
        RECT 65.065 173.570 65.325 173.830 ;
        RECT 82.295 173.570 82.555 173.830 ;
        RECT 82.615 173.570 82.875 173.830 ;
        RECT 82.935 173.570 83.195 173.830 ;
        RECT 83.255 173.570 83.515 173.830 ;
        RECT 83.575 173.570 83.835 173.830 ;
        RECT 46.900 173.060 47.160 173.320 ;
        RECT 48.280 173.060 48.540 173.320 ;
        RECT 52.880 173.060 53.140 173.320 ;
        RECT 48.740 172.720 49.000 172.980 ;
        RECT 51.960 172.720 52.220 172.980 ;
        RECT 74.500 173.060 74.760 173.320 ;
        RECT 75.420 173.060 75.680 173.320 ;
        RECT 38.160 172.040 38.420 172.300 ;
        RECT 44.600 172.040 44.860 172.300 ;
        RECT 58.860 172.380 59.120 172.640 ;
        RECT 69.900 172.720 70.160 172.980 ;
        RECT 72.660 172.720 72.920 172.980 ;
        RECT 47.360 172.040 47.620 172.300 ;
        RECT 51.500 172.040 51.760 172.300 ;
        RECT 57.020 172.040 57.280 172.300 ;
        RECT 58.400 172.040 58.660 172.300 ;
        RECT 42.300 171.360 42.560 171.620 ;
        RECT 45.060 171.360 45.320 171.620 ;
        RECT 45.980 171.360 46.240 171.620 ;
        RECT 52.420 171.360 52.680 171.620 ;
        RECT 52.880 171.360 53.140 171.620 ;
        RECT 58.860 171.700 59.120 171.960 ;
        RECT 61.160 172.040 61.420 172.300 ;
        RECT 79.560 173.060 79.820 173.320 ;
        RECT 81.400 173.060 81.660 173.320 ;
        RECT 69.440 172.040 69.700 172.300 ;
        RECT 78.180 172.380 78.440 172.640 ;
        RECT 90.600 172.380 90.860 172.640 ;
        RECT 63.920 171.700 64.180 171.960 ;
        RECT 60.700 171.360 60.960 171.620 ;
        RECT 72.660 171.360 72.920 171.620 ;
        RECT 74.040 172.040 74.300 172.300 ;
        RECT 85.080 172.040 85.340 172.300 ;
        RECT 91.060 172.040 91.320 172.300 ;
        RECT 78.640 171.360 78.900 171.620 ;
        RECT 79.560 171.360 79.820 171.620 ;
        RECT 81.400 171.360 81.660 171.620 ;
        RECT 83.700 171.360 83.960 171.620 ;
        RECT 36.020 170.850 36.280 171.110 ;
        RECT 36.340 170.850 36.600 171.110 ;
        RECT 36.660 170.850 36.920 171.110 ;
        RECT 36.980 170.850 37.240 171.110 ;
        RECT 37.300 170.850 37.560 171.110 ;
        RECT 54.530 170.850 54.790 171.110 ;
        RECT 54.850 170.850 55.110 171.110 ;
        RECT 55.170 170.850 55.430 171.110 ;
        RECT 55.490 170.850 55.750 171.110 ;
        RECT 55.810 170.850 56.070 171.110 ;
        RECT 73.040 170.850 73.300 171.110 ;
        RECT 73.360 170.850 73.620 171.110 ;
        RECT 73.680 170.850 73.940 171.110 ;
        RECT 74.000 170.850 74.260 171.110 ;
        RECT 74.320 170.850 74.580 171.110 ;
        RECT 91.550 170.850 91.810 171.110 ;
        RECT 91.870 170.850 92.130 171.110 ;
        RECT 92.190 170.850 92.450 171.110 ;
        RECT 92.510 170.850 92.770 171.110 ;
        RECT 92.830 170.850 93.090 171.110 ;
        RECT 38.160 170.340 38.420 170.600 ;
        RECT 40.460 169.660 40.720 169.920 ;
        RECT 42.300 169.660 42.560 169.920 ;
        RECT 44.140 169.660 44.400 169.920 ;
        RECT 45.060 170.000 45.320 170.260 ;
        RECT 49.200 170.000 49.460 170.260 ;
        RECT 45.980 169.660 46.240 169.920 ;
        RECT 47.360 169.660 47.620 169.920 ;
        RECT 47.820 169.660 48.080 169.920 ;
        RECT 53.340 170.340 53.600 170.600 ;
        RECT 57.480 170.340 57.740 170.600 ;
        RECT 60.700 170.340 60.960 170.600 ;
        RECT 63.920 170.340 64.180 170.600 ;
        RECT 50.580 170.000 50.840 170.260 ;
        RECT 38.160 168.640 38.420 168.900 ;
        RECT 44.140 168.980 44.400 169.240 ;
        RECT 59.780 169.660 60.040 169.920 ;
        RECT 71.740 170.000 72.000 170.260 ;
        RECT 67.600 169.660 67.860 169.920 ;
        RECT 72.660 169.660 72.920 169.920 ;
        RECT 60.700 169.320 60.960 169.580 ;
        RECT 62.080 169.320 62.340 169.580 ;
        RECT 72.200 169.320 72.460 169.580 ;
        RECT 76.800 169.660 77.060 169.920 ;
        RECT 79.560 169.660 79.820 169.920 ;
        RECT 83.700 169.660 83.960 169.920 ;
        RECT 81.860 169.320 82.120 169.580 ;
        RECT 62.540 168.980 62.800 169.240 ;
        RECT 51.960 168.640 52.220 168.900 ;
        RECT 76.340 168.640 76.600 168.900 ;
        RECT 91.060 168.640 91.320 168.900 ;
        RECT 26.765 168.130 27.025 168.390 ;
        RECT 27.085 168.130 27.345 168.390 ;
        RECT 27.405 168.130 27.665 168.390 ;
        RECT 27.725 168.130 27.985 168.390 ;
        RECT 28.045 168.130 28.305 168.390 ;
        RECT 45.275 168.130 45.535 168.390 ;
        RECT 45.595 168.130 45.855 168.390 ;
        RECT 45.915 168.130 46.175 168.390 ;
        RECT 46.235 168.130 46.495 168.390 ;
        RECT 46.555 168.130 46.815 168.390 ;
        RECT 63.785 168.130 64.045 168.390 ;
        RECT 64.105 168.130 64.365 168.390 ;
        RECT 64.425 168.130 64.685 168.390 ;
        RECT 64.745 168.130 65.005 168.390 ;
        RECT 65.065 168.130 65.325 168.390 ;
        RECT 82.295 168.130 82.555 168.390 ;
        RECT 82.615 168.130 82.875 168.390 ;
        RECT 82.935 168.130 83.195 168.390 ;
        RECT 83.255 168.130 83.515 168.390 ;
        RECT 83.575 168.130 83.835 168.390 ;
        RECT 61.160 167.620 61.420 167.880 ;
        RECT 80.940 167.280 81.200 167.540 ;
        RECT 51.960 166.940 52.220 167.200 ;
        RECT 53.800 166.600 54.060 166.860 ;
        RECT 57.020 166.940 57.280 167.200 ;
        RECT 67.600 166.940 67.860 167.200 ;
        RECT 68.060 166.940 68.320 167.200 ;
        RECT 56.560 166.600 56.820 166.860 ;
        RECT 59.780 166.600 60.040 166.860 ;
        RECT 75.880 166.600 76.140 166.860 ;
        RECT 78.640 166.940 78.900 167.200 ;
        RECT 76.800 166.600 77.060 166.860 ;
        RECT 57.020 166.260 57.280 166.520 ;
        RECT 59.320 166.260 59.580 166.520 ;
        RECT 66.680 166.260 66.940 166.520 ;
        RECT 46.900 165.920 47.160 166.180 ;
        RECT 48.740 165.920 49.000 166.180 ;
        RECT 57.480 165.920 57.740 166.180 ;
        RECT 68.060 165.920 68.320 166.180 ;
        RECT 78.640 166.260 78.900 166.520 ;
        RECT 81.400 166.600 81.660 166.860 ;
        RECT 90.140 166.600 90.400 166.860 ;
        RECT 36.020 165.410 36.280 165.670 ;
        RECT 36.340 165.410 36.600 165.670 ;
        RECT 36.660 165.410 36.920 165.670 ;
        RECT 36.980 165.410 37.240 165.670 ;
        RECT 37.300 165.410 37.560 165.670 ;
        RECT 54.530 165.410 54.790 165.670 ;
        RECT 54.850 165.410 55.110 165.670 ;
        RECT 55.170 165.410 55.430 165.670 ;
        RECT 55.490 165.410 55.750 165.670 ;
        RECT 55.810 165.410 56.070 165.670 ;
        RECT 73.040 165.410 73.300 165.670 ;
        RECT 73.360 165.410 73.620 165.670 ;
        RECT 73.680 165.410 73.940 165.670 ;
        RECT 74.000 165.410 74.260 165.670 ;
        RECT 74.320 165.410 74.580 165.670 ;
        RECT 91.550 165.410 91.810 165.670 ;
        RECT 91.870 165.410 92.130 165.670 ;
        RECT 92.190 165.410 92.450 165.670 ;
        RECT 92.510 165.410 92.770 165.670 ;
        RECT 92.830 165.410 93.090 165.670 ;
        RECT 47.820 164.900 48.080 165.160 ;
        RECT 53.800 164.900 54.060 165.160 ;
        RECT 57.020 164.900 57.280 165.160 ;
        RECT 57.480 164.900 57.740 165.160 ;
        RECT 42.760 164.220 43.020 164.480 ;
        RECT 50.580 164.560 50.840 164.820 ;
        RECT 46.900 164.220 47.160 164.480 ;
        RECT 47.820 164.220 48.080 164.480 ;
        RECT 56.560 164.560 56.820 164.820 ;
        RECT 47.360 163.880 47.620 164.140 ;
        RECT 53.800 164.220 54.060 164.480 ;
        RECT 37.700 163.200 37.960 163.460 ;
        RECT 59.780 164.900 60.040 165.160 ;
        RECT 74.040 164.900 74.300 165.160 ;
        RECT 75.880 164.900 76.140 165.160 ;
        RECT 63.000 164.220 63.260 164.480 ;
        RECT 77.720 164.560 77.980 164.820 ;
        RECT 66.680 164.220 66.940 164.480 ;
        RECT 68.060 164.220 68.320 164.480 ;
        RECT 68.520 164.220 68.780 164.480 ;
        RECT 69.440 164.220 69.700 164.480 ;
        RECT 78.640 164.220 78.900 164.480 ;
        RECT 85.080 164.900 85.340 165.160 ;
        RECT 81.860 164.560 82.120 164.820 ;
        RECT 80.940 164.220 81.200 164.480 ;
        RECT 86.000 164.220 86.260 164.480 ;
        RECT 60.700 163.540 60.960 163.800 ;
        RECT 84.160 163.880 84.420 164.140 ;
        RECT 79.560 163.540 79.820 163.800 ;
        RECT 58.400 163.200 58.660 163.460 ;
        RECT 78.180 163.200 78.440 163.460 ;
        RECT 81.400 163.200 81.660 163.460 ;
        RECT 87.840 163.540 88.100 163.800 ;
        RECT 90.600 163.200 90.860 163.460 ;
        RECT 26.765 162.690 27.025 162.950 ;
        RECT 27.085 162.690 27.345 162.950 ;
        RECT 27.405 162.690 27.665 162.950 ;
        RECT 27.725 162.690 27.985 162.950 ;
        RECT 28.045 162.690 28.305 162.950 ;
        RECT 45.275 162.690 45.535 162.950 ;
        RECT 45.595 162.690 45.855 162.950 ;
        RECT 45.915 162.690 46.175 162.950 ;
        RECT 46.235 162.690 46.495 162.950 ;
        RECT 46.555 162.690 46.815 162.950 ;
        RECT 63.785 162.690 64.045 162.950 ;
        RECT 64.105 162.690 64.365 162.950 ;
        RECT 64.425 162.690 64.685 162.950 ;
        RECT 64.745 162.690 65.005 162.950 ;
        RECT 65.065 162.690 65.325 162.950 ;
        RECT 82.295 162.690 82.555 162.950 ;
        RECT 82.615 162.690 82.875 162.950 ;
        RECT 82.935 162.690 83.195 162.950 ;
        RECT 83.255 162.690 83.515 162.950 ;
        RECT 83.575 162.690 83.835 162.950 ;
        RECT 47.820 162.180 48.080 162.440 ;
        RECT 63.000 162.180 63.260 162.440 ;
        RECT 68.520 162.180 68.780 162.440 ;
        RECT 52.880 161.840 53.140 162.100 ;
        RECT 53.340 161.840 53.600 162.100 ;
        RECT 84.160 162.180 84.420 162.440 ;
        RECT 37.700 160.820 37.960 161.080 ;
        RECT 50.580 161.160 50.840 161.420 ;
        RECT 50.120 160.820 50.380 161.080 ;
        RECT 74.960 161.500 75.220 161.760 ;
        RECT 58.400 161.160 58.660 161.420 ;
        RECT 38.160 160.480 38.420 160.740 ;
        RECT 51.960 160.480 52.220 160.740 ;
        RECT 56.560 160.820 56.820 161.080 ;
        RECT 68.060 160.820 68.320 161.080 ;
        RECT 68.980 160.820 69.240 161.080 ;
        RECT 76.340 161.160 76.600 161.420 ;
        RECT 80.480 161.840 80.740 162.100 ;
        RECT 72.200 160.820 72.460 161.080 ;
        RECT 74.040 160.820 74.300 161.080 ;
        RECT 54.260 160.480 54.520 160.740 ;
        RECT 69.900 160.480 70.160 160.740 ;
        RECT 74.960 160.480 75.220 160.740 ;
        RECT 78.180 161.160 78.440 161.420 ;
        RECT 80.020 161.160 80.280 161.420 ;
        RECT 80.940 161.160 81.200 161.420 ;
        RECT 81.400 161.160 81.660 161.420 ;
        RECT 85.080 161.160 85.340 161.420 ;
        RECT 36.020 159.970 36.280 160.230 ;
        RECT 36.340 159.970 36.600 160.230 ;
        RECT 36.660 159.970 36.920 160.230 ;
        RECT 36.980 159.970 37.240 160.230 ;
        RECT 37.300 159.970 37.560 160.230 ;
        RECT 54.530 159.970 54.790 160.230 ;
        RECT 54.850 159.970 55.110 160.230 ;
        RECT 55.170 159.970 55.430 160.230 ;
        RECT 55.490 159.970 55.750 160.230 ;
        RECT 55.810 159.970 56.070 160.230 ;
        RECT 73.040 159.970 73.300 160.230 ;
        RECT 73.360 159.970 73.620 160.230 ;
        RECT 73.680 159.970 73.940 160.230 ;
        RECT 74.000 159.970 74.260 160.230 ;
        RECT 74.320 159.970 74.580 160.230 ;
        RECT 91.550 159.970 91.810 160.230 ;
        RECT 91.870 159.970 92.130 160.230 ;
        RECT 92.190 159.970 92.450 160.230 ;
        RECT 92.510 159.970 92.770 160.230 ;
        RECT 92.830 159.970 93.090 160.230 ;
        RECT 69.440 159.460 69.700 159.720 ;
        RECT 75.420 159.460 75.680 159.720 ;
        RECT 60.240 159.120 60.500 159.380 ;
        RECT 43.220 158.780 43.480 159.040 ;
        RECT 52.420 158.780 52.680 159.040 ;
        RECT 56.560 158.780 56.820 159.040 ;
        RECT 55.640 158.440 55.900 158.700 ;
        RECT 80.480 158.440 80.740 158.700 ;
        RECT 81.860 158.440 82.120 158.700 ;
        RECT 38.160 157.760 38.420 158.020 ;
        RECT 47.360 158.100 47.620 158.360 ;
        RECT 50.120 157.760 50.380 158.020 ;
        RECT 56.560 157.760 56.820 158.020 ;
        RECT 69.900 157.760 70.160 158.020 ;
        RECT 75.880 157.760 76.140 158.020 ;
        RECT 87.840 157.760 88.100 158.020 ;
        RECT 26.765 157.250 27.025 157.510 ;
        RECT 27.085 157.250 27.345 157.510 ;
        RECT 27.405 157.250 27.665 157.510 ;
        RECT 27.725 157.250 27.985 157.510 ;
        RECT 28.045 157.250 28.305 157.510 ;
        RECT 45.275 157.250 45.535 157.510 ;
        RECT 45.595 157.250 45.855 157.510 ;
        RECT 45.915 157.250 46.175 157.510 ;
        RECT 46.235 157.250 46.495 157.510 ;
        RECT 46.555 157.250 46.815 157.510 ;
        RECT 63.785 157.250 64.045 157.510 ;
        RECT 64.105 157.250 64.365 157.510 ;
        RECT 64.425 157.250 64.685 157.510 ;
        RECT 64.745 157.250 65.005 157.510 ;
        RECT 65.065 157.250 65.325 157.510 ;
        RECT 82.295 157.250 82.555 157.510 ;
        RECT 82.615 157.250 82.875 157.510 ;
        RECT 82.935 157.250 83.195 157.510 ;
        RECT 83.255 157.250 83.515 157.510 ;
        RECT 83.575 157.250 83.835 157.510 ;
        RECT 43.220 156.740 43.480 157.000 ;
        RECT 56.560 156.400 56.820 156.660 ;
        RECT 72.200 156.740 72.460 157.000 ;
        RECT 77.720 156.740 77.980 157.000 ;
        RECT 50.120 156.060 50.380 156.320 ;
        RECT 55.640 156.060 55.900 156.320 ;
        RECT 43.680 155.720 43.940 155.980 ;
        RECT 44.600 155.720 44.860 155.980 ;
        RECT 45.520 155.720 45.780 155.980 ;
        RECT 57.020 155.720 57.280 155.980 ;
        RECT 54.260 155.380 54.520 155.640 ;
        RECT 48.280 155.040 48.540 155.300 ;
        RECT 51.960 155.040 52.220 155.300 ;
        RECT 52.880 155.040 53.140 155.300 ;
        RECT 53.800 155.040 54.060 155.300 ;
        RECT 67.600 155.720 67.860 155.980 ;
        RECT 68.520 156.060 68.780 156.320 ;
        RECT 68.980 155.720 69.240 155.980 ;
        RECT 69.440 155.720 69.700 155.980 ;
        RECT 75.880 156.060 76.140 156.320 ;
        RECT 74.960 155.720 75.220 155.980 ;
        RECT 71.740 155.380 72.000 155.640 ;
        RECT 77.260 155.720 77.520 155.980 ;
        RECT 77.720 155.720 77.980 155.980 ;
        RECT 65.300 155.040 65.560 155.300 ;
        RECT 65.760 155.040 66.020 155.300 ;
        RECT 72.660 155.040 72.920 155.300 ;
        RECT 74.960 155.040 75.220 155.300 ;
        RECT 82.320 155.380 82.580 155.640 ;
        RECT 36.020 154.530 36.280 154.790 ;
        RECT 36.340 154.530 36.600 154.790 ;
        RECT 36.660 154.530 36.920 154.790 ;
        RECT 36.980 154.530 37.240 154.790 ;
        RECT 37.300 154.530 37.560 154.790 ;
        RECT 54.530 154.530 54.790 154.790 ;
        RECT 54.850 154.530 55.110 154.790 ;
        RECT 55.170 154.530 55.430 154.790 ;
        RECT 55.490 154.530 55.750 154.790 ;
        RECT 55.810 154.530 56.070 154.790 ;
        RECT 73.040 154.530 73.300 154.790 ;
        RECT 73.360 154.530 73.620 154.790 ;
        RECT 73.680 154.530 73.940 154.790 ;
        RECT 74.000 154.530 74.260 154.790 ;
        RECT 74.320 154.530 74.580 154.790 ;
        RECT 91.550 154.530 91.810 154.790 ;
        RECT 91.870 154.530 92.130 154.790 ;
        RECT 92.190 154.530 92.450 154.790 ;
        RECT 92.510 154.530 92.770 154.790 ;
        RECT 92.830 154.530 93.090 154.790 ;
        RECT 45.520 154.020 45.780 154.280 ;
        RECT 48.280 154.020 48.540 154.280 ;
        RECT 53.340 154.020 53.600 154.280 ;
        RECT 53.800 154.020 54.060 154.280 ;
        RECT 57.020 154.020 57.280 154.280 ;
        RECT 46.900 153.680 47.160 153.940 ;
        RECT 40.460 153.340 40.720 153.600 ;
        RECT 42.300 153.340 42.560 153.600 ;
        RECT 41.840 152.320 42.100 152.580 ;
        RECT 47.360 153.340 47.620 153.600 ;
        RECT 48.740 153.340 49.000 153.600 ;
        RECT 54.720 153.680 54.980 153.940 ;
        RECT 52.420 153.340 52.680 153.600 ;
        RECT 51.960 153.000 52.220 153.260 ;
        RECT 53.340 153.340 53.600 153.600 ;
        RECT 52.880 152.660 53.140 152.920 ;
        RECT 51.500 152.320 51.760 152.580 ;
        RECT 55.180 153.340 55.440 153.600 ;
        RECT 65.760 153.340 66.020 153.600 ;
        RECT 69.900 154.020 70.160 154.280 ;
        RECT 71.740 154.020 72.000 154.280 ;
        RECT 72.200 154.020 72.460 154.280 ;
        RECT 77.260 154.020 77.520 154.280 ;
        RECT 82.320 154.020 82.580 154.280 ;
        RECT 74.500 153.680 74.760 153.940 ;
        RECT 56.100 153.000 56.360 153.260 ;
        RECT 72.200 153.340 72.460 153.600 ;
        RECT 72.660 153.340 72.920 153.600 ;
        RECT 75.420 153.340 75.680 153.600 ;
        RECT 68.980 152.660 69.240 152.920 ;
        RECT 69.440 152.660 69.700 152.920 ;
        RECT 73.120 152.660 73.380 152.920 ;
        RECT 63.000 152.320 63.260 152.580 ;
        RECT 71.740 152.320 72.000 152.580 ;
        RECT 26.765 151.810 27.025 152.070 ;
        RECT 27.085 151.810 27.345 152.070 ;
        RECT 27.405 151.810 27.665 152.070 ;
        RECT 27.725 151.810 27.985 152.070 ;
        RECT 28.045 151.810 28.305 152.070 ;
        RECT 45.275 151.810 45.535 152.070 ;
        RECT 45.595 151.810 45.855 152.070 ;
        RECT 45.915 151.810 46.175 152.070 ;
        RECT 46.235 151.810 46.495 152.070 ;
        RECT 46.555 151.810 46.815 152.070 ;
        RECT 63.785 151.810 64.045 152.070 ;
        RECT 64.105 151.810 64.365 152.070 ;
        RECT 64.425 151.810 64.685 152.070 ;
        RECT 64.745 151.810 65.005 152.070 ;
        RECT 65.065 151.810 65.325 152.070 ;
        RECT 82.295 151.810 82.555 152.070 ;
        RECT 82.615 151.810 82.875 152.070 ;
        RECT 82.935 151.810 83.195 152.070 ;
        RECT 83.255 151.810 83.515 152.070 ;
        RECT 83.575 151.810 83.835 152.070 ;
        RECT 42.300 151.300 42.560 151.560 ;
        RECT 46.900 151.300 47.160 151.560 ;
        RECT 52.880 151.300 53.140 151.560 ;
        RECT 72.200 151.300 72.460 151.560 ;
        RECT 74.500 151.300 74.760 151.560 ;
        RECT 74.960 151.300 75.220 151.560 ;
        RECT 59.320 150.960 59.580 151.220 ;
        RECT 60.240 150.960 60.500 151.220 ;
        RECT 56.100 150.620 56.360 150.880 ;
        RECT 41.840 150.280 42.100 150.540 ;
        RECT 44.140 150.280 44.400 150.540 ;
        RECT 48.740 149.940 49.000 150.200 ;
        RECT 38.160 149.600 38.420 149.860 ;
        RECT 55.180 150.280 55.440 150.540 ;
        RECT 56.560 150.280 56.820 150.540 ;
        RECT 53.800 149.940 54.060 150.200 ;
        RECT 54.720 149.940 54.980 150.200 ;
        RECT 61.620 150.280 61.880 150.540 ;
        RECT 63.000 150.280 63.260 150.540 ;
        RECT 67.600 150.280 67.860 150.540 ;
        RECT 68.060 150.280 68.320 150.540 ;
        RECT 71.740 150.280 72.000 150.540 ;
        RECT 74.960 150.280 75.220 150.540 ;
        RECT 80.020 150.280 80.280 150.540 ;
        RECT 59.320 149.940 59.580 150.200 ;
        RECT 53.340 149.600 53.600 149.860 ;
        RECT 61.160 149.600 61.420 149.860 ;
        RECT 62.540 149.600 62.800 149.860 ;
        RECT 72.200 149.600 72.460 149.860 ;
        RECT 36.020 149.090 36.280 149.350 ;
        RECT 36.340 149.090 36.600 149.350 ;
        RECT 36.660 149.090 36.920 149.350 ;
        RECT 36.980 149.090 37.240 149.350 ;
        RECT 37.300 149.090 37.560 149.350 ;
        RECT 54.530 149.090 54.790 149.350 ;
        RECT 54.850 149.090 55.110 149.350 ;
        RECT 55.170 149.090 55.430 149.350 ;
        RECT 55.490 149.090 55.750 149.350 ;
        RECT 55.810 149.090 56.070 149.350 ;
        RECT 73.040 149.090 73.300 149.350 ;
        RECT 73.360 149.090 73.620 149.350 ;
        RECT 73.680 149.090 73.940 149.350 ;
        RECT 74.000 149.090 74.260 149.350 ;
        RECT 74.320 149.090 74.580 149.350 ;
        RECT 91.550 149.090 91.810 149.350 ;
        RECT 91.870 149.090 92.130 149.350 ;
        RECT 92.190 149.090 92.450 149.350 ;
        RECT 92.510 149.090 92.770 149.350 ;
        RECT 92.830 149.090 93.090 149.350 ;
        RECT 53.340 148.580 53.600 148.840 ;
        RECT 61.160 148.580 61.420 148.840 ;
        RECT 61.620 148.580 61.880 148.840 ;
        RECT 66.680 148.580 66.940 148.840 ;
        RECT 55.180 148.240 55.440 148.500 ;
        RECT 54.260 147.560 54.520 147.820 ;
        RECT 48.740 147.220 49.000 147.480 ;
        RECT 61.160 147.900 61.420 148.160 ;
        RECT 62.540 147.900 62.800 148.160 ;
        RECT 68.060 148.240 68.320 148.500 ;
        RECT 71.740 148.580 72.000 148.840 ;
        RECT 74.960 148.580 75.220 148.840 ;
        RECT 72.200 147.900 72.460 148.160 ;
        RECT 59.320 147.560 59.580 147.820 ;
        RECT 60.700 147.220 60.960 147.480 ;
        RECT 53.340 146.880 53.600 147.140 ;
        RECT 57.020 146.880 57.280 147.140 ;
        RECT 70.360 146.880 70.620 147.140 ;
        RECT 131.200 147.000 131.805 147.605 ;
        RECT 26.765 146.370 27.025 146.630 ;
        RECT 27.085 146.370 27.345 146.630 ;
        RECT 27.405 146.370 27.665 146.630 ;
        RECT 27.725 146.370 27.985 146.630 ;
        RECT 28.045 146.370 28.305 146.630 ;
        RECT 45.275 146.370 45.535 146.630 ;
        RECT 45.595 146.370 45.855 146.630 ;
        RECT 45.915 146.370 46.175 146.630 ;
        RECT 46.235 146.370 46.495 146.630 ;
        RECT 46.555 146.370 46.815 146.630 ;
        RECT 63.785 146.370 64.045 146.630 ;
        RECT 64.105 146.370 64.365 146.630 ;
        RECT 64.425 146.370 64.685 146.630 ;
        RECT 64.745 146.370 65.005 146.630 ;
        RECT 65.065 146.370 65.325 146.630 ;
        RECT 82.295 146.370 82.555 146.630 ;
        RECT 82.615 146.370 82.875 146.630 ;
        RECT 82.935 146.370 83.195 146.630 ;
        RECT 83.255 146.370 83.515 146.630 ;
        RECT 83.575 146.370 83.835 146.630 ;
        RECT 53.800 145.860 54.060 146.120 ;
        RECT 59.320 145.860 59.580 146.120 ;
        RECT 71.740 145.860 72.000 146.120 ;
        RECT 38.160 145.180 38.420 145.440 ;
        RECT 55.180 145.180 55.440 145.440 ;
        RECT 75.420 145.180 75.680 145.440 ;
        RECT 113.200 145.800 113.800 146.400 ;
        RECT 116.400 145.900 117.000 146.500 ;
        RECT 119.300 146.000 119.900 146.600 ;
        RECT 48.740 144.840 49.000 145.100 ;
        RECT 53.340 144.840 53.600 145.100 ;
        RECT 45.060 144.500 45.320 144.760 ;
        RECT 50.120 144.160 50.380 144.420 ;
        RECT 56.560 144.840 56.820 145.100 ;
        RECT 60.240 144.840 60.500 145.100 ;
        RECT 122.300 145.900 122.900 146.500 ;
        RECT 125.300 145.900 125.900 146.500 ;
        RECT 128.300 145.900 128.900 146.500 ;
        RECT 67.140 144.500 67.400 144.760 ;
        RECT 36.020 143.650 36.280 143.910 ;
        RECT 36.340 143.650 36.600 143.910 ;
        RECT 36.660 143.650 36.920 143.910 ;
        RECT 36.980 143.650 37.240 143.910 ;
        RECT 37.300 143.650 37.560 143.910 ;
        RECT 54.530 143.650 54.790 143.910 ;
        RECT 54.850 143.650 55.110 143.910 ;
        RECT 55.170 143.650 55.430 143.910 ;
        RECT 55.490 143.650 55.750 143.910 ;
        RECT 55.810 143.650 56.070 143.910 ;
        RECT 73.040 143.650 73.300 143.910 ;
        RECT 73.360 143.650 73.620 143.910 ;
        RECT 73.680 143.650 73.940 143.910 ;
        RECT 74.000 143.650 74.260 143.910 ;
        RECT 74.320 143.650 74.580 143.910 ;
        RECT 91.550 143.650 91.810 143.910 ;
        RECT 91.870 143.650 92.130 143.910 ;
        RECT 92.190 143.650 92.450 143.910 ;
        RECT 92.510 143.650 92.770 143.910 ;
        RECT 92.830 143.650 93.090 143.910 ;
        RECT 45.060 143.140 45.320 143.400 ;
        RECT 67.140 143.140 67.400 143.400 ;
        RECT 44.600 142.460 44.860 142.720 ;
        RECT 50.120 142.460 50.380 142.720 ;
        RECT 66.680 142.460 66.940 142.720 ;
        RECT 70.360 142.460 70.620 142.720 ;
        RECT 26.765 140.930 27.025 141.190 ;
        RECT 27.085 140.930 27.345 141.190 ;
        RECT 27.405 140.930 27.665 141.190 ;
        RECT 27.725 140.930 27.985 141.190 ;
        RECT 28.045 140.930 28.305 141.190 ;
        RECT 45.275 140.930 45.535 141.190 ;
        RECT 45.595 140.930 45.855 141.190 ;
        RECT 45.915 140.930 46.175 141.190 ;
        RECT 46.235 140.930 46.495 141.190 ;
        RECT 46.555 140.930 46.815 141.190 ;
        RECT 63.785 140.930 64.045 141.190 ;
        RECT 64.105 140.930 64.365 141.190 ;
        RECT 64.425 140.930 64.685 141.190 ;
        RECT 64.745 140.930 65.005 141.190 ;
        RECT 65.065 140.930 65.325 141.190 ;
        RECT 82.295 140.930 82.555 141.190 ;
        RECT 82.615 140.930 82.875 141.190 ;
        RECT 82.935 140.930 83.195 141.190 ;
        RECT 83.255 140.930 83.515 141.190 ;
        RECT 83.575 140.930 83.835 141.190 ;
        RECT 36.020 138.210 36.280 138.470 ;
        RECT 36.340 138.210 36.600 138.470 ;
        RECT 36.660 138.210 36.920 138.470 ;
        RECT 36.980 138.210 37.240 138.470 ;
        RECT 37.300 138.210 37.560 138.470 ;
        RECT 54.530 138.210 54.790 138.470 ;
        RECT 54.850 138.210 55.110 138.470 ;
        RECT 55.170 138.210 55.430 138.470 ;
        RECT 55.490 138.210 55.750 138.470 ;
        RECT 55.810 138.210 56.070 138.470 ;
        RECT 73.040 138.210 73.300 138.470 ;
        RECT 73.360 138.210 73.620 138.470 ;
        RECT 73.680 138.210 73.940 138.470 ;
        RECT 74.000 138.210 74.260 138.470 ;
        RECT 74.320 138.210 74.580 138.470 ;
        RECT 91.550 138.210 91.810 138.470 ;
        RECT 91.870 138.210 92.130 138.470 ;
        RECT 92.190 138.210 92.450 138.470 ;
        RECT 92.510 138.210 92.770 138.470 ;
        RECT 92.830 138.210 93.090 138.470 ;
        RECT 26.765 135.490 27.025 135.750 ;
        RECT 27.085 135.490 27.345 135.750 ;
        RECT 27.405 135.490 27.665 135.750 ;
        RECT 27.725 135.490 27.985 135.750 ;
        RECT 28.045 135.490 28.305 135.750 ;
        RECT 45.275 135.490 45.535 135.750 ;
        RECT 45.595 135.490 45.855 135.750 ;
        RECT 45.915 135.490 46.175 135.750 ;
        RECT 46.235 135.490 46.495 135.750 ;
        RECT 46.555 135.490 46.815 135.750 ;
        RECT 63.785 135.490 64.045 135.750 ;
        RECT 64.105 135.490 64.365 135.750 ;
        RECT 64.425 135.490 64.685 135.750 ;
        RECT 64.745 135.490 65.005 135.750 ;
        RECT 65.065 135.490 65.325 135.750 ;
        RECT 82.295 135.490 82.555 135.750 ;
        RECT 82.615 135.490 82.875 135.750 ;
        RECT 82.935 135.490 83.195 135.750 ;
        RECT 83.255 135.490 83.515 135.750 ;
        RECT 83.575 135.490 83.835 135.750 ;
        RECT 36.020 132.770 36.280 133.030 ;
        RECT 36.340 132.770 36.600 133.030 ;
        RECT 36.660 132.770 36.920 133.030 ;
        RECT 36.980 132.770 37.240 133.030 ;
        RECT 37.300 132.770 37.560 133.030 ;
        RECT 54.530 132.770 54.790 133.030 ;
        RECT 54.850 132.770 55.110 133.030 ;
        RECT 55.170 132.770 55.430 133.030 ;
        RECT 55.490 132.770 55.750 133.030 ;
        RECT 55.810 132.770 56.070 133.030 ;
        RECT 73.040 132.770 73.300 133.030 ;
        RECT 73.360 132.770 73.620 133.030 ;
        RECT 73.680 132.770 73.940 133.030 ;
        RECT 74.000 132.770 74.260 133.030 ;
        RECT 74.320 132.770 74.580 133.030 ;
        RECT 91.550 132.770 91.810 133.030 ;
        RECT 91.870 132.770 92.130 133.030 ;
        RECT 92.190 132.770 92.450 133.030 ;
        RECT 92.510 132.770 92.770 133.030 ;
        RECT 92.830 132.770 93.090 133.030 ;
        RECT 103.000 77.700 104.000 78.700 ;
        RECT 137.900 35.700 138.500 36.300 ;
      LAYER met2 ;
        RECT 19.740 222.345 20.040 222.735 ;
        RECT 19.750 208.180 20.030 222.345 ;
        RECT 26.250 221.695 26.550 221.705 ;
        RECT 26.215 221.415 26.585 221.695 ;
        RECT 26.250 210.180 26.550 221.415 ;
        RECT 32.575 220.445 32.965 220.745 ;
        RECT 26.190 208.515 26.550 210.180 ;
        RECT 26.190 208.180 26.470 208.515 ;
        RECT 32.630 208.180 32.910 220.445 ;
        RECT 39.045 219.655 39.345 219.665 ;
        RECT 39.010 219.375 39.380 219.655 ;
        RECT 39.045 210.180 39.345 219.375 ;
        RECT 45.480 218.500 45.760 218.535 ;
        RECT 45.470 210.180 45.770 218.500 ;
        RECT 51.940 216.915 52.240 217.305 ;
        RECT 39.045 208.635 39.350 210.180 ;
        RECT 45.470 209.075 45.790 210.180 ;
        RECT 39.070 208.180 39.350 208.635 ;
        RECT 45.510 208.180 45.790 209.075 ;
        RECT 51.950 208.180 52.230 216.915 ;
        RECT 58.400 216.010 58.700 216.020 ;
        RECT 58.365 215.730 58.735 216.010 ;
        RECT 58.400 210.180 58.700 215.730 ;
        RECT 64.820 214.715 65.120 215.105 ;
        RECT 58.390 208.835 58.700 210.180 ;
        RECT 58.390 208.180 58.670 208.835 ;
        RECT 64.830 208.180 65.110 214.715 ;
        RECT 71.210 213.930 71.510 213.940 ;
        RECT 71.175 213.650 71.545 213.930 ;
        RECT 71.210 210.180 71.510 213.650 ;
        RECT 77.700 212.625 78.000 213.015 ;
        RECT 71.210 208.795 71.550 210.180 ;
        RECT 71.270 208.180 71.550 208.795 ;
        RECT 77.710 208.180 77.990 212.625 ;
        RECT 84.130 211.985 84.430 211.995 ;
        RECT 84.095 211.705 84.465 211.985 ;
        RECT 84.130 209.175 84.430 211.705 ;
        RECT 90.535 210.720 90.925 211.020 ;
        RECT 84.150 208.180 84.430 209.175 ;
        RECT 90.590 208.180 90.870 210.720 ;
        RECT 19.820 204.970 19.960 208.180 ;
        RECT 26.260 204.970 26.400 208.180 ;
        RECT 26.765 206.155 28.305 206.525 ;
        RECT 32.700 204.970 32.840 208.180 ;
        RECT 19.760 204.650 20.020 204.970 ;
        RECT 26.200 204.650 26.460 204.970 ;
        RECT 32.640 204.650 32.900 204.970 ;
        RECT 39.140 204.630 39.280 208.180 ;
        RECT 45.580 207.430 45.720 208.180 ;
        RECT 44.660 207.290 45.720 207.430 ;
        RECT 40.000 205.670 40.260 205.990 ;
        RECT 39.540 204.990 39.800 205.310 ;
        RECT 39.080 204.310 39.340 204.630 ;
        RECT 37.700 203.970 37.960 204.290 ;
        RECT 38.620 203.970 38.880 204.290 ;
        RECT 36.020 203.435 37.560 203.805 ;
        RECT 26.765 200.715 28.305 201.085 ;
        RECT 36.020 197.995 37.560 198.365 ;
        RECT 37.760 197.740 37.900 203.970 ;
        RECT 38.680 199.870 38.820 203.970 ;
        RECT 39.600 201.570 39.740 204.990 ;
        RECT 39.540 201.250 39.800 201.570 ;
        RECT 38.620 199.550 38.880 199.870 ;
        RECT 38.160 199.210 38.420 199.530 ;
        RECT 37.300 197.600 37.900 197.740 ;
        RECT 36.320 196.490 36.580 196.810 ;
        RECT 26.765 195.275 28.305 195.645 ;
        RECT 36.380 194.510 36.520 196.490 ;
        RECT 37.300 196.470 37.440 197.600 ;
        RECT 38.220 197.150 38.360 199.210 ;
        RECT 38.160 196.830 38.420 197.150 ;
        RECT 37.240 196.150 37.500 196.470 ;
        RECT 38.160 195.810 38.420 196.130 ;
        RECT 36.380 194.370 37.900 194.510 ;
        RECT 31.720 193.090 31.980 193.410 ;
        RECT 26.765 189.835 28.305 190.205 ;
        RECT 31.780 188.990 31.920 193.090 ;
        RECT 36.020 192.555 37.560 192.925 ;
        RECT 37.760 192.390 37.900 194.370 ;
        RECT 38.220 194.090 38.360 195.810 ;
        RECT 38.160 193.770 38.420 194.090 ;
        RECT 37.700 192.070 37.960 192.390 ;
        RECT 34.940 190.370 35.200 190.690 ;
        RECT 35.400 190.370 35.660 190.690 ;
        RECT 35.000 188.990 35.140 190.370 ;
        RECT 31.720 188.670 31.980 188.990 ;
        RECT 34.940 188.670 35.200 188.990 ;
        RECT 35.000 185.250 35.140 188.670 ;
        RECT 35.460 188.650 35.600 190.370 ;
        RECT 35.400 188.330 35.660 188.650 ;
        RECT 38.620 188.330 38.880 188.650 ;
        RECT 35.460 186.950 35.600 188.330 ;
        RECT 36.020 187.115 37.560 187.485 ;
        RECT 38.680 186.950 38.820 188.330 ;
        RECT 35.400 186.630 35.660 186.950 ;
        RECT 38.620 186.630 38.880 186.950 ;
        RECT 37.240 185.950 37.500 186.270 ;
        RECT 34.940 184.930 35.200 185.250 ;
        RECT 26.765 184.395 28.305 184.765 ;
        RECT 37.300 183.550 37.440 185.950 ;
        RECT 39.600 185.250 39.740 201.250 ;
        RECT 40.060 200.550 40.200 205.670 ;
        RECT 43.220 205.330 43.480 205.650 ;
        RECT 40.920 204.880 41.180 204.970 ;
        RECT 40.920 204.740 41.580 204.880 ;
        RECT 40.920 204.650 41.180 204.740 ;
        RECT 41.440 202.590 41.580 204.740 ;
        RECT 42.760 203.970 43.020 204.290 ;
        RECT 41.840 202.610 42.100 202.930 ;
        RECT 40.460 202.270 40.720 202.590 ;
        RECT 41.380 202.270 41.640 202.590 ;
        RECT 40.520 200.550 40.660 202.270 ;
        RECT 41.380 201.250 41.640 201.570 ;
        RECT 40.000 200.230 40.260 200.550 ;
        RECT 40.460 200.230 40.720 200.550 ;
        RECT 40.060 190.690 40.200 200.230 ;
        RECT 41.440 199.870 41.580 201.250 ;
        RECT 41.380 199.550 41.640 199.870 ;
        RECT 41.900 194.430 42.040 202.610 ;
        RECT 42.300 201.250 42.560 201.570 ;
        RECT 41.840 194.110 42.100 194.430 ;
        RECT 40.000 190.370 40.260 190.690 ;
        RECT 40.460 188.670 40.720 188.990 ;
        RECT 40.520 185.250 40.660 188.670 ;
        RECT 41.380 185.610 41.640 185.930 ;
        RECT 39.540 184.930 39.800 185.250 ;
        RECT 40.460 184.930 40.720 185.250 ;
        RECT 39.600 183.890 39.740 184.930 ;
        RECT 41.440 184.230 41.580 185.610 ;
        RECT 41.900 184.230 42.040 194.110 ;
        RECT 42.360 192.050 42.500 201.250 ;
        RECT 42.820 199.190 42.960 203.970 ;
        RECT 42.760 198.870 43.020 199.190 ;
        RECT 42.300 191.730 42.560 192.050 ;
        RECT 42.300 188.330 42.560 188.650 ;
        RECT 42.360 186.950 42.500 188.330 ;
        RECT 42.300 186.630 42.560 186.950 ;
        RECT 41.380 183.910 41.640 184.230 ;
        RECT 41.840 183.910 42.100 184.230 ;
        RECT 39.540 183.570 39.800 183.890 ;
        RECT 37.240 183.230 37.500 183.550 ;
        RECT 36.020 181.675 37.560 182.045 ;
        RECT 41.380 179.490 41.640 179.810 ;
        RECT 26.765 178.955 28.305 179.325 ;
        RECT 41.440 177.770 41.580 179.490 ;
        RECT 41.900 178.790 42.040 183.910 ;
        RECT 43.280 181.510 43.420 205.330 ;
        RECT 44.660 204.970 44.800 207.290 ;
        RECT 45.275 206.155 46.815 206.525 ;
        RECT 52.020 204.970 52.160 208.180 ;
        RECT 58.460 205.310 58.600 208.180 ;
        RECT 64.900 207.430 65.040 208.180 ;
        RECT 64.900 207.290 65.960 207.430 ;
        RECT 63.785 206.155 65.325 206.525 ;
        RECT 58.400 204.990 58.660 205.310 ;
        RECT 65.820 204.970 65.960 207.290 ;
        RECT 69.900 205.670 70.160 205.990 ;
        RECT 44.600 204.650 44.860 204.970 ;
        RECT 51.960 204.650 52.220 204.970 ;
        RECT 53.340 204.650 53.600 204.970 ;
        RECT 60.240 204.650 60.500 204.970 ;
        RECT 65.760 204.650 66.020 204.970 ;
        RECT 46.900 203.970 47.160 204.290 ;
        RECT 45.275 200.715 46.815 201.085 ;
        RECT 46.440 199.890 46.700 200.210 ;
        RECT 46.500 198.850 46.640 199.890 ;
        RECT 46.440 198.530 46.700 198.850 ;
        RECT 46.960 196.810 47.100 203.970 ;
        RECT 52.880 202.950 53.140 203.270 ;
        RECT 50.120 202.270 50.380 202.590 ;
        RECT 50.180 200.550 50.320 202.270 ;
        RECT 51.960 201.250 52.220 201.570 ;
        RECT 52.420 201.250 52.680 201.570 ;
        RECT 50.120 200.230 50.380 200.550 ;
        RECT 52.020 199.870 52.160 201.250 ;
        RECT 51.960 199.550 52.220 199.870 ;
        RECT 52.480 198.850 52.620 201.250 ;
        RECT 52.420 198.530 52.680 198.850 ;
        RECT 46.900 196.490 47.160 196.810 ;
        RECT 47.820 196.490 48.080 196.810 ;
        RECT 44.600 195.810 44.860 196.130 ;
        RECT 44.660 194.090 44.800 195.810 ;
        RECT 45.275 195.275 46.815 195.645 ;
        RECT 47.880 195.110 48.020 196.490 ;
        RECT 52.420 195.810 52.680 196.130 ;
        RECT 47.820 194.790 48.080 195.110 ;
        RECT 51.960 194.790 52.220 195.110 ;
        RECT 44.600 193.770 44.860 194.090 ;
        RECT 52.020 193.410 52.160 194.790 ;
        RECT 52.480 194.430 52.620 195.810 ;
        RECT 52.420 194.110 52.680 194.430 ;
        RECT 50.120 193.090 50.380 193.410 ;
        RECT 51.960 193.090 52.220 193.410 ;
        RECT 45.275 189.835 46.815 190.205 ;
        RECT 50.180 189.330 50.320 193.090 ;
        RECT 50.580 191.390 50.840 191.710 ;
        RECT 50.120 189.010 50.380 189.330 ;
        RECT 43.680 187.990 43.940 188.310 ;
        RECT 46.900 187.990 47.160 188.310 ;
        RECT 43.220 181.190 43.480 181.510 ;
        RECT 43.740 181.170 43.880 187.990 ;
        RECT 44.140 187.650 44.400 187.970 ;
        RECT 45.520 187.650 45.780 187.970 ;
        RECT 44.200 186.270 44.340 187.650 ;
        RECT 45.580 186.270 45.720 187.650 ;
        RECT 44.140 185.950 44.400 186.270 ;
        RECT 45.520 185.950 45.780 186.270 ;
        RECT 45.275 184.395 46.815 184.765 ;
        RECT 43.680 180.850 43.940 181.170 ;
        RECT 46.960 180.830 47.100 187.990 ;
        RECT 50.180 185.590 50.320 189.010 ;
        RECT 50.640 188.650 50.780 191.390 ;
        RECT 52.020 189.330 52.160 193.090 ;
        RECT 52.480 191.370 52.620 194.110 ;
        RECT 52.420 191.050 52.680 191.370 ;
        RECT 52.480 189.670 52.620 191.050 ;
        RECT 52.420 189.350 52.680 189.670 ;
        RECT 51.960 189.010 52.220 189.330 ;
        RECT 52.940 188.650 53.080 202.950 ;
        RECT 53.400 202.590 53.540 204.650 ;
        RECT 53.800 203.970 54.060 204.290 ;
        RECT 57.480 203.970 57.740 204.290 ;
        RECT 53.340 202.270 53.600 202.590 ;
        RECT 53.400 195.110 53.540 202.270 ;
        RECT 53.860 199.530 54.000 203.970 ;
        RECT 54.530 203.435 56.070 203.805 ;
        RECT 56.560 202.950 56.820 203.270 ;
        RECT 53.800 199.210 54.060 199.530 ;
        RECT 53.800 198.530 54.060 198.850 ;
        RECT 53.860 195.110 54.000 198.530 ;
        RECT 54.530 197.995 56.070 198.365 ;
        RECT 53.340 194.790 53.600 195.110 ;
        RECT 53.800 194.790 54.060 195.110 ;
        RECT 54.530 192.555 56.070 192.925 ;
        RECT 56.620 191.710 56.760 202.950 ;
        RECT 57.540 199.870 57.680 203.970 ;
        RECT 60.300 203.270 60.440 204.650 ;
        RECT 68.060 204.310 68.320 204.630 ;
        RECT 60.700 203.970 60.960 204.290 ;
        RECT 60.240 202.950 60.500 203.270 ;
        RECT 57.940 201.930 58.200 202.250 ;
        RECT 58.000 199.950 58.140 201.930 ;
        RECT 57.480 199.550 57.740 199.870 ;
        RECT 58.000 199.810 58.600 199.950 ;
        RECT 59.320 199.890 59.580 200.210 ;
        RECT 58.460 196.810 58.600 199.810 ;
        RECT 58.860 196.830 59.120 197.150 ;
        RECT 58.400 196.490 58.660 196.810 ;
        RECT 58.920 195.110 59.060 196.830 ;
        RECT 58.860 194.790 59.120 195.110 ;
        RECT 59.380 194.430 59.520 199.890 ;
        RECT 59.780 199.210 60.040 199.530 ;
        RECT 59.320 194.110 59.580 194.430 ;
        RECT 59.840 192.390 59.980 199.210 ;
        RECT 60.760 194.090 60.900 203.970 ;
        RECT 61.620 202.270 61.880 202.590 ;
        RECT 61.160 201.250 61.420 201.570 ;
        RECT 60.700 193.770 60.960 194.090 ;
        RECT 59.780 192.070 60.040 192.390 ;
        RECT 56.100 191.390 56.360 191.710 ;
        RECT 56.560 191.390 56.820 191.710 ;
        RECT 50.580 188.560 50.840 188.650 ;
        RECT 52.880 188.560 53.140 188.650 ;
        RECT 50.580 188.420 51.240 188.560 ;
        RECT 50.580 188.330 50.840 188.420 ;
        RECT 50.580 185.950 50.840 186.270 ;
        RECT 50.120 185.270 50.380 185.590 ;
        RECT 47.360 184.930 47.620 185.250 ;
        RECT 44.600 180.510 44.860 180.830 ;
        RECT 46.900 180.510 47.160 180.830 ;
        RECT 42.760 180.170 43.020 180.490 ;
        RECT 41.840 178.470 42.100 178.790 ;
        RECT 41.380 177.450 41.640 177.770 ;
        RECT 36.020 176.235 37.560 176.605 ;
        RECT 41.900 176.070 42.040 178.470 ;
        RECT 42.820 176.070 42.960 180.170 ;
        RECT 44.660 178.790 44.800 180.510 ;
        RECT 45.275 178.955 46.815 179.325 ;
        RECT 44.600 178.470 44.860 178.790 ;
        RECT 46.960 178.450 47.100 180.510 ;
        RECT 46.900 178.130 47.160 178.450 ;
        RECT 41.840 175.750 42.100 176.070 ;
        RECT 42.760 175.750 43.020 176.070 ;
        RECT 26.765 173.515 28.305 173.885 ;
        RECT 38.160 172.010 38.420 172.330 ;
        RECT 36.020 170.795 37.560 171.165 ;
        RECT 38.220 170.630 38.360 172.010 ;
        RECT 42.300 171.330 42.560 171.650 ;
        RECT 38.160 170.310 38.420 170.630 ;
        RECT 42.360 169.950 42.500 171.330 ;
        RECT 40.460 169.630 40.720 169.950 ;
        RECT 42.300 169.630 42.560 169.950 ;
        RECT 38.160 168.610 38.420 168.930 ;
        RECT 26.765 168.075 28.305 168.445 ;
        RECT 36.020 165.355 37.560 165.725 ;
        RECT 37.700 163.170 37.960 163.490 ;
        RECT 26.765 162.635 28.305 163.005 ;
        RECT 37.760 161.110 37.900 163.170 ;
        RECT 37.700 160.790 37.960 161.110 ;
        RECT 38.220 160.770 38.360 168.610 ;
        RECT 38.160 160.450 38.420 160.770 ;
        RECT 36.020 159.915 37.560 160.285 ;
        RECT 38.220 158.050 38.360 160.450 ;
        RECT 38.160 157.730 38.420 158.050 ;
        RECT 26.765 157.195 28.305 157.565 ;
        RECT 36.020 154.475 37.560 154.845 ;
        RECT 26.765 151.755 28.305 152.125 ;
        RECT 38.220 149.890 38.360 157.730 ;
        RECT 40.520 153.630 40.660 169.630 ;
        RECT 42.820 164.510 42.960 175.750 ;
        RECT 46.900 174.390 47.160 174.710 ;
        RECT 44.600 174.050 44.860 174.370 ;
        RECT 44.660 172.330 44.800 174.050 ;
        RECT 45.275 173.515 46.815 173.885 ;
        RECT 46.960 173.350 47.100 174.390 ;
        RECT 46.900 173.030 47.160 173.350 ;
        RECT 47.420 172.330 47.560 184.930 ;
        RECT 48.280 182.210 48.540 182.530 ;
        RECT 48.340 181.510 48.480 182.210 ;
        RECT 50.640 181.510 50.780 185.950 ;
        RECT 48.280 181.190 48.540 181.510 ;
        RECT 50.580 181.190 50.840 181.510 ;
        RECT 50.120 180.170 50.380 180.490 ;
        RECT 48.740 179.490 49.000 179.810 ;
        RECT 47.820 176.770 48.080 177.090 ;
        RECT 47.880 175.730 48.020 176.770 ;
        RECT 47.820 175.410 48.080 175.730 ;
        RECT 44.600 172.010 44.860 172.330 ;
        RECT 47.360 172.010 47.620 172.330 ;
        RECT 45.060 171.330 45.320 171.650 ;
        RECT 45.980 171.330 46.240 171.650 ;
        RECT 47.880 171.390 48.020 175.410 ;
        RECT 48.280 175.070 48.540 175.390 ;
        RECT 48.340 173.350 48.480 175.070 ;
        RECT 48.800 174.710 48.940 179.490 ;
        RECT 50.180 177.090 50.320 180.170 ;
        RECT 50.580 177.450 50.840 177.770 ;
        RECT 50.120 176.770 50.380 177.090 ;
        RECT 50.180 175.730 50.320 176.770 ;
        RECT 50.120 175.410 50.380 175.730 ;
        RECT 50.640 175.050 50.780 177.450 ;
        RECT 51.100 176.070 51.240 188.420 ;
        RECT 52.480 188.420 53.140 188.560 ;
        RECT 52.480 186.950 52.620 188.420 ;
        RECT 52.880 188.330 53.140 188.420 ;
        RECT 56.160 188.390 56.300 191.390 ;
        RECT 56.620 189.670 56.760 191.390 ;
        RECT 58.400 191.050 58.660 191.370 ;
        RECT 59.780 191.050 60.040 191.370 ;
        RECT 57.480 190.370 57.740 190.690 ;
        RECT 56.560 189.350 56.820 189.670 ;
        RECT 57.020 188.670 57.280 188.990 ;
        RECT 56.160 188.310 56.760 188.390 ;
        RECT 56.100 188.250 56.760 188.310 ;
        RECT 56.100 187.990 56.360 188.250 ;
        RECT 52.880 187.650 53.140 187.970 ;
        RECT 53.340 187.650 53.600 187.970 ;
        RECT 53.800 187.650 54.060 187.970 ;
        RECT 52.420 186.630 52.680 186.950 ;
        RECT 52.940 186.270 53.080 187.650 ;
        RECT 53.400 186.270 53.540 187.650 ;
        RECT 53.860 186.270 54.000 187.650 ;
        RECT 54.530 187.115 56.070 187.485 ;
        RECT 52.880 185.950 53.140 186.270 ;
        RECT 53.340 185.950 53.600 186.270 ;
        RECT 53.800 185.950 54.060 186.270 ;
        RECT 51.500 184.930 51.760 185.250 ;
        RECT 51.040 175.750 51.300 176.070 ;
        RECT 50.580 174.730 50.840 175.050 ;
        RECT 48.740 174.390 49.000 174.710 ;
        RECT 48.280 173.030 48.540 173.350 ;
        RECT 48.800 173.010 48.940 174.390 ;
        RECT 49.200 174.050 49.460 174.370 ;
        RECT 48.740 172.690 49.000 173.010 ;
        RECT 45.120 170.290 45.260 171.330 ;
        RECT 45.060 169.970 45.320 170.290 ;
        RECT 46.040 169.950 46.180 171.330 ;
        RECT 47.420 171.250 48.020 171.390 ;
        RECT 47.420 169.950 47.560 171.250 ;
        RECT 44.140 169.630 44.400 169.950 ;
        RECT 45.980 169.630 46.240 169.950 ;
        RECT 47.360 169.630 47.620 169.950 ;
        RECT 47.820 169.630 48.080 169.950 ;
        RECT 44.200 169.270 44.340 169.630 ;
        RECT 44.140 168.950 44.400 169.270 ;
        RECT 42.760 164.420 43.020 164.510 ;
        RECT 42.760 164.280 43.880 164.420 ;
        RECT 42.760 164.190 43.020 164.280 ;
        RECT 43.220 158.750 43.480 159.070 ;
        RECT 43.280 157.030 43.420 158.750 ;
        RECT 43.220 156.710 43.480 157.030 ;
        RECT 43.740 156.010 43.880 164.280 ;
        RECT 43.680 155.690 43.940 156.010 ;
        RECT 40.460 153.310 40.720 153.630 ;
        RECT 42.300 153.310 42.560 153.630 ;
        RECT 41.840 152.290 42.100 152.610 ;
        RECT 41.900 150.570 42.040 152.290 ;
        RECT 42.360 151.590 42.500 153.310 ;
        RECT 42.300 151.270 42.560 151.590 ;
        RECT 44.200 150.570 44.340 168.950 ;
        RECT 45.275 168.075 46.815 168.445 ;
        RECT 46.900 165.890 47.160 166.210 ;
        RECT 46.960 164.510 47.100 165.890 ;
        RECT 46.900 164.190 47.160 164.510 ;
        RECT 47.420 164.170 47.560 169.630 ;
        RECT 47.880 165.190 48.020 169.630 ;
        RECT 48.800 166.210 48.940 172.690 ;
        RECT 49.260 170.290 49.400 174.050 ;
        RECT 51.560 172.330 51.700 184.930 ;
        RECT 53.860 181.510 54.000 185.950 ;
        RECT 54.530 181.675 56.070 182.045 ;
        RECT 52.420 181.190 52.680 181.510 ;
        RECT 53.800 181.190 54.060 181.510 ;
        RECT 52.480 177.770 52.620 181.190 ;
        RECT 53.340 180.850 53.600 181.170 ;
        RECT 53.400 178.790 53.540 180.850 ;
        RECT 54.260 180.510 54.520 180.830 ;
        RECT 54.320 178.790 54.460 180.510 ;
        RECT 53.340 178.470 53.600 178.790 ;
        RECT 54.260 178.470 54.520 178.790 ;
        RECT 51.960 177.450 52.220 177.770 ;
        RECT 52.420 177.450 52.680 177.770 ;
        RECT 52.020 173.010 52.160 177.450 ;
        RECT 52.880 176.770 53.140 177.090 ;
        RECT 52.940 175.390 53.080 176.770 ;
        RECT 54.530 176.235 56.070 176.605 ;
        RECT 56.620 176.070 56.760 188.250 ;
        RECT 57.080 177.430 57.220 188.670 ;
        RECT 57.540 186.270 57.680 190.370 ;
        RECT 58.460 188.390 58.600 191.050 ;
        RECT 58.860 190.710 59.120 191.030 ;
        RECT 59.320 190.710 59.580 191.030 ;
        RECT 58.920 189.670 59.060 190.710 ;
        RECT 58.860 189.350 59.120 189.670 ;
        RECT 58.460 188.250 59.060 188.390 ;
        RECT 58.400 187.650 58.660 187.970 ;
        RECT 58.460 186.950 58.600 187.650 ;
        RECT 58.400 186.630 58.660 186.950 ;
        RECT 58.920 186.610 59.060 188.250 ;
        RECT 58.860 186.290 59.120 186.610 ;
        RECT 57.480 185.950 57.740 186.270 ;
        RECT 57.480 185.270 57.740 185.590 ;
        RECT 57.020 177.110 57.280 177.430 ;
        RECT 56.560 175.750 56.820 176.070 ;
        RECT 52.880 175.070 53.140 175.390 ;
        RECT 53.340 175.070 53.600 175.390 ;
        RECT 52.940 173.350 53.080 175.070 ;
        RECT 52.880 173.030 53.140 173.350 ;
        RECT 51.960 172.690 52.220 173.010 ;
        RECT 51.500 172.010 51.760 172.330 ;
        RECT 52.940 171.650 53.080 173.030 ;
        RECT 52.420 171.330 52.680 171.650 ;
        RECT 52.880 171.330 53.140 171.650 ;
        RECT 49.200 169.970 49.460 170.290 ;
        RECT 50.580 169.970 50.840 170.290 ;
        RECT 48.740 165.890 49.000 166.210 ;
        RECT 47.820 164.870 48.080 165.190 ;
        RECT 47.820 164.190 48.080 164.510 ;
        RECT 47.360 163.850 47.620 164.170 ;
        RECT 45.275 162.635 46.815 163.005 ;
        RECT 47.420 158.390 47.560 163.850 ;
        RECT 47.880 162.470 48.020 164.190 ;
        RECT 47.820 162.150 48.080 162.470 ;
        RECT 47.360 158.070 47.620 158.390 ;
        RECT 45.275 157.195 46.815 157.565 ;
        RECT 44.600 155.690 44.860 156.010 ;
        RECT 45.520 155.690 45.780 156.010 ;
        RECT 41.840 150.250 42.100 150.570 ;
        RECT 44.140 150.250 44.400 150.570 ;
        RECT 38.160 149.570 38.420 149.890 ;
        RECT 36.020 149.035 37.560 149.405 ;
        RECT 26.765 146.315 28.305 146.685 ;
        RECT 38.220 145.470 38.360 149.570 ;
        RECT 38.160 145.150 38.420 145.470 ;
        RECT 36.020 143.595 37.560 143.965 ;
        RECT 44.660 142.750 44.800 155.690 ;
        RECT 45.580 154.310 45.720 155.690 ;
        RECT 45.520 153.990 45.780 154.310 ;
        RECT 46.900 153.650 47.160 153.970 ;
        RECT 45.275 151.755 46.815 152.125 ;
        RECT 46.960 151.590 47.100 153.650 ;
        RECT 47.420 153.630 47.560 158.070 ;
        RECT 48.280 155.010 48.540 155.330 ;
        RECT 48.340 154.310 48.480 155.010 ;
        RECT 48.280 153.990 48.540 154.310 ;
        RECT 48.800 153.630 48.940 165.890 ;
        RECT 50.640 164.850 50.780 169.970 ;
        RECT 51.960 168.610 52.220 168.930 ;
        RECT 52.020 167.230 52.160 168.610 ;
        RECT 51.960 166.910 52.220 167.230 ;
        RECT 50.580 164.530 50.840 164.850 ;
        RECT 50.640 161.450 50.780 164.530 ;
        RECT 50.580 161.130 50.840 161.450 ;
        RECT 50.120 160.790 50.380 161.110 ;
        RECT 50.180 158.050 50.320 160.790 ;
        RECT 52.020 160.770 52.160 166.910 ;
        RECT 51.960 160.450 52.220 160.770 ;
        RECT 52.480 159.070 52.620 171.330 ;
        RECT 52.940 162.130 53.080 171.330 ;
        RECT 53.400 170.630 53.540 175.070 ;
        RECT 57.020 172.010 57.280 172.330 ;
        RECT 54.530 170.795 56.070 171.165 ;
        RECT 53.340 170.310 53.600 170.630 ;
        RECT 57.080 167.230 57.220 172.010 ;
        RECT 57.540 170.630 57.680 185.270 ;
        RECT 59.380 185.250 59.520 190.710 ;
        RECT 59.320 184.930 59.580 185.250 ;
        RECT 58.400 183.570 58.660 183.890 ;
        RECT 58.460 181.510 58.600 183.570 ;
        RECT 58.860 183.230 59.120 183.550 ;
        RECT 58.920 181.510 59.060 183.230 ;
        RECT 58.400 181.190 58.660 181.510 ;
        RECT 58.860 181.190 59.120 181.510 ;
        RECT 58.920 180.830 59.060 181.190 ;
        RECT 57.940 180.510 58.200 180.830 ;
        RECT 58.860 180.510 59.120 180.830 ;
        RECT 58.000 178.790 58.140 180.510 ;
        RECT 58.920 178.790 59.060 180.510 ;
        RECT 57.940 178.470 58.200 178.790 ;
        RECT 58.400 178.470 58.660 178.790 ;
        RECT 58.860 178.470 59.120 178.790 ;
        RECT 58.460 178.110 58.600 178.470 ;
        RECT 58.400 177.790 58.660 178.110 ;
        RECT 58.460 175.390 58.600 177.790 ;
        RECT 58.400 175.070 58.660 175.390 ;
        RECT 58.460 172.330 58.600 175.070 ;
        RECT 58.860 172.350 59.120 172.670 ;
        RECT 58.400 172.010 58.660 172.330 ;
        RECT 58.920 171.990 59.060 172.350 ;
        RECT 58.860 171.670 59.120 171.990 ;
        RECT 57.480 170.310 57.740 170.630 ;
        RECT 57.020 166.910 57.280 167.230 ;
        RECT 53.800 166.570 54.060 166.890 ;
        RECT 56.560 166.570 56.820 166.890 ;
        RECT 58.920 166.630 59.060 171.670 ;
        RECT 59.840 169.950 59.980 191.050 ;
        RECT 60.240 187.990 60.500 188.310 ;
        RECT 60.300 186.950 60.440 187.990 ;
        RECT 60.240 186.630 60.500 186.950 ;
        RECT 60.240 182.550 60.500 182.870 ;
        RECT 60.300 174.370 60.440 182.550 ;
        RECT 60.760 177.430 60.900 193.770 ;
        RECT 61.220 191.030 61.360 201.250 ;
        RECT 61.680 200.550 61.820 202.270 ;
        RECT 63.000 201.930 63.260 202.250 ;
        RECT 66.220 201.930 66.480 202.250 ;
        RECT 66.680 201.930 66.940 202.250 ;
        RECT 61.620 200.230 61.880 200.550 ;
        RECT 62.080 196.830 62.340 197.150 ;
        RECT 62.140 195.110 62.280 196.830 ;
        RECT 62.080 194.790 62.340 195.110 ;
        RECT 61.160 190.710 61.420 191.030 ;
        RECT 61.620 190.370 61.880 190.690 ;
        RECT 62.540 190.370 62.800 190.690 ;
        RECT 61.680 188.650 61.820 190.370 ;
        RECT 62.080 189.350 62.340 189.670 ;
        RECT 61.620 188.330 61.880 188.650 ;
        RECT 62.140 183.210 62.280 189.350 ;
        RECT 62.600 188.650 62.740 190.370 ;
        RECT 63.060 188.990 63.200 201.930 ;
        RECT 63.785 200.715 65.325 201.085 ;
        RECT 66.280 200.550 66.420 201.930 ;
        RECT 66.220 200.230 66.480 200.550 ;
        RECT 66.740 199.530 66.880 201.930 ;
        RECT 66.680 199.210 66.940 199.530 ;
        RECT 63.785 195.275 65.325 195.645 ;
        RECT 66.740 194.430 66.880 199.210 ;
        RECT 67.600 195.810 67.860 196.130 ;
        RECT 66.680 194.110 66.940 194.430 ;
        RECT 67.660 194.090 67.800 195.810 ;
        RECT 67.600 193.770 67.860 194.090 ;
        RECT 67.660 191.030 67.800 193.770 ;
        RECT 68.120 193.410 68.260 204.310 ;
        RECT 69.440 203.970 69.700 204.290 ;
        RECT 69.500 200.210 69.640 203.970 ;
        RECT 69.960 200.550 70.100 205.670 ;
        RECT 71.340 204.970 71.480 208.180 ;
        RECT 77.780 204.970 77.920 208.180 ;
        RECT 82.295 206.155 83.835 206.525 ;
        RECT 84.220 204.970 84.360 208.180 ;
        RECT 71.280 204.650 71.540 204.970 ;
        RECT 77.720 204.650 77.980 204.970 ;
        RECT 84.160 204.650 84.420 204.970 ;
        RECT 72.200 203.970 72.460 204.290 ;
        RECT 79.560 203.970 79.820 204.290 ;
        RECT 85.540 203.970 85.800 204.290 ;
        RECT 72.260 202.250 72.400 203.970 ;
        RECT 73.040 203.435 74.580 203.805 ;
        RECT 79.620 202.930 79.760 203.970 ;
        RECT 85.600 203.270 85.740 203.970 ;
        RECT 85.540 202.950 85.800 203.270 ;
        RECT 79.560 202.610 79.820 202.930 ;
        RECT 77.720 202.270 77.980 202.590 ;
        RECT 72.200 201.930 72.460 202.250 ;
        RECT 70.360 201.250 70.620 201.570 ;
        RECT 69.900 200.230 70.160 200.550 ;
        RECT 69.440 199.890 69.700 200.210 ;
        RECT 68.980 194.790 69.240 195.110 ;
        RECT 68.060 193.090 68.320 193.410 ;
        RECT 67.600 190.710 67.860 191.030 ;
        RECT 63.785 189.835 65.325 190.205 ;
        RECT 63.000 188.670 63.260 188.990 ;
        RECT 62.540 188.330 62.800 188.650 ;
        RECT 63.920 187.990 64.180 188.310 ;
        RECT 63.980 186.950 64.120 187.990 ;
        RECT 63.920 186.630 64.180 186.950 ;
        RECT 66.220 185.950 66.480 186.270 ;
        RECT 63.000 185.270 63.260 185.590 ;
        RECT 65.760 185.270 66.020 185.590 ;
        RECT 62.540 184.930 62.800 185.250 ;
        RECT 62.080 182.890 62.340 183.210 ;
        RECT 62.600 182.270 62.740 184.930 ;
        RECT 62.140 182.130 62.740 182.270 ;
        RECT 62.140 180.150 62.280 182.130 ;
        RECT 63.060 181.590 63.200 185.270 ;
        RECT 63.785 184.395 65.325 184.765 ;
        RECT 62.600 181.450 63.200 181.590 ;
        RECT 62.600 180.830 62.740 181.450 ;
        RECT 62.540 180.510 62.800 180.830 ;
        RECT 62.080 179.830 62.340 180.150 ;
        RECT 60.700 177.110 60.960 177.430 ;
        RECT 61.160 176.770 61.420 177.090 ;
        RECT 60.240 174.050 60.500 174.370 ;
        RECT 59.780 169.630 60.040 169.950 ;
        RECT 59.840 166.890 59.980 169.630 ;
        RECT 53.860 165.190 54.000 166.570 ;
        RECT 54.530 165.355 56.070 165.725 ;
        RECT 53.800 164.870 54.060 165.190 ;
        RECT 53.860 164.510 54.000 164.870 ;
        RECT 56.620 164.850 56.760 166.570 ;
        RECT 58.920 166.550 59.520 166.630 ;
        RECT 59.780 166.570 60.040 166.890 ;
        RECT 57.020 166.230 57.280 166.550 ;
        RECT 58.920 166.490 59.580 166.550 ;
        RECT 59.320 166.230 59.580 166.490 ;
        RECT 57.080 165.190 57.220 166.230 ;
        RECT 57.480 165.890 57.740 166.210 ;
        RECT 57.540 165.190 57.680 165.890 ;
        RECT 59.840 165.190 59.980 166.570 ;
        RECT 57.020 164.870 57.280 165.190 ;
        RECT 57.480 164.870 57.740 165.190 ;
        RECT 59.780 164.870 60.040 165.190 ;
        RECT 56.560 164.530 56.820 164.850 ;
        RECT 53.800 164.190 54.060 164.510 ;
        RECT 52.880 161.810 53.140 162.130 ;
        RECT 53.340 161.810 53.600 162.130 ;
        RECT 52.870 160.935 53.150 161.305 ;
        RECT 52.420 158.750 52.680 159.070 ;
        RECT 52.480 158.470 52.620 158.750 ;
        RECT 51.560 158.330 52.620 158.470 ;
        RECT 50.120 157.730 50.380 158.050 ;
        RECT 50.180 156.350 50.320 157.730 ;
        RECT 50.120 156.030 50.380 156.350 ;
        RECT 47.360 153.310 47.620 153.630 ;
        RECT 48.740 153.310 49.000 153.630 ;
        RECT 51.560 152.610 51.700 158.330 ;
        RECT 52.940 157.850 53.080 160.935 ;
        RECT 52.480 157.710 53.080 157.850 ;
        RECT 51.960 155.010 52.220 155.330 ;
        RECT 52.020 153.290 52.160 155.010 ;
        RECT 52.480 153.630 52.620 157.710 ;
        RECT 52.880 155.010 53.140 155.330 ;
        RECT 52.940 153.710 53.080 155.010 ;
        RECT 53.400 154.310 53.540 161.810 ;
        RECT 53.860 157.850 54.000 164.190 ;
        RECT 58.400 163.170 58.660 163.490 ;
        RECT 58.460 161.450 58.600 163.170 ;
        RECT 54.250 160.935 54.530 161.305 ;
        RECT 58.400 161.130 58.660 161.450 ;
        RECT 54.320 160.770 54.460 160.935 ;
        RECT 56.560 160.790 56.820 161.110 ;
        RECT 54.260 160.450 54.520 160.770 ;
        RECT 54.530 159.915 56.070 160.285 ;
        RECT 56.620 159.070 56.760 160.790 ;
        RECT 60.300 159.410 60.440 174.050 ;
        RECT 61.220 172.330 61.360 176.770 ;
        RECT 61.160 172.010 61.420 172.330 ;
        RECT 60.700 171.330 60.960 171.650 ;
        RECT 60.760 170.630 60.900 171.330 ;
        RECT 60.700 170.310 60.960 170.630 ;
        RECT 60.700 169.290 60.960 169.610 ;
        RECT 60.760 163.830 60.900 169.290 ;
        RECT 61.220 167.910 61.360 172.010 ;
        RECT 62.140 169.610 62.280 179.830 ;
        RECT 62.600 177.090 62.740 180.510 ;
        RECT 65.820 179.810 65.960 185.270 ;
        RECT 66.280 184.230 66.420 185.950 ;
        RECT 67.140 184.930 67.400 185.250 ;
        RECT 66.220 183.910 66.480 184.230 ;
        RECT 66.220 182.890 66.480 183.210 ;
        RECT 66.280 181.170 66.420 182.890 ;
        RECT 66.680 182.210 66.940 182.530 ;
        RECT 66.740 181.170 66.880 182.210 ;
        RECT 66.220 180.850 66.480 181.170 ;
        RECT 66.680 180.850 66.940 181.170 ;
        RECT 67.200 180.830 67.340 184.930 ;
        RECT 67.140 180.510 67.400 180.830 ;
        RECT 66.220 179.830 66.480 180.150 ;
        RECT 65.760 179.490 66.020 179.810 ;
        RECT 63.785 178.955 65.325 179.325 ;
        RECT 66.280 177.770 66.420 179.830 ;
        RECT 66.220 177.450 66.480 177.770 ;
        RECT 62.540 176.770 62.800 177.090 ;
        RECT 62.080 169.290 62.340 169.610 ;
        RECT 62.600 169.270 62.740 176.770 ;
        RECT 63.785 173.515 65.325 173.885 ;
        RECT 63.920 171.670 64.180 171.990 ;
        RECT 63.980 170.630 64.120 171.670 ;
        RECT 63.920 170.310 64.180 170.630 ;
        RECT 67.600 169.630 67.860 169.950 ;
        RECT 62.540 168.950 62.800 169.270 ;
        RECT 63.785 168.075 65.325 168.445 ;
        RECT 61.160 167.590 61.420 167.910 ;
        RECT 67.660 167.230 67.800 169.630 ;
        RECT 68.120 167.230 68.260 193.090 ;
        RECT 69.040 175.050 69.180 194.790 ;
        RECT 69.500 177.770 69.640 199.890 ;
        RECT 70.420 199.530 70.560 201.250 ;
        RECT 70.820 200.230 71.080 200.550 ;
        RECT 70.360 199.210 70.620 199.530 ;
        RECT 70.880 195.110 71.020 200.230 ;
        RECT 71.740 196.490 72.000 196.810 ;
        RECT 70.820 194.790 71.080 195.110 ;
        RECT 71.800 193.410 71.940 196.490 ;
        RECT 71.740 193.090 72.000 193.410 ;
        RECT 71.800 188.650 71.940 193.090 ;
        RECT 71.740 188.330 72.000 188.650 ;
        RECT 71.280 187.650 71.540 187.970 ;
        RECT 71.340 186.270 71.480 187.650 ;
        RECT 71.280 185.950 71.540 186.270 ;
        RECT 69.900 181.190 70.160 181.510 ;
        RECT 69.960 178.450 70.100 181.190 ;
        RECT 71.280 180.850 71.540 181.170 ;
        RECT 70.820 180.170 71.080 180.490 ;
        RECT 69.900 178.130 70.160 178.450 ;
        RECT 69.960 177.770 70.100 178.130 ;
        RECT 69.440 177.450 69.700 177.770 ;
        RECT 69.900 177.450 70.160 177.770 ;
        RECT 69.960 177.090 70.100 177.450 ;
        RECT 69.900 176.770 70.160 177.090 ;
        RECT 70.360 176.770 70.620 177.090 ;
        RECT 70.420 175.390 70.560 176.770 ;
        RECT 70.360 175.070 70.620 175.390 ;
        RECT 68.980 174.730 69.240 175.050 ;
        RECT 70.880 174.960 71.020 180.170 ;
        RECT 71.340 177.770 71.480 180.850 ;
        RECT 71.800 178.790 71.940 188.330 ;
        RECT 71.740 178.470 72.000 178.790 ;
        RECT 71.280 177.450 71.540 177.770 ;
        RECT 71.800 177.625 71.940 178.470 ;
        RECT 71.730 177.255 72.010 177.625 ;
        RECT 71.280 174.960 71.540 175.050 ;
        RECT 70.880 174.820 71.540 174.960 ;
        RECT 71.280 174.730 71.540 174.820 ;
        RECT 67.600 166.910 67.860 167.230 ;
        RECT 68.060 166.910 68.320 167.230 ;
        RECT 66.680 166.230 66.940 166.550 ;
        RECT 66.740 164.510 66.880 166.230 ;
        RECT 68.060 165.890 68.320 166.210 ;
        RECT 68.120 164.510 68.260 165.890 ;
        RECT 63.000 164.190 63.260 164.510 ;
        RECT 66.680 164.190 66.940 164.510 ;
        RECT 68.060 164.190 68.320 164.510 ;
        RECT 68.520 164.190 68.780 164.510 ;
        RECT 60.700 163.510 60.960 163.830 ;
        RECT 63.060 162.470 63.200 164.190 ;
        RECT 63.785 162.635 65.325 163.005 ;
        RECT 68.580 162.470 68.720 164.190 ;
        RECT 63.000 162.150 63.260 162.470 ;
        RECT 68.520 162.150 68.780 162.470 ;
        RECT 69.040 161.110 69.180 174.730 ;
        RECT 69.900 172.690 70.160 173.010 ;
        RECT 69.440 172.010 69.700 172.330 ;
        RECT 69.500 164.510 69.640 172.010 ;
        RECT 69.440 164.190 69.700 164.510 ;
        RECT 68.060 160.790 68.320 161.110 ;
        RECT 68.980 160.790 69.240 161.110 ;
        RECT 60.240 159.090 60.500 159.410 ;
        RECT 56.560 158.750 56.820 159.070 ;
        RECT 55.640 158.410 55.900 158.730 ;
        RECT 53.860 157.710 54.460 157.850 ;
        RECT 54.320 155.670 54.460 157.710 ;
        RECT 55.700 156.350 55.840 158.410 ;
        RECT 56.560 157.730 56.820 158.050 ;
        RECT 56.620 156.690 56.760 157.730 ;
        RECT 63.785 157.195 65.325 157.565 ;
        RECT 56.560 156.370 56.820 156.690 ;
        RECT 55.640 156.030 55.900 156.350 ;
        RECT 54.260 155.350 54.520 155.670 ;
        RECT 53.800 155.010 54.060 155.330 ;
        RECT 53.860 154.310 54.000 155.010 ;
        RECT 54.530 154.475 56.070 154.845 ;
        RECT 53.340 153.990 53.600 154.310 ;
        RECT 53.800 153.990 54.060 154.310 ;
        RECT 52.940 153.630 53.540 153.710 ;
        RECT 54.720 153.650 54.980 153.970 ;
        RECT 56.620 153.710 56.760 156.370 ;
        RECT 57.020 155.690 57.280 156.010 ;
        RECT 67.600 155.690 67.860 156.010 ;
        RECT 57.080 154.310 57.220 155.690 ;
        RECT 65.300 155.010 65.560 155.330 ;
        RECT 65.760 155.010 66.020 155.330 ;
        RECT 57.020 153.990 57.280 154.310 ;
        RECT 52.420 153.310 52.680 153.630 ;
        RECT 52.940 153.570 53.600 153.630 ;
        RECT 53.340 153.310 53.600 153.570 ;
        RECT 51.960 152.970 52.220 153.290 ;
        RECT 52.880 152.630 53.140 152.950 ;
        RECT 51.500 152.290 51.760 152.610 ;
        RECT 52.940 151.590 53.080 152.630 ;
        RECT 46.900 151.270 47.160 151.590 ;
        RECT 52.880 151.270 53.140 151.590 ;
        RECT 48.740 149.910 49.000 150.230 ;
        RECT 48.800 147.510 48.940 149.910 ;
        RECT 53.400 149.890 53.540 153.310 ;
        RECT 54.780 150.230 54.920 153.650 ;
        RECT 55.180 153.310 55.440 153.630 ;
        RECT 56.620 153.570 57.220 153.710 ;
        RECT 55.240 150.570 55.380 153.310 ;
        RECT 56.100 152.970 56.360 153.290 ;
        RECT 56.160 150.910 56.300 152.970 ;
        RECT 56.100 150.590 56.360 150.910 ;
        RECT 55.180 150.250 55.440 150.570 ;
        RECT 56.560 150.250 56.820 150.570 ;
        RECT 53.800 149.910 54.060 150.230 ;
        RECT 54.720 149.910 54.980 150.230 ;
        RECT 53.340 149.570 53.600 149.890 ;
        RECT 53.400 148.870 53.540 149.570 ;
        RECT 53.340 148.550 53.600 148.870 ;
        RECT 53.860 147.590 54.000 149.910 ;
        RECT 54.530 149.035 56.070 149.405 ;
        RECT 55.180 148.210 55.440 148.530 ;
        RECT 54.260 147.590 54.520 147.850 ;
        RECT 53.860 147.530 54.520 147.590 ;
        RECT 48.740 147.190 49.000 147.510 ;
        RECT 53.860 147.450 54.460 147.530 ;
        RECT 45.275 146.315 46.815 146.685 ;
        RECT 48.800 145.130 48.940 147.190 ;
        RECT 53.340 146.850 53.600 147.170 ;
        RECT 53.400 145.130 53.540 146.850 ;
        RECT 53.860 146.150 54.000 147.450 ;
        RECT 53.800 145.830 54.060 146.150 ;
        RECT 55.240 145.470 55.380 148.210 ;
        RECT 55.180 145.150 55.440 145.470 ;
        RECT 56.620 145.130 56.760 150.250 ;
        RECT 57.080 147.170 57.220 153.570 ;
        RECT 65.360 153.030 65.500 155.010 ;
        RECT 65.820 153.630 65.960 155.010 ;
        RECT 65.760 153.310 66.020 153.630 ;
        RECT 67.660 153.145 67.800 155.690 ;
        RECT 65.360 152.890 66.880 153.030 ;
        RECT 63.000 152.290 63.260 152.610 ;
        RECT 59.320 150.930 59.580 151.250 ;
        RECT 60.240 150.930 60.500 151.250 ;
        RECT 59.380 150.230 59.520 150.930 ;
        RECT 59.320 149.910 59.580 150.230 ;
        RECT 59.320 147.530 59.580 147.850 ;
        RECT 57.020 146.850 57.280 147.170 ;
        RECT 59.380 146.150 59.520 147.530 ;
        RECT 59.320 145.830 59.580 146.150 ;
        RECT 60.300 145.130 60.440 150.930 ;
        RECT 63.060 150.570 63.200 152.290 ;
        RECT 63.785 151.755 65.325 152.125 ;
        RECT 61.620 150.250 61.880 150.570 ;
        RECT 63.000 150.250 63.260 150.570 ;
        RECT 61.160 149.570 61.420 149.890 ;
        RECT 61.220 148.870 61.360 149.570 ;
        RECT 61.680 148.870 61.820 150.250 ;
        RECT 62.540 149.570 62.800 149.890 ;
        RECT 61.160 148.550 61.420 148.870 ;
        RECT 61.620 148.550 61.880 148.870 ;
        RECT 62.600 148.190 62.740 149.570 ;
        RECT 66.740 148.870 66.880 152.890 ;
        RECT 67.590 152.775 67.870 153.145 ;
        RECT 67.660 150.570 67.800 152.775 ;
        RECT 68.120 150.570 68.260 160.790 ;
        RECT 69.500 159.750 69.640 164.190 ;
        RECT 69.960 160.770 70.100 172.690 ;
        RECT 71.800 170.290 71.940 177.255 ;
        RECT 71.740 169.970 72.000 170.290 ;
        RECT 72.260 169.610 72.400 201.930 ;
        RECT 75.880 200.230 76.140 200.550 ;
        RECT 75.940 199.530 76.080 200.230 ;
        RECT 74.960 199.210 75.220 199.530 ;
        RECT 75.880 199.210 76.140 199.530 ;
        RECT 76.340 199.210 76.600 199.530 ;
        RECT 77.260 199.385 77.520 199.530 ;
        RECT 72.660 198.870 72.920 199.190 ;
        RECT 72.720 194.090 72.860 198.870 ;
        RECT 73.040 197.995 74.580 198.365 ;
        RECT 75.020 197.830 75.160 199.210 ;
        RECT 74.960 197.510 75.220 197.830 ;
        RECT 75.880 197.170 76.140 197.490 ;
        RECT 74.500 196.830 74.760 197.150 ;
        RECT 74.960 196.830 75.220 197.150 ;
        RECT 74.560 195.110 74.700 196.830 ;
        RECT 74.500 194.790 74.760 195.110 ;
        RECT 75.020 194.430 75.160 196.830 ;
        RECT 74.960 194.110 75.220 194.430 ;
        RECT 72.660 193.770 72.920 194.090 ;
        RECT 75.420 193.090 75.680 193.410 ;
        RECT 73.040 192.555 74.580 192.925 ;
        RECT 75.480 192.390 75.620 193.090 ;
        RECT 74.960 192.070 75.220 192.390 ;
        RECT 75.420 192.070 75.680 192.390 ;
        RECT 72.660 191.050 72.920 191.370 ;
        RECT 72.720 185.930 72.860 191.050 ;
        RECT 73.040 187.115 74.580 187.485 ;
        RECT 75.020 186.950 75.160 192.070 ;
        RECT 74.960 186.630 75.220 186.950 ;
        RECT 75.940 186.270 76.080 197.170 ;
        RECT 75.880 185.950 76.140 186.270 ;
        RECT 72.660 185.610 72.920 185.930 ;
        RECT 72.720 173.010 72.860 185.610 ;
        RECT 75.880 182.550 76.140 182.870 ;
        RECT 73.040 181.675 74.580 182.045 ;
        RECT 75.940 178.110 76.080 182.550 ;
        RECT 76.400 181.170 76.540 199.210 ;
        RECT 77.250 199.015 77.530 199.385 ;
        RECT 76.800 198.530 77.060 198.850 ;
        RECT 76.860 197.830 77.000 198.530 ;
        RECT 77.780 197.830 77.920 202.270 ;
        RECT 86.460 201.250 86.720 201.570 ;
        RECT 82.295 200.715 83.835 201.085 ;
        RECT 85.080 200.230 85.340 200.550 ;
        RECT 80.020 199.890 80.280 200.210 ;
        RECT 78.640 199.210 78.900 199.530 ;
        RECT 78.700 197.830 78.840 199.210 ;
        RECT 79.560 198.530 79.820 198.850 ;
        RECT 76.800 197.510 77.060 197.830 ;
        RECT 77.720 197.510 77.980 197.830 ;
        RECT 78.640 197.510 78.900 197.830 ;
        RECT 79.620 197.150 79.760 198.530 ;
        RECT 80.080 197.150 80.220 199.890 ;
        RECT 80.480 198.870 80.740 199.190 ;
        RECT 77.260 196.830 77.520 197.150 ;
        RECT 79.560 196.830 79.820 197.150 ;
        RECT 80.020 196.830 80.280 197.150 ;
        RECT 77.320 194.430 77.460 196.830 ;
        RECT 78.180 195.810 78.440 196.130 ;
        RECT 77.260 194.110 77.520 194.430 ;
        RECT 76.800 193.430 77.060 193.750 ;
        RECT 76.860 191.370 77.000 193.430 ;
        RECT 76.800 191.050 77.060 191.370 ;
        RECT 77.320 186.270 77.460 194.110 ;
        RECT 78.240 192.390 78.380 195.810 ;
        RECT 78.640 194.450 78.900 194.770 ;
        RECT 80.020 194.450 80.280 194.770 ;
        RECT 78.700 193.750 78.840 194.450 ;
        RECT 80.080 193.750 80.220 194.450 ;
        RECT 78.640 193.430 78.900 193.750 ;
        RECT 80.020 193.430 80.280 193.750 ;
        RECT 78.180 192.070 78.440 192.390 ;
        RECT 78.700 189.670 78.840 193.430 ;
        RECT 78.640 189.350 78.900 189.670 ;
        RECT 80.020 189.350 80.280 189.670 ;
        RECT 80.080 188.390 80.220 189.350 ;
        RECT 79.620 188.250 80.220 188.390 ;
        RECT 77.720 187.650 77.980 187.970 ;
        RECT 77.780 186.270 77.920 187.650 ;
        RECT 77.260 185.950 77.520 186.270 ;
        RECT 77.720 185.950 77.980 186.270 ;
        RECT 78.640 185.950 78.900 186.270 ;
        RECT 79.100 185.950 79.360 186.270 ;
        RECT 77.320 183.550 77.460 185.950 ;
        RECT 77.720 184.930 77.980 185.250 ;
        RECT 77.260 183.230 77.520 183.550 ;
        RECT 76.340 180.850 76.600 181.170 ;
        RECT 75.880 177.790 76.140 178.110 ;
        RECT 73.040 176.235 74.580 176.605 ;
        RECT 73.120 175.750 73.380 176.070 ;
        RECT 74.040 175.750 74.300 176.070 ;
        RECT 73.180 175.470 73.320 175.750 ;
        RECT 74.100 175.470 74.240 175.750 ;
        RECT 76.400 175.730 76.540 180.850 ;
        RECT 77.320 180.230 77.460 183.230 ;
        RECT 77.780 180.830 77.920 184.930 ;
        RECT 78.700 184.230 78.840 185.950 ;
        RECT 78.640 183.910 78.900 184.230 ;
        RECT 77.720 180.510 77.980 180.830 ;
        RECT 77.320 180.090 77.920 180.230 ;
        RECT 77.780 179.810 77.920 180.090 ;
        RECT 77.720 179.490 77.980 179.810 ;
        RECT 77.780 177.770 77.920 179.490 ;
        RECT 78.640 178.190 78.900 178.450 ;
        RECT 79.160 178.190 79.300 185.950 ;
        RECT 79.620 183.890 79.760 188.250 ;
        RECT 80.020 187.650 80.280 187.970 ;
        RECT 79.560 183.570 79.820 183.890 ;
        RECT 79.620 180.910 79.760 183.570 ;
        RECT 80.080 183.210 80.220 187.650 ;
        RECT 80.020 182.890 80.280 183.210 ;
        RECT 80.020 182.210 80.280 182.530 ;
        RECT 80.080 181.025 80.220 182.210 ;
        RECT 80.010 180.910 80.290 181.025 ;
        RECT 79.620 180.830 80.290 180.910 ;
        RECT 79.560 180.770 80.290 180.830 ;
        RECT 79.560 180.510 79.820 180.770 ;
        RECT 80.010 180.655 80.290 180.770 ;
        RECT 79.550 179.975 79.830 180.345 ;
        RECT 79.560 179.830 79.820 179.975 ;
        RECT 78.640 178.130 79.300 178.190 ;
        RECT 78.700 178.050 79.300 178.130 ;
        RECT 77.720 177.450 77.980 177.770 ;
        RECT 78.640 177.450 78.900 177.770 ;
        RECT 79.160 177.680 79.300 178.050 ;
        RECT 79.560 177.680 79.820 177.770 ;
        RECT 79.160 177.540 79.820 177.680 ;
        RECT 79.560 177.450 79.820 177.540 ;
        RECT 73.180 175.330 74.240 175.470 ;
        RECT 76.340 175.410 76.600 175.730 ;
        RECT 75.420 175.070 75.680 175.390 ;
        RECT 73.120 174.960 73.380 175.050 ;
        RECT 74.040 174.960 74.300 175.050 ;
        RECT 73.120 174.820 74.300 174.960 ;
        RECT 73.120 174.730 73.380 174.820 ;
        RECT 74.040 174.730 74.300 174.820 ;
        RECT 74.040 174.050 74.300 174.370 ;
        RECT 74.500 174.050 74.760 174.370 ;
        RECT 72.660 172.690 72.920 173.010 ;
        RECT 74.100 172.330 74.240 174.050 ;
        RECT 74.560 173.350 74.700 174.050 ;
        RECT 75.480 173.350 75.620 175.070 ;
        RECT 74.500 173.030 74.760 173.350 ;
        RECT 75.420 173.030 75.680 173.350 ;
        RECT 74.040 172.010 74.300 172.330 ;
        RECT 72.660 171.330 72.920 171.650 ;
        RECT 72.720 169.950 72.860 171.330 ;
        RECT 73.040 170.795 74.580 171.165 ;
        RECT 72.660 169.630 72.920 169.950 ;
        RECT 76.800 169.630 77.060 169.950 ;
        RECT 72.200 169.290 72.460 169.610 ;
        RECT 76.340 168.610 76.600 168.930 ;
        RECT 75.880 166.570 76.140 166.890 ;
        RECT 73.040 165.355 74.580 165.725 ;
        RECT 75.940 165.190 76.080 166.570 ;
        RECT 74.040 164.870 74.300 165.190 ;
        RECT 75.880 164.870 76.140 165.190 ;
        RECT 74.100 161.110 74.240 164.870 ;
        RECT 74.960 161.470 75.220 161.790 ;
        RECT 72.200 160.790 72.460 161.110 ;
        RECT 74.040 160.790 74.300 161.110 ;
        RECT 69.900 160.450 70.160 160.770 ;
        RECT 69.440 159.430 69.700 159.750 ;
        RECT 69.960 158.050 70.100 160.450 ;
        RECT 69.900 157.850 70.160 158.050 ;
        RECT 69.040 157.730 70.160 157.850 ;
        RECT 69.040 157.710 70.100 157.730 ;
        RECT 69.040 157.110 69.180 157.710 ;
        RECT 68.580 156.970 69.180 157.110 ;
        RECT 72.260 157.030 72.400 160.790 ;
        RECT 75.020 160.770 75.160 161.470 ;
        RECT 76.400 161.450 76.540 168.610 ;
        RECT 76.860 166.890 77.000 169.630 ;
        RECT 76.800 166.570 77.060 166.890 ;
        RECT 77.780 164.850 77.920 177.450 ;
        RECT 78.700 175.730 78.840 177.450 ;
        RECT 78.640 175.410 78.900 175.730 ;
        RECT 78.180 175.070 78.440 175.390 ;
        RECT 78.240 172.670 78.380 175.070 ;
        RECT 79.560 173.030 79.820 173.350 ;
        RECT 78.180 172.350 78.440 172.670 ;
        RECT 79.620 171.650 79.760 173.030 ;
        RECT 78.640 171.330 78.900 171.650 ;
        RECT 79.560 171.330 79.820 171.650 ;
        RECT 78.700 167.230 78.840 171.330 ;
        RECT 79.620 169.950 79.760 171.330 ;
        RECT 79.560 169.630 79.820 169.950 ;
        RECT 78.640 166.910 78.900 167.230 ;
        RECT 78.640 166.230 78.900 166.550 ;
        RECT 77.720 164.530 77.980 164.850 ;
        RECT 78.700 164.510 78.840 166.230 ;
        RECT 78.640 164.190 78.900 164.510 ;
        RECT 79.620 163.830 79.760 169.630 ;
        RECT 79.560 163.510 79.820 163.830 ;
        RECT 78.180 163.170 78.440 163.490 ;
        RECT 80.540 163.230 80.680 198.870 ;
        RECT 81.860 197.170 82.120 197.490 ;
        RECT 81.920 191.710 82.060 197.170 ;
        RECT 82.295 195.275 83.835 195.645 ;
        RECT 85.140 194.090 85.280 200.230 ;
        RECT 86.520 199.870 86.660 201.250 ;
        RECT 86.460 199.550 86.720 199.870 ;
        RECT 87.840 199.385 88.100 199.530 ;
        RECT 87.830 199.015 88.110 199.385 ;
        RECT 88.760 198.530 89.020 198.850 ;
        RECT 88.820 194.090 88.960 198.530 ;
        RECT 85.080 193.770 85.340 194.090 ;
        RECT 86.460 193.770 86.720 194.090 ;
        RECT 88.760 193.770 89.020 194.090 ;
        RECT 83.700 193.090 83.960 193.410 ;
        RECT 83.760 191.710 83.900 193.090 ;
        RECT 81.860 191.390 82.120 191.710 ;
        RECT 83.700 191.390 83.960 191.710 ;
        RECT 80.940 187.990 81.200 188.310 ;
        RECT 81.000 185.590 81.140 187.990 ;
        RECT 81.920 186.270 82.060 191.390 ;
        RECT 82.295 189.835 83.835 190.205 ;
        RECT 85.140 188.650 85.280 193.770 ;
        RECT 86.520 188.650 86.660 193.770 ;
        RECT 85.080 188.330 85.340 188.650 ;
        RECT 85.540 188.330 85.800 188.650 ;
        RECT 86.460 188.330 86.720 188.650 ;
        RECT 83.700 187.650 83.960 187.970 ;
        RECT 83.760 186.270 83.900 187.650 ;
        RECT 81.860 185.950 82.120 186.270 ;
        RECT 83.700 185.950 83.960 186.270 ;
        RECT 81.400 185.610 81.660 185.930 ;
        RECT 80.940 185.270 81.200 185.590 ;
        RECT 81.000 184.230 81.140 185.270 ;
        RECT 81.460 184.230 81.600 185.610 ;
        RECT 80.940 183.910 81.200 184.230 ;
        RECT 81.400 183.910 81.660 184.230 ;
        RECT 80.940 182.890 81.200 183.210 ;
        RECT 81.000 182.530 81.140 182.890 ;
        RECT 81.920 182.870 82.060 185.950 ;
        RECT 82.295 184.395 83.835 184.765 ;
        RECT 81.860 182.550 82.120 182.870 ;
        RECT 80.940 182.210 81.200 182.530 ;
        RECT 81.000 177.000 81.140 182.210 ;
        RECT 81.920 180.230 82.060 182.550 ;
        RECT 82.780 180.510 83.040 180.830 ;
        RECT 82.320 180.230 82.580 180.490 ;
        RECT 82.840 180.345 82.980 180.510 ;
        RECT 81.920 180.170 82.580 180.230 ;
        RECT 81.400 179.830 81.660 180.150 ;
        RECT 81.920 180.090 82.520 180.170 ;
        RECT 81.460 178.790 81.600 179.830 ;
        RECT 81.400 178.470 81.660 178.790 ;
        RECT 81.400 177.625 81.660 177.770 ;
        RECT 81.390 177.255 81.670 177.625 ;
        RECT 81.400 177.000 81.660 177.090 ;
        RECT 81.000 176.860 81.660 177.000 ;
        RECT 81.400 176.770 81.660 176.860 ;
        RECT 81.460 173.350 81.600 176.770 ;
        RECT 81.920 175.730 82.060 180.090 ;
        RECT 82.770 179.975 83.050 180.345 ;
        RECT 82.295 178.955 83.835 179.325 ;
        RECT 85.140 177.770 85.280 188.330 ;
        RECT 85.600 186.950 85.740 188.330 ;
        RECT 85.540 186.630 85.800 186.950 ;
        RECT 86.520 185.450 86.660 188.330 ;
        RECT 86.060 185.310 86.660 185.450 ;
        RECT 86.060 181.510 86.200 185.310 ;
        RECT 86.000 181.190 86.260 181.510 ;
        RECT 86.060 177.770 86.200 181.190 ;
        RECT 85.080 177.450 85.340 177.770 ;
        RECT 86.000 177.450 86.260 177.770 ;
        RECT 90.140 177.450 90.400 177.770 ;
        RECT 83.700 176.770 83.960 177.090 ;
        RECT 81.860 175.410 82.120 175.730 ;
        RECT 83.760 175.390 83.900 176.770 ;
        RECT 85.140 175.390 85.280 177.450 ;
        RECT 83.700 175.070 83.960 175.390 ;
        RECT 85.080 175.070 85.340 175.390 ;
        RECT 82.295 173.515 83.835 173.885 ;
        RECT 81.400 173.030 81.660 173.350 ;
        RECT 85.140 172.330 85.280 175.070 ;
        RECT 85.080 172.010 85.340 172.330 ;
        RECT 81.400 171.330 81.660 171.650 ;
        RECT 83.700 171.330 83.960 171.650 ;
        RECT 80.940 167.250 81.200 167.570 ;
        RECT 81.000 164.510 81.140 167.250 ;
        RECT 81.460 166.890 81.600 171.330 ;
        RECT 83.760 169.950 83.900 171.330 ;
        RECT 83.700 169.630 83.960 169.950 ;
        RECT 81.860 169.290 82.120 169.610 ;
        RECT 81.400 166.570 81.660 166.890 ;
        RECT 81.920 164.850 82.060 169.290 ;
        RECT 82.295 168.075 83.835 168.445 ;
        RECT 85.140 165.190 85.280 172.010 ;
        RECT 85.080 164.870 85.340 165.190 ;
        RECT 81.860 164.530 82.120 164.850 ;
        RECT 80.940 164.190 81.200 164.510 ;
        RECT 78.240 161.450 78.380 163.170 ;
        RECT 80.080 163.090 80.680 163.230 ;
        RECT 80.080 161.450 80.220 163.090 ;
        RECT 80.480 161.810 80.740 162.130 ;
        RECT 76.340 161.130 76.600 161.450 ;
        RECT 78.180 161.130 78.440 161.450 ;
        RECT 80.020 161.130 80.280 161.450 ;
        RECT 74.960 160.450 75.220 160.770 ;
        RECT 73.040 159.915 74.580 160.285 ;
        RECT 75.420 159.430 75.680 159.750 ;
        RECT 68.580 156.350 68.720 156.970 ;
        RECT 72.200 156.710 72.460 157.030 ;
        RECT 68.520 156.030 68.780 156.350 ;
        RECT 68.980 155.690 69.240 156.010 ;
        RECT 69.440 155.690 69.700 156.010 ;
        RECT 69.040 152.950 69.180 155.690 ;
        RECT 69.500 152.950 69.640 155.690 ;
        RECT 69.890 155.495 70.170 155.865 ;
        RECT 69.960 154.310 70.100 155.495 ;
        RECT 71.740 155.350 72.000 155.670 ;
        RECT 71.800 154.310 71.940 155.350 ;
        RECT 72.260 154.310 72.400 156.710 ;
        RECT 74.960 155.865 75.220 156.010 ;
        RECT 74.950 155.495 75.230 155.865 ;
        RECT 72.660 155.010 72.920 155.330 ;
        RECT 74.960 155.010 75.220 155.330 ;
        RECT 69.900 153.990 70.160 154.310 ;
        RECT 71.740 153.990 72.000 154.310 ;
        RECT 72.200 153.990 72.460 154.310 ;
        RECT 68.980 152.630 69.240 152.950 ;
        RECT 69.440 152.630 69.700 152.950 ;
        RECT 71.800 152.610 71.940 153.990 ;
        RECT 72.260 153.630 72.400 153.990 ;
        RECT 72.720 153.630 72.860 155.010 ;
        RECT 73.040 154.475 74.580 154.845 ;
        RECT 74.500 153.650 74.760 153.970 ;
        RECT 72.200 153.310 72.460 153.630 ;
        RECT 72.660 153.310 72.920 153.630 ;
        RECT 71.740 152.290 72.000 152.610 ;
        RECT 71.800 150.570 71.940 152.290 ;
        RECT 72.260 151.590 72.400 153.310 ;
        RECT 73.110 152.775 73.390 153.145 ;
        RECT 73.120 152.630 73.380 152.775 ;
        RECT 74.560 151.590 74.700 153.650 ;
        RECT 75.020 151.590 75.160 155.010 ;
        RECT 75.480 153.630 75.620 159.430 ;
        RECT 75.880 157.730 76.140 158.050 ;
        RECT 75.940 156.350 76.080 157.730 ;
        RECT 77.720 156.710 77.980 157.030 ;
        RECT 75.880 156.030 76.140 156.350 ;
        RECT 77.780 156.010 77.920 156.710 ;
        RECT 77.260 155.690 77.520 156.010 ;
        RECT 77.720 155.690 77.980 156.010 ;
        RECT 77.320 154.310 77.460 155.690 ;
        RECT 77.260 153.990 77.520 154.310 ;
        RECT 75.420 153.310 75.680 153.630 ;
        RECT 72.200 151.270 72.460 151.590 ;
        RECT 74.500 151.270 74.760 151.590 ;
        RECT 74.960 151.270 75.220 151.590 ;
        RECT 67.600 150.250 67.860 150.570 ;
        RECT 68.060 150.250 68.320 150.570 ;
        RECT 71.740 150.250 72.000 150.570 ;
        RECT 74.960 150.250 75.220 150.570 ;
        RECT 66.680 148.550 66.940 148.870 ;
        RECT 61.160 147.870 61.420 148.190 ;
        RECT 62.540 147.870 62.800 148.190 ;
        RECT 61.220 147.590 61.360 147.870 ;
        RECT 60.760 147.510 61.360 147.590 ;
        RECT 60.700 147.450 61.360 147.510 ;
        RECT 60.700 147.190 60.960 147.450 ;
        RECT 63.785 146.315 65.325 146.685 ;
        RECT 48.740 144.810 49.000 145.130 ;
        RECT 53.340 144.810 53.600 145.130 ;
        RECT 56.560 144.810 56.820 145.130 ;
        RECT 60.240 144.810 60.500 145.130 ;
        RECT 45.060 144.470 45.320 144.790 ;
        RECT 45.120 143.430 45.260 144.470 ;
        RECT 50.120 144.130 50.380 144.450 ;
        RECT 45.060 143.110 45.320 143.430 ;
        RECT 50.180 142.750 50.320 144.130 ;
        RECT 54.530 143.595 56.070 143.965 ;
        RECT 66.740 142.750 66.880 148.550 ;
        RECT 68.120 148.530 68.260 150.250 ;
        RECT 71.800 148.870 71.940 150.250 ;
        RECT 72.200 149.570 72.460 149.890 ;
        RECT 71.740 148.550 72.000 148.870 ;
        RECT 68.060 148.210 68.320 148.530 ;
        RECT 70.360 146.850 70.620 147.170 ;
        RECT 67.140 144.470 67.400 144.790 ;
        RECT 67.200 143.430 67.340 144.470 ;
        RECT 67.140 143.110 67.400 143.430 ;
        RECT 70.420 142.750 70.560 146.850 ;
        RECT 71.800 146.150 71.940 148.550 ;
        RECT 72.260 148.190 72.400 149.570 ;
        RECT 73.040 149.035 74.580 149.405 ;
        RECT 75.020 148.870 75.160 150.250 ;
        RECT 74.960 148.550 75.220 148.870 ;
        RECT 72.200 147.870 72.460 148.190 ;
        RECT 71.740 145.830 72.000 146.150 ;
        RECT 75.480 145.470 75.620 153.310 ;
        RECT 80.080 150.570 80.220 161.130 ;
        RECT 80.540 158.730 80.680 161.810 ;
        RECT 81.000 161.450 81.140 164.190 ;
        RECT 81.400 163.170 81.660 163.490 ;
        RECT 81.460 161.450 81.600 163.170 ;
        RECT 80.940 161.130 81.200 161.450 ;
        RECT 81.400 161.130 81.660 161.450 ;
        RECT 81.920 158.730 82.060 164.530 ;
        RECT 84.160 163.850 84.420 164.170 ;
        RECT 82.295 162.635 83.835 163.005 ;
        RECT 84.220 162.470 84.360 163.850 ;
        RECT 84.160 162.150 84.420 162.470 ;
        RECT 85.140 161.450 85.280 164.870 ;
        RECT 86.060 164.510 86.200 177.450 ;
        RECT 90.200 175.470 90.340 177.450 ;
        RECT 90.660 176.070 90.800 208.180 ;
        RECT 91.550 203.435 93.090 203.805 ;
        RECT 91.050 202.415 91.330 202.785 ;
        RECT 91.120 199.530 91.260 202.415 ;
        RECT 91.060 199.210 91.320 199.530 ;
        RECT 91.120 197.830 91.260 199.210 ;
        RECT 91.550 197.995 93.090 198.365 ;
        RECT 91.060 197.510 91.320 197.830 ;
        RECT 91.060 193.770 91.320 194.090 ;
        RECT 91.120 192.050 91.260 193.770 ;
        RECT 91.550 192.555 93.090 192.925 ;
        RECT 91.060 191.905 91.320 192.050 ;
        RECT 91.050 191.535 91.330 191.905 ;
        RECT 91.550 187.115 93.090 187.485 ;
        RECT 91.060 185.610 91.320 185.930 ;
        RECT 91.120 185.250 91.260 185.610 ;
        RECT 91.060 184.930 91.320 185.250 ;
        RECT 91.120 183.745 91.260 184.930 ;
        RECT 91.050 183.375 91.330 183.745 ;
        RECT 91.550 181.675 93.090 182.045 ;
        RECT 91.050 180.655 91.330 181.025 ;
        RECT 91.120 179.810 91.260 180.655 ;
        RECT 91.060 179.490 91.320 179.810 ;
        RECT 90.600 175.750 90.860 176.070 ;
        RECT 90.200 175.330 90.800 175.470 ;
        RECT 90.660 174.370 90.800 175.330 ;
        RECT 90.600 174.050 90.860 174.370 ;
        RECT 91.120 174.225 91.260 179.490 ;
        RECT 91.550 176.235 93.090 176.605 ;
        RECT 90.660 172.670 90.800 174.050 ;
        RECT 91.050 173.855 91.330 174.225 ;
        RECT 90.600 172.350 90.860 172.670 ;
        RECT 90.140 166.570 90.400 166.890 ;
        RECT 86.000 164.190 86.260 164.510 ;
        RECT 90.200 163.910 90.340 166.570 ;
        RECT 90.660 164.705 90.800 172.350 ;
        RECT 91.060 172.010 91.320 172.330 ;
        RECT 91.120 168.930 91.260 172.010 ;
        RECT 91.550 170.795 93.090 171.165 ;
        RECT 91.060 168.610 91.320 168.930 ;
        RECT 90.590 164.335 90.870 164.705 ;
        RECT 87.840 163.510 88.100 163.830 ;
        RECT 90.200 163.770 90.800 163.910 ;
        RECT 85.080 161.130 85.340 161.450 ;
        RECT 80.480 158.410 80.740 158.730 ;
        RECT 81.860 158.410 82.120 158.730 ;
        RECT 87.900 158.050 88.040 163.510 ;
        RECT 90.660 163.490 90.800 163.770 ;
        RECT 90.600 163.170 90.860 163.490 ;
        RECT 87.840 157.730 88.100 158.050 ;
        RECT 82.295 157.195 83.835 157.565 ;
        RECT 82.320 155.350 82.580 155.670 ;
        RECT 82.380 154.310 82.520 155.350 ;
        RECT 82.320 153.990 82.580 154.310 ;
        RECT 82.295 151.755 83.835 152.125 ;
        RECT 80.020 150.250 80.280 150.570 ;
        RECT 82.295 146.315 83.835 146.685 ;
        RECT 87.900 145.665 88.040 157.730 ;
        RECT 75.420 145.150 75.680 145.470 ;
        RECT 87.830 145.295 88.110 145.665 ;
        RECT 73.040 143.595 74.580 143.965 ;
        RECT 44.600 142.430 44.860 142.750 ;
        RECT 50.120 142.430 50.380 142.750 ;
        RECT 66.680 142.430 66.940 142.750 ;
        RECT 70.360 142.430 70.620 142.750 ;
        RECT 26.765 140.875 28.305 141.245 ;
        RECT 45.275 140.875 46.815 141.245 ;
        RECT 63.785 140.875 65.325 141.245 ;
        RECT 82.295 140.875 83.835 141.245 ;
        RECT 36.020 138.155 37.560 138.525 ;
        RECT 54.530 138.155 56.070 138.525 ;
        RECT 73.040 138.155 74.580 138.525 ;
        RECT 90.660 136.145 90.800 163.170 ;
        RECT 91.120 157.905 91.260 168.610 ;
        RECT 91.550 165.355 93.090 165.725 ;
        RECT 91.550 159.915 93.090 160.285 ;
        RECT 91.050 157.535 91.330 157.905 ;
        RECT 91.550 154.475 93.090 154.845 ;
        RECT 91.550 149.035 93.090 149.405 ;
        RECT 131.200 148.780 131.805 148.805 ;
        RECT 131.180 148.225 131.825 148.780 ;
        RECT 113.200 147.475 113.800 147.500 ;
        RECT 116.400 147.475 117.000 147.500 ;
        RECT 119.300 147.475 119.900 147.500 ;
        RECT 122.300 147.475 122.900 147.500 ;
        RECT 125.300 147.475 125.900 147.500 ;
        RECT 128.300 147.475 128.900 147.500 ;
        RECT 113.180 146.925 113.820 147.475 ;
        RECT 116.380 146.925 117.020 147.475 ;
        RECT 119.280 146.925 119.920 147.475 ;
        RECT 122.280 146.925 122.920 147.475 ;
        RECT 125.280 146.925 125.920 147.475 ;
        RECT 128.280 146.925 128.920 147.475 ;
        RECT 131.200 146.970 131.805 148.225 ;
        RECT 107.325 145.830 107.875 145.850 ;
        RECT 107.300 145.230 109.330 145.830 ;
        RECT 113.200 145.770 113.800 146.925 ;
        RECT 116.400 145.870 117.000 146.925 ;
        RECT 119.300 145.970 119.900 146.925 ;
        RECT 122.300 145.870 122.900 146.925 ;
        RECT 125.300 145.870 125.900 146.925 ;
        RECT 128.300 145.870 128.900 146.925 ;
        RECT 107.325 145.210 107.875 145.230 ;
        RECT 91.550 143.595 93.090 143.965 ;
        RECT 91.550 138.155 93.090 138.525 ;
        RECT 26.765 135.435 28.305 135.805 ;
        RECT 45.275 135.435 46.815 135.805 ;
        RECT 63.785 135.435 65.325 135.805 ;
        RECT 82.295 135.435 83.835 135.805 ;
        RECT 90.590 135.775 90.870 136.145 ;
        RECT 36.020 132.715 37.560 133.085 ;
        RECT 54.530 132.715 56.070 133.085 ;
        RECT 73.040 132.715 74.580 133.085 ;
        RECT 91.550 132.715 93.090 133.085 ;
        RECT 103.000 81.975 104.000 82.000 ;
        RECT 102.980 81.025 104.020 81.975 ;
        RECT 103.000 77.670 104.000 81.025 ;
        RECT 137.870 35.700 138.530 36.300 ;
        RECT 137.900 26.400 138.500 35.700 ;
        RECT 147.325 26.400 147.875 26.420 ;
        RECT 137.900 25.800 147.900 26.400 ;
        RECT 147.325 25.780 147.875 25.800 ;
      LAYER via2 ;
        RECT 19.740 222.390 20.040 222.690 ;
        RECT 26.260 221.415 26.540 221.695 ;
        RECT 32.620 220.445 32.920 220.745 ;
        RECT 39.055 219.375 39.335 219.655 ;
        RECT 45.480 218.210 45.760 218.490 ;
        RECT 51.940 216.960 52.240 217.260 ;
        RECT 58.410 215.730 58.690 216.010 ;
        RECT 64.820 214.760 65.120 215.060 ;
        RECT 71.220 213.650 71.500 213.930 ;
        RECT 77.700 212.670 78.000 212.970 ;
        RECT 84.140 211.705 84.420 211.985 ;
        RECT 90.580 210.720 90.880 211.020 ;
        RECT 26.795 206.200 27.075 206.480 ;
        RECT 27.195 206.200 27.475 206.480 ;
        RECT 27.595 206.200 27.875 206.480 ;
        RECT 27.995 206.200 28.275 206.480 ;
        RECT 36.050 203.480 36.330 203.760 ;
        RECT 36.450 203.480 36.730 203.760 ;
        RECT 36.850 203.480 37.130 203.760 ;
        RECT 37.250 203.480 37.530 203.760 ;
        RECT 26.795 200.760 27.075 201.040 ;
        RECT 27.195 200.760 27.475 201.040 ;
        RECT 27.595 200.760 27.875 201.040 ;
        RECT 27.995 200.760 28.275 201.040 ;
        RECT 36.050 198.040 36.330 198.320 ;
        RECT 36.450 198.040 36.730 198.320 ;
        RECT 36.850 198.040 37.130 198.320 ;
        RECT 37.250 198.040 37.530 198.320 ;
        RECT 26.795 195.320 27.075 195.600 ;
        RECT 27.195 195.320 27.475 195.600 ;
        RECT 27.595 195.320 27.875 195.600 ;
        RECT 27.995 195.320 28.275 195.600 ;
        RECT 26.795 189.880 27.075 190.160 ;
        RECT 27.195 189.880 27.475 190.160 ;
        RECT 27.595 189.880 27.875 190.160 ;
        RECT 27.995 189.880 28.275 190.160 ;
        RECT 36.050 192.600 36.330 192.880 ;
        RECT 36.450 192.600 36.730 192.880 ;
        RECT 36.850 192.600 37.130 192.880 ;
        RECT 37.250 192.600 37.530 192.880 ;
        RECT 36.050 187.160 36.330 187.440 ;
        RECT 36.450 187.160 36.730 187.440 ;
        RECT 36.850 187.160 37.130 187.440 ;
        RECT 37.250 187.160 37.530 187.440 ;
        RECT 26.795 184.440 27.075 184.720 ;
        RECT 27.195 184.440 27.475 184.720 ;
        RECT 27.595 184.440 27.875 184.720 ;
        RECT 27.995 184.440 28.275 184.720 ;
        RECT 36.050 181.720 36.330 182.000 ;
        RECT 36.450 181.720 36.730 182.000 ;
        RECT 36.850 181.720 37.130 182.000 ;
        RECT 37.250 181.720 37.530 182.000 ;
        RECT 26.795 179.000 27.075 179.280 ;
        RECT 27.195 179.000 27.475 179.280 ;
        RECT 27.595 179.000 27.875 179.280 ;
        RECT 27.995 179.000 28.275 179.280 ;
        RECT 45.305 206.200 45.585 206.480 ;
        RECT 45.705 206.200 45.985 206.480 ;
        RECT 46.105 206.200 46.385 206.480 ;
        RECT 46.505 206.200 46.785 206.480 ;
        RECT 63.815 206.200 64.095 206.480 ;
        RECT 64.215 206.200 64.495 206.480 ;
        RECT 64.615 206.200 64.895 206.480 ;
        RECT 65.015 206.200 65.295 206.480 ;
        RECT 45.305 200.760 45.585 201.040 ;
        RECT 45.705 200.760 45.985 201.040 ;
        RECT 46.105 200.760 46.385 201.040 ;
        RECT 46.505 200.760 46.785 201.040 ;
        RECT 45.305 195.320 45.585 195.600 ;
        RECT 45.705 195.320 45.985 195.600 ;
        RECT 46.105 195.320 46.385 195.600 ;
        RECT 46.505 195.320 46.785 195.600 ;
        RECT 45.305 189.880 45.585 190.160 ;
        RECT 45.705 189.880 45.985 190.160 ;
        RECT 46.105 189.880 46.385 190.160 ;
        RECT 46.505 189.880 46.785 190.160 ;
        RECT 45.305 184.440 45.585 184.720 ;
        RECT 45.705 184.440 45.985 184.720 ;
        RECT 46.105 184.440 46.385 184.720 ;
        RECT 46.505 184.440 46.785 184.720 ;
        RECT 54.560 203.480 54.840 203.760 ;
        RECT 54.960 203.480 55.240 203.760 ;
        RECT 55.360 203.480 55.640 203.760 ;
        RECT 55.760 203.480 56.040 203.760 ;
        RECT 54.560 198.040 54.840 198.320 ;
        RECT 54.960 198.040 55.240 198.320 ;
        RECT 55.360 198.040 55.640 198.320 ;
        RECT 55.760 198.040 56.040 198.320 ;
        RECT 54.560 192.600 54.840 192.880 ;
        RECT 54.960 192.600 55.240 192.880 ;
        RECT 55.360 192.600 55.640 192.880 ;
        RECT 55.760 192.600 56.040 192.880 ;
        RECT 36.050 176.280 36.330 176.560 ;
        RECT 36.450 176.280 36.730 176.560 ;
        RECT 36.850 176.280 37.130 176.560 ;
        RECT 37.250 176.280 37.530 176.560 ;
        RECT 45.305 179.000 45.585 179.280 ;
        RECT 45.705 179.000 45.985 179.280 ;
        RECT 46.105 179.000 46.385 179.280 ;
        RECT 46.505 179.000 46.785 179.280 ;
        RECT 26.795 173.560 27.075 173.840 ;
        RECT 27.195 173.560 27.475 173.840 ;
        RECT 27.595 173.560 27.875 173.840 ;
        RECT 27.995 173.560 28.275 173.840 ;
        RECT 36.050 170.840 36.330 171.120 ;
        RECT 36.450 170.840 36.730 171.120 ;
        RECT 36.850 170.840 37.130 171.120 ;
        RECT 37.250 170.840 37.530 171.120 ;
        RECT 26.795 168.120 27.075 168.400 ;
        RECT 27.195 168.120 27.475 168.400 ;
        RECT 27.595 168.120 27.875 168.400 ;
        RECT 27.995 168.120 28.275 168.400 ;
        RECT 36.050 165.400 36.330 165.680 ;
        RECT 36.450 165.400 36.730 165.680 ;
        RECT 36.850 165.400 37.130 165.680 ;
        RECT 37.250 165.400 37.530 165.680 ;
        RECT 26.795 162.680 27.075 162.960 ;
        RECT 27.195 162.680 27.475 162.960 ;
        RECT 27.595 162.680 27.875 162.960 ;
        RECT 27.995 162.680 28.275 162.960 ;
        RECT 36.050 159.960 36.330 160.240 ;
        RECT 36.450 159.960 36.730 160.240 ;
        RECT 36.850 159.960 37.130 160.240 ;
        RECT 37.250 159.960 37.530 160.240 ;
        RECT 26.795 157.240 27.075 157.520 ;
        RECT 27.195 157.240 27.475 157.520 ;
        RECT 27.595 157.240 27.875 157.520 ;
        RECT 27.995 157.240 28.275 157.520 ;
        RECT 36.050 154.520 36.330 154.800 ;
        RECT 36.450 154.520 36.730 154.800 ;
        RECT 36.850 154.520 37.130 154.800 ;
        RECT 37.250 154.520 37.530 154.800 ;
        RECT 26.795 151.800 27.075 152.080 ;
        RECT 27.195 151.800 27.475 152.080 ;
        RECT 27.595 151.800 27.875 152.080 ;
        RECT 27.995 151.800 28.275 152.080 ;
        RECT 45.305 173.560 45.585 173.840 ;
        RECT 45.705 173.560 45.985 173.840 ;
        RECT 46.105 173.560 46.385 173.840 ;
        RECT 46.505 173.560 46.785 173.840 ;
        RECT 54.560 187.160 54.840 187.440 ;
        RECT 54.960 187.160 55.240 187.440 ;
        RECT 55.360 187.160 55.640 187.440 ;
        RECT 55.760 187.160 56.040 187.440 ;
        RECT 45.305 168.120 45.585 168.400 ;
        RECT 45.705 168.120 45.985 168.400 ;
        RECT 46.105 168.120 46.385 168.400 ;
        RECT 46.505 168.120 46.785 168.400 ;
        RECT 54.560 181.720 54.840 182.000 ;
        RECT 54.960 181.720 55.240 182.000 ;
        RECT 55.360 181.720 55.640 182.000 ;
        RECT 55.760 181.720 56.040 182.000 ;
        RECT 54.560 176.280 54.840 176.560 ;
        RECT 54.960 176.280 55.240 176.560 ;
        RECT 55.360 176.280 55.640 176.560 ;
        RECT 55.760 176.280 56.040 176.560 ;
        RECT 45.305 162.680 45.585 162.960 ;
        RECT 45.705 162.680 45.985 162.960 ;
        RECT 46.105 162.680 46.385 162.960 ;
        RECT 46.505 162.680 46.785 162.960 ;
        RECT 45.305 157.240 45.585 157.520 ;
        RECT 45.705 157.240 45.985 157.520 ;
        RECT 46.105 157.240 46.385 157.520 ;
        RECT 46.505 157.240 46.785 157.520 ;
        RECT 36.050 149.080 36.330 149.360 ;
        RECT 36.450 149.080 36.730 149.360 ;
        RECT 36.850 149.080 37.130 149.360 ;
        RECT 37.250 149.080 37.530 149.360 ;
        RECT 26.795 146.360 27.075 146.640 ;
        RECT 27.195 146.360 27.475 146.640 ;
        RECT 27.595 146.360 27.875 146.640 ;
        RECT 27.995 146.360 28.275 146.640 ;
        RECT 36.050 143.640 36.330 143.920 ;
        RECT 36.450 143.640 36.730 143.920 ;
        RECT 36.850 143.640 37.130 143.920 ;
        RECT 37.250 143.640 37.530 143.920 ;
        RECT 45.305 151.800 45.585 152.080 ;
        RECT 45.705 151.800 45.985 152.080 ;
        RECT 46.105 151.800 46.385 152.080 ;
        RECT 46.505 151.800 46.785 152.080 ;
        RECT 54.560 170.840 54.840 171.120 ;
        RECT 54.960 170.840 55.240 171.120 ;
        RECT 55.360 170.840 55.640 171.120 ;
        RECT 55.760 170.840 56.040 171.120 ;
        RECT 63.815 200.760 64.095 201.040 ;
        RECT 64.215 200.760 64.495 201.040 ;
        RECT 64.615 200.760 64.895 201.040 ;
        RECT 65.015 200.760 65.295 201.040 ;
        RECT 63.815 195.320 64.095 195.600 ;
        RECT 64.215 195.320 64.495 195.600 ;
        RECT 64.615 195.320 64.895 195.600 ;
        RECT 65.015 195.320 65.295 195.600 ;
        RECT 82.325 206.200 82.605 206.480 ;
        RECT 82.725 206.200 83.005 206.480 ;
        RECT 83.125 206.200 83.405 206.480 ;
        RECT 83.525 206.200 83.805 206.480 ;
        RECT 73.070 203.480 73.350 203.760 ;
        RECT 73.470 203.480 73.750 203.760 ;
        RECT 73.870 203.480 74.150 203.760 ;
        RECT 74.270 203.480 74.550 203.760 ;
        RECT 63.815 189.880 64.095 190.160 ;
        RECT 64.215 189.880 64.495 190.160 ;
        RECT 64.615 189.880 64.895 190.160 ;
        RECT 65.015 189.880 65.295 190.160 ;
        RECT 63.815 184.440 64.095 184.720 ;
        RECT 64.215 184.440 64.495 184.720 ;
        RECT 64.615 184.440 64.895 184.720 ;
        RECT 65.015 184.440 65.295 184.720 ;
        RECT 54.560 165.400 54.840 165.680 ;
        RECT 54.960 165.400 55.240 165.680 ;
        RECT 55.360 165.400 55.640 165.680 ;
        RECT 55.760 165.400 56.040 165.680 ;
        RECT 52.870 160.980 53.150 161.260 ;
        RECT 54.250 160.980 54.530 161.260 ;
        RECT 54.560 159.960 54.840 160.240 ;
        RECT 54.960 159.960 55.240 160.240 ;
        RECT 55.360 159.960 55.640 160.240 ;
        RECT 55.760 159.960 56.040 160.240 ;
        RECT 63.815 179.000 64.095 179.280 ;
        RECT 64.215 179.000 64.495 179.280 ;
        RECT 64.615 179.000 64.895 179.280 ;
        RECT 65.015 179.000 65.295 179.280 ;
        RECT 63.815 173.560 64.095 173.840 ;
        RECT 64.215 173.560 64.495 173.840 ;
        RECT 64.615 173.560 64.895 173.840 ;
        RECT 65.015 173.560 65.295 173.840 ;
        RECT 63.815 168.120 64.095 168.400 ;
        RECT 64.215 168.120 64.495 168.400 ;
        RECT 64.615 168.120 64.895 168.400 ;
        RECT 65.015 168.120 65.295 168.400 ;
        RECT 71.730 177.300 72.010 177.580 ;
        RECT 63.815 162.680 64.095 162.960 ;
        RECT 64.215 162.680 64.495 162.960 ;
        RECT 64.615 162.680 64.895 162.960 ;
        RECT 65.015 162.680 65.295 162.960 ;
        RECT 63.815 157.240 64.095 157.520 ;
        RECT 64.215 157.240 64.495 157.520 ;
        RECT 64.615 157.240 64.895 157.520 ;
        RECT 65.015 157.240 65.295 157.520 ;
        RECT 54.560 154.520 54.840 154.800 ;
        RECT 54.960 154.520 55.240 154.800 ;
        RECT 55.360 154.520 55.640 154.800 ;
        RECT 55.760 154.520 56.040 154.800 ;
        RECT 54.560 149.080 54.840 149.360 ;
        RECT 54.960 149.080 55.240 149.360 ;
        RECT 55.360 149.080 55.640 149.360 ;
        RECT 55.760 149.080 56.040 149.360 ;
        RECT 45.305 146.360 45.585 146.640 ;
        RECT 45.705 146.360 45.985 146.640 ;
        RECT 46.105 146.360 46.385 146.640 ;
        RECT 46.505 146.360 46.785 146.640 ;
        RECT 63.815 151.800 64.095 152.080 ;
        RECT 64.215 151.800 64.495 152.080 ;
        RECT 64.615 151.800 64.895 152.080 ;
        RECT 65.015 151.800 65.295 152.080 ;
        RECT 67.590 152.820 67.870 153.100 ;
        RECT 73.070 198.040 73.350 198.320 ;
        RECT 73.470 198.040 73.750 198.320 ;
        RECT 73.870 198.040 74.150 198.320 ;
        RECT 74.270 198.040 74.550 198.320 ;
        RECT 73.070 192.600 73.350 192.880 ;
        RECT 73.470 192.600 73.750 192.880 ;
        RECT 73.870 192.600 74.150 192.880 ;
        RECT 74.270 192.600 74.550 192.880 ;
        RECT 73.070 187.160 73.350 187.440 ;
        RECT 73.470 187.160 73.750 187.440 ;
        RECT 73.870 187.160 74.150 187.440 ;
        RECT 74.270 187.160 74.550 187.440 ;
        RECT 73.070 181.720 73.350 182.000 ;
        RECT 73.470 181.720 73.750 182.000 ;
        RECT 73.870 181.720 74.150 182.000 ;
        RECT 74.270 181.720 74.550 182.000 ;
        RECT 77.250 199.060 77.530 199.340 ;
        RECT 82.325 200.760 82.605 201.040 ;
        RECT 82.725 200.760 83.005 201.040 ;
        RECT 83.125 200.760 83.405 201.040 ;
        RECT 83.525 200.760 83.805 201.040 ;
        RECT 73.070 176.280 73.350 176.560 ;
        RECT 73.470 176.280 73.750 176.560 ;
        RECT 73.870 176.280 74.150 176.560 ;
        RECT 74.270 176.280 74.550 176.560 ;
        RECT 80.010 180.700 80.290 180.980 ;
        RECT 79.550 180.020 79.830 180.300 ;
        RECT 73.070 170.840 73.350 171.120 ;
        RECT 73.470 170.840 73.750 171.120 ;
        RECT 73.870 170.840 74.150 171.120 ;
        RECT 74.270 170.840 74.550 171.120 ;
        RECT 73.070 165.400 73.350 165.680 ;
        RECT 73.470 165.400 73.750 165.680 ;
        RECT 73.870 165.400 74.150 165.680 ;
        RECT 74.270 165.400 74.550 165.680 ;
        RECT 82.325 195.320 82.605 195.600 ;
        RECT 82.725 195.320 83.005 195.600 ;
        RECT 83.125 195.320 83.405 195.600 ;
        RECT 83.525 195.320 83.805 195.600 ;
        RECT 87.830 199.060 88.110 199.340 ;
        RECT 82.325 189.880 82.605 190.160 ;
        RECT 82.725 189.880 83.005 190.160 ;
        RECT 83.125 189.880 83.405 190.160 ;
        RECT 83.525 189.880 83.805 190.160 ;
        RECT 82.325 184.440 82.605 184.720 ;
        RECT 82.725 184.440 83.005 184.720 ;
        RECT 83.125 184.440 83.405 184.720 ;
        RECT 83.525 184.440 83.805 184.720 ;
        RECT 81.390 177.300 81.670 177.580 ;
        RECT 82.770 180.020 83.050 180.300 ;
        RECT 82.325 179.000 82.605 179.280 ;
        RECT 82.725 179.000 83.005 179.280 ;
        RECT 83.125 179.000 83.405 179.280 ;
        RECT 83.525 179.000 83.805 179.280 ;
        RECT 82.325 173.560 82.605 173.840 ;
        RECT 82.725 173.560 83.005 173.840 ;
        RECT 83.125 173.560 83.405 173.840 ;
        RECT 83.525 173.560 83.805 173.840 ;
        RECT 82.325 168.120 82.605 168.400 ;
        RECT 82.725 168.120 83.005 168.400 ;
        RECT 83.125 168.120 83.405 168.400 ;
        RECT 83.525 168.120 83.805 168.400 ;
        RECT 73.070 159.960 73.350 160.240 ;
        RECT 73.470 159.960 73.750 160.240 ;
        RECT 73.870 159.960 74.150 160.240 ;
        RECT 74.270 159.960 74.550 160.240 ;
        RECT 69.890 155.540 70.170 155.820 ;
        RECT 74.950 155.540 75.230 155.820 ;
        RECT 73.070 154.520 73.350 154.800 ;
        RECT 73.470 154.520 73.750 154.800 ;
        RECT 73.870 154.520 74.150 154.800 ;
        RECT 74.270 154.520 74.550 154.800 ;
        RECT 73.110 152.820 73.390 153.100 ;
        RECT 63.815 146.360 64.095 146.640 ;
        RECT 64.215 146.360 64.495 146.640 ;
        RECT 64.615 146.360 64.895 146.640 ;
        RECT 65.015 146.360 65.295 146.640 ;
        RECT 54.560 143.640 54.840 143.920 ;
        RECT 54.960 143.640 55.240 143.920 ;
        RECT 55.360 143.640 55.640 143.920 ;
        RECT 55.760 143.640 56.040 143.920 ;
        RECT 73.070 149.080 73.350 149.360 ;
        RECT 73.470 149.080 73.750 149.360 ;
        RECT 73.870 149.080 74.150 149.360 ;
        RECT 74.270 149.080 74.550 149.360 ;
        RECT 82.325 162.680 82.605 162.960 ;
        RECT 82.725 162.680 83.005 162.960 ;
        RECT 83.125 162.680 83.405 162.960 ;
        RECT 83.525 162.680 83.805 162.960 ;
        RECT 91.580 203.480 91.860 203.760 ;
        RECT 91.980 203.480 92.260 203.760 ;
        RECT 92.380 203.480 92.660 203.760 ;
        RECT 92.780 203.480 93.060 203.760 ;
        RECT 91.050 202.460 91.330 202.740 ;
        RECT 91.580 198.040 91.860 198.320 ;
        RECT 91.980 198.040 92.260 198.320 ;
        RECT 92.380 198.040 92.660 198.320 ;
        RECT 92.780 198.040 93.060 198.320 ;
        RECT 91.580 192.600 91.860 192.880 ;
        RECT 91.980 192.600 92.260 192.880 ;
        RECT 92.380 192.600 92.660 192.880 ;
        RECT 92.780 192.600 93.060 192.880 ;
        RECT 91.050 191.580 91.330 191.860 ;
        RECT 91.580 187.160 91.860 187.440 ;
        RECT 91.980 187.160 92.260 187.440 ;
        RECT 92.380 187.160 92.660 187.440 ;
        RECT 92.780 187.160 93.060 187.440 ;
        RECT 91.050 183.420 91.330 183.700 ;
        RECT 91.580 181.720 91.860 182.000 ;
        RECT 91.980 181.720 92.260 182.000 ;
        RECT 92.380 181.720 92.660 182.000 ;
        RECT 92.780 181.720 93.060 182.000 ;
        RECT 91.050 180.700 91.330 180.980 ;
        RECT 91.580 176.280 91.860 176.560 ;
        RECT 91.980 176.280 92.260 176.560 ;
        RECT 92.380 176.280 92.660 176.560 ;
        RECT 92.780 176.280 93.060 176.560 ;
        RECT 91.050 173.900 91.330 174.180 ;
        RECT 91.580 170.840 91.860 171.120 ;
        RECT 91.980 170.840 92.260 171.120 ;
        RECT 92.380 170.840 92.660 171.120 ;
        RECT 92.780 170.840 93.060 171.120 ;
        RECT 90.590 164.380 90.870 164.660 ;
        RECT 82.325 157.240 82.605 157.520 ;
        RECT 82.725 157.240 83.005 157.520 ;
        RECT 83.125 157.240 83.405 157.520 ;
        RECT 83.525 157.240 83.805 157.520 ;
        RECT 82.325 151.800 82.605 152.080 ;
        RECT 82.725 151.800 83.005 152.080 ;
        RECT 83.125 151.800 83.405 152.080 ;
        RECT 83.525 151.800 83.805 152.080 ;
        RECT 82.325 146.360 82.605 146.640 ;
        RECT 82.725 146.360 83.005 146.640 ;
        RECT 83.125 146.360 83.405 146.640 ;
        RECT 83.525 146.360 83.805 146.640 ;
        RECT 87.830 145.340 88.110 145.620 ;
        RECT 73.070 143.640 73.350 143.920 ;
        RECT 73.470 143.640 73.750 143.920 ;
        RECT 73.870 143.640 74.150 143.920 ;
        RECT 74.270 143.640 74.550 143.920 ;
        RECT 26.795 140.920 27.075 141.200 ;
        RECT 27.195 140.920 27.475 141.200 ;
        RECT 27.595 140.920 27.875 141.200 ;
        RECT 27.995 140.920 28.275 141.200 ;
        RECT 45.305 140.920 45.585 141.200 ;
        RECT 45.705 140.920 45.985 141.200 ;
        RECT 46.105 140.920 46.385 141.200 ;
        RECT 46.505 140.920 46.785 141.200 ;
        RECT 63.815 140.920 64.095 141.200 ;
        RECT 64.215 140.920 64.495 141.200 ;
        RECT 64.615 140.920 64.895 141.200 ;
        RECT 65.015 140.920 65.295 141.200 ;
        RECT 82.325 140.920 82.605 141.200 ;
        RECT 82.725 140.920 83.005 141.200 ;
        RECT 83.125 140.920 83.405 141.200 ;
        RECT 83.525 140.920 83.805 141.200 ;
        RECT 36.050 138.200 36.330 138.480 ;
        RECT 36.450 138.200 36.730 138.480 ;
        RECT 36.850 138.200 37.130 138.480 ;
        RECT 37.250 138.200 37.530 138.480 ;
        RECT 54.560 138.200 54.840 138.480 ;
        RECT 54.960 138.200 55.240 138.480 ;
        RECT 55.360 138.200 55.640 138.480 ;
        RECT 55.760 138.200 56.040 138.480 ;
        RECT 73.070 138.200 73.350 138.480 ;
        RECT 73.470 138.200 73.750 138.480 ;
        RECT 73.870 138.200 74.150 138.480 ;
        RECT 74.270 138.200 74.550 138.480 ;
        RECT 91.580 165.400 91.860 165.680 ;
        RECT 91.980 165.400 92.260 165.680 ;
        RECT 92.380 165.400 92.660 165.680 ;
        RECT 92.780 165.400 93.060 165.680 ;
        RECT 91.580 159.960 91.860 160.240 ;
        RECT 91.980 159.960 92.260 160.240 ;
        RECT 92.380 159.960 92.660 160.240 ;
        RECT 92.780 159.960 93.060 160.240 ;
        RECT 91.050 157.580 91.330 157.860 ;
        RECT 91.580 154.520 91.860 154.800 ;
        RECT 91.980 154.520 92.260 154.800 ;
        RECT 92.380 154.520 92.660 154.800 ;
        RECT 92.780 154.520 93.060 154.800 ;
        RECT 91.580 149.080 91.860 149.360 ;
        RECT 91.980 149.080 92.260 149.360 ;
        RECT 92.380 149.080 92.660 149.360 ;
        RECT 92.780 149.080 93.060 149.360 ;
        RECT 131.225 148.225 131.780 148.780 ;
        RECT 113.225 146.925 113.775 147.475 ;
        RECT 116.425 146.925 116.975 147.475 ;
        RECT 119.325 146.925 119.875 147.475 ;
        RECT 122.325 146.925 122.875 147.475 ;
        RECT 125.325 146.925 125.875 147.475 ;
        RECT 128.325 146.925 128.875 147.475 ;
        RECT 107.325 145.255 107.875 145.805 ;
        RECT 91.580 143.640 91.860 143.920 ;
        RECT 91.980 143.640 92.260 143.920 ;
        RECT 92.380 143.640 92.660 143.920 ;
        RECT 92.780 143.640 93.060 143.920 ;
        RECT 91.580 138.200 91.860 138.480 ;
        RECT 91.980 138.200 92.260 138.480 ;
        RECT 92.380 138.200 92.660 138.480 ;
        RECT 92.780 138.200 93.060 138.480 ;
        RECT 90.590 135.820 90.870 136.100 ;
        RECT 26.795 135.480 27.075 135.760 ;
        RECT 27.195 135.480 27.475 135.760 ;
        RECT 27.595 135.480 27.875 135.760 ;
        RECT 27.995 135.480 28.275 135.760 ;
        RECT 45.305 135.480 45.585 135.760 ;
        RECT 45.705 135.480 45.985 135.760 ;
        RECT 46.105 135.480 46.385 135.760 ;
        RECT 46.505 135.480 46.785 135.760 ;
        RECT 63.815 135.480 64.095 135.760 ;
        RECT 64.215 135.480 64.495 135.760 ;
        RECT 64.615 135.480 64.895 135.760 ;
        RECT 65.015 135.480 65.295 135.760 ;
        RECT 82.325 135.480 82.605 135.760 ;
        RECT 82.725 135.480 83.005 135.760 ;
        RECT 83.125 135.480 83.405 135.760 ;
        RECT 83.525 135.480 83.805 135.760 ;
        RECT 36.050 132.760 36.330 133.040 ;
        RECT 36.450 132.760 36.730 133.040 ;
        RECT 36.850 132.760 37.130 133.040 ;
        RECT 37.250 132.760 37.530 133.040 ;
        RECT 54.560 132.760 54.840 133.040 ;
        RECT 54.960 132.760 55.240 133.040 ;
        RECT 55.360 132.760 55.640 133.040 ;
        RECT 55.760 132.760 56.040 133.040 ;
        RECT 73.070 132.760 73.350 133.040 ;
        RECT 73.470 132.760 73.750 133.040 ;
        RECT 73.870 132.760 74.150 133.040 ;
        RECT 74.270 132.760 74.550 133.040 ;
        RECT 91.580 132.760 91.860 133.040 ;
        RECT 91.980 132.760 92.260 133.040 ;
        RECT 92.380 132.760 92.660 133.040 ;
        RECT 92.780 132.760 93.060 133.040 ;
        RECT 103.025 81.025 103.975 81.975 ;
        RECT 147.325 25.825 147.875 26.375 ;
      LAYER met3 ;
        RECT 19.715 222.690 20.065 222.715 ;
        RECT 114.350 222.690 114.730 222.700 ;
        RECT 19.715 222.390 114.730 222.690 ;
        RECT 19.715 222.365 20.065 222.390 ;
        RECT 114.350 222.380 114.730 222.390 ;
        RECT 26.235 221.705 26.565 221.720 ;
        RECT 118.060 221.705 118.380 221.745 ;
        RECT 26.235 221.405 118.380 221.705 ;
        RECT 26.235 221.390 26.565 221.405 ;
        RECT 118.060 221.365 118.380 221.405 ;
        RECT 32.595 220.745 32.945 220.770 ;
        RECT 121.725 220.745 122.045 220.785 ;
        RECT 32.595 220.445 122.045 220.745 ;
        RECT 32.595 220.420 32.945 220.445 ;
        RECT 121.725 220.405 122.045 220.445 ;
        RECT 39.030 219.665 39.360 219.680 ;
        RECT 125.420 219.665 125.740 219.705 ;
        RECT 39.030 219.365 125.740 219.665 ;
        RECT 39.030 219.350 39.360 219.365 ;
        RECT 125.420 219.325 125.740 219.365 ;
        RECT 45.455 218.500 45.785 218.515 ;
        RECT 129.070 218.500 129.450 218.510 ;
        RECT 45.455 218.200 129.450 218.500 ;
        RECT 45.455 218.185 45.785 218.200 ;
        RECT 129.070 218.190 129.450 218.200 ;
        RECT 51.915 217.260 52.265 217.285 ;
        RECT 132.760 217.260 133.080 217.300 ;
        RECT 51.915 216.960 133.080 217.260 ;
        RECT 51.915 216.935 52.265 216.960 ;
        RECT 132.760 216.920 133.080 216.960 ;
        RECT 58.385 216.020 58.715 216.035 ;
        RECT 136.460 216.020 136.780 216.060 ;
        RECT 58.385 215.720 136.780 216.020 ;
        RECT 58.385 215.705 58.715 215.720 ;
        RECT 136.460 215.680 136.780 215.720 ;
        RECT 64.795 215.060 65.145 215.085 ;
        RECT 140.090 215.060 140.470 215.070 ;
        RECT 64.795 214.760 140.470 215.060 ;
        RECT 64.795 214.735 65.145 214.760 ;
        RECT 140.090 214.750 140.470 214.760 ;
        RECT 71.195 213.940 71.525 213.955 ;
        RECT 143.820 213.940 144.140 213.980 ;
        RECT 71.195 213.640 144.140 213.940 ;
        RECT 71.195 213.625 71.525 213.640 ;
        RECT 143.820 213.600 144.140 213.640 ;
        RECT 77.675 212.970 78.025 212.995 ;
        RECT 147.430 212.970 147.810 212.980 ;
        RECT 77.675 212.670 147.810 212.970 ;
        RECT 77.675 212.645 78.025 212.670 ;
        RECT 147.430 212.660 147.810 212.670 ;
        RECT 84.115 211.995 84.445 212.010 ;
        RECT 151.180 211.995 151.500 212.035 ;
        RECT 84.115 211.695 151.500 211.995 ;
        RECT 84.115 211.680 84.445 211.695 ;
        RECT 151.180 211.655 151.500 211.695 ;
        RECT 90.555 211.020 90.905 211.045 ;
        RECT 154.865 211.020 155.185 211.060 ;
        RECT 90.555 210.720 155.185 211.020 ;
        RECT 90.555 210.695 90.905 210.720 ;
        RECT 154.865 210.680 155.185 210.720 ;
        RECT 26.745 206.175 28.325 206.505 ;
        RECT 45.255 206.175 46.835 206.505 ;
        RECT 63.765 206.175 65.345 206.505 ;
        RECT 82.275 206.175 83.855 206.505 ;
        RECT 36.000 203.455 37.580 203.785 ;
        RECT 54.510 203.455 56.090 203.785 ;
        RECT 73.020 203.455 74.600 203.785 ;
        RECT 91.530 203.455 93.110 203.785 ;
        RECT 91.025 202.750 91.355 202.765 ;
        RECT 93.520 202.750 131.800 202.900 ;
        RECT 91.025 202.450 131.800 202.750 ;
        RECT 91.025 202.435 91.355 202.450 ;
        RECT 93.520 202.300 131.800 202.450 ;
        RECT 26.745 200.735 28.325 201.065 ;
        RECT 45.255 200.735 46.835 201.065 ;
        RECT 63.765 200.735 65.345 201.065 ;
        RECT 82.275 200.735 83.855 201.065 ;
        RECT 77.225 199.350 77.555 199.365 ;
        RECT 87.805 199.350 88.135 199.365 ;
        RECT 77.225 199.050 88.135 199.350 ;
        RECT 77.225 199.035 77.555 199.050 ;
        RECT 87.805 199.035 88.135 199.050 ;
        RECT 36.000 198.015 37.580 198.345 ;
        RECT 54.510 198.015 56.090 198.345 ;
        RECT 73.020 198.015 74.600 198.345 ;
        RECT 91.530 198.015 93.110 198.345 ;
        RECT 26.745 195.295 28.325 195.625 ;
        RECT 45.255 195.295 46.835 195.625 ;
        RECT 63.765 195.295 65.345 195.625 ;
        RECT 82.275 195.295 83.855 195.625 ;
        RECT 36.000 192.575 37.580 192.905 ;
        RECT 54.510 192.575 56.090 192.905 ;
        RECT 73.020 192.575 74.600 192.905 ;
        RECT 91.530 192.575 93.110 192.905 ;
        RECT 93.520 192.780 128.900 193.380 ;
        RECT 91.025 191.870 91.355 191.885 ;
        RECT 94.030 191.870 94.330 192.780 ;
        RECT 91.025 191.570 94.330 191.870 ;
        RECT 91.025 191.555 91.355 191.570 ;
        RECT 26.745 189.855 28.325 190.185 ;
        RECT 45.255 189.855 46.835 190.185 ;
        RECT 63.765 189.855 65.345 190.185 ;
        RECT 82.275 189.855 83.855 190.185 ;
        RECT 36.000 187.135 37.580 187.465 ;
        RECT 54.510 187.135 56.090 187.465 ;
        RECT 73.020 187.135 74.600 187.465 ;
        RECT 91.530 187.135 93.110 187.465 ;
        RECT 26.745 184.415 28.325 184.745 ;
        RECT 45.255 184.415 46.835 184.745 ;
        RECT 63.765 184.415 65.345 184.745 ;
        RECT 82.275 184.415 83.855 184.745 ;
        RECT 91.025 183.710 91.355 183.725 ;
        RECT 93.520 183.710 125.900 183.860 ;
        RECT 91.025 183.410 125.900 183.710 ;
        RECT 91.025 183.395 91.355 183.410 ;
        RECT 93.520 183.260 125.900 183.410 ;
        RECT 36.000 181.695 37.580 182.025 ;
        RECT 54.510 181.695 56.090 182.025 ;
        RECT 73.020 181.695 74.600 182.025 ;
        RECT 91.530 181.695 93.110 182.025 ;
        RECT 79.985 180.990 80.315 181.005 ;
        RECT 91.025 180.990 91.355 181.005 ;
        RECT 79.985 180.690 91.355 180.990 ;
        RECT 79.985 180.675 80.315 180.690 ;
        RECT 91.025 180.675 91.355 180.690 ;
        RECT 79.525 180.310 79.855 180.325 ;
        RECT 82.745 180.310 83.075 180.325 ;
        RECT 79.525 180.010 83.075 180.310 ;
        RECT 79.525 179.995 79.855 180.010 ;
        RECT 82.745 179.995 83.075 180.010 ;
        RECT 26.745 178.975 28.325 179.305 ;
        RECT 45.255 178.975 46.835 179.305 ;
        RECT 63.765 178.975 65.345 179.305 ;
        RECT 82.275 178.975 83.855 179.305 ;
        RECT 71.705 177.590 72.035 177.605 ;
        RECT 81.365 177.590 81.695 177.605 ;
        RECT 71.705 177.290 81.695 177.590 ;
        RECT 71.705 177.275 72.035 177.290 ;
        RECT 81.365 177.275 81.695 177.290 ;
        RECT 36.000 176.255 37.580 176.585 ;
        RECT 54.510 176.255 56.090 176.585 ;
        RECT 73.020 176.255 74.600 176.585 ;
        RECT 91.530 176.255 93.110 176.585 ;
        RECT 91.025 174.190 91.355 174.205 ;
        RECT 93.520 174.190 122.900 174.340 ;
        RECT 91.025 173.890 122.900 174.190 ;
        RECT 91.025 173.875 91.355 173.890 ;
        RECT 26.745 173.535 28.325 173.865 ;
        RECT 45.255 173.535 46.835 173.865 ;
        RECT 63.765 173.535 65.345 173.865 ;
        RECT 82.275 173.535 83.855 173.865 ;
        RECT 93.520 173.740 122.900 173.890 ;
        RECT 36.000 170.815 37.580 171.145 ;
        RECT 54.510 170.815 56.090 171.145 ;
        RECT 73.020 170.815 74.600 171.145 ;
        RECT 91.530 170.815 93.110 171.145 ;
        RECT 26.745 168.095 28.325 168.425 ;
        RECT 45.255 168.095 46.835 168.425 ;
        RECT 63.765 168.095 65.345 168.425 ;
        RECT 82.275 168.095 83.855 168.425 ;
        RECT 36.000 165.375 37.580 165.705 ;
        RECT 54.510 165.375 56.090 165.705 ;
        RECT 73.020 165.375 74.600 165.705 ;
        RECT 91.530 165.375 93.110 165.705 ;
        RECT 90.565 164.670 90.895 164.685 ;
        RECT 93.520 164.670 119.900 164.820 ;
        RECT 90.565 164.370 119.900 164.670 ;
        RECT 90.565 164.355 90.895 164.370 ;
        RECT 93.520 164.220 119.900 164.370 ;
        RECT 26.745 162.655 28.325 162.985 ;
        RECT 45.255 162.655 46.835 162.985 ;
        RECT 63.765 162.655 65.345 162.985 ;
        RECT 82.275 162.655 83.855 162.985 ;
        RECT 52.845 161.270 53.175 161.285 ;
        RECT 54.225 161.270 54.555 161.285 ;
        RECT 52.845 160.970 54.555 161.270 ;
        RECT 52.845 160.955 53.175 160.970 ;
        RECT 54.225 160.955 54.555 160.970 ;
        RECT 36.000 159.935 37.580 160.265 ;
        RECT 54.510 159.935 56.090 160.265 ;
        RECT 73.020 159.935 74.600 160.265 ;
        RECT 91.530 159.935 93.110 160.265 ;
        RECT 91.025 157.870 91.355 157.885 ;
        RECT 91.025 157.570 94.330 157.870 ;
        RECT 91.025 157.555 91.355 157.570 ;
        RECT 26.745 157.215 28.325 157.545 ;
        RECT 45.255 157.215 46.835 157.545 ;
        RECT 63.765 157.215 65.345 157.545 ;
        RECT 82.275 157.215 83.855 157.545 ;
        RECT 69.865 155.830 70.195 155.845 ;
        RECT 74.925 155.830 75.255 155.845 ;
        RECT 69.865 155.530 75.255 155.830 ;
        RECT 69.865 155.515 70.195 155.530 ;
        RECT 74.925 155.515 75.255 155.530 ;
        RECT 94.030 155.300 94.330 157.570 ;
        RECT 36.000 154.495 37.580 154.825 ;
        RECT 54.510 154.495 56.090 154.825 ;
        RECT 73.020 154.495 74.600 154.825 ;
        RECT 91.530 154.495 93.110 154.825 ;
        RECT 93.520 154.700 117.000 155.300 ;
        RECT 67.565 153.110 67.895 153.125 ;
        RECT 73.085 153.110 73.415 153.125 ;
        RECT 67.565 152.810 73.415 153.110 ;
        RECT 67.565 152.795 67.895 152.810 ;
        RECT 73.085 152.795 73.415 152.810 ;
        RECT 26.745 151.775 28.325 152.105 ;
        RECT 45.255 151.775 46.835 152.105 ;
        RECT 63.765 151.775 65.345 152.105 ;
        RECT 82.275 151.775 83.855 152.105 ;
        RECT 36.000 149.055 37.580 149.385 ;
        RECT 54.510 149.055 56.090 149.385 ;
        RECT 73.020 149.055 74.600 149.385 ;
        RECT 91.530 149.055 93.110 149.385 ;
        RECT 99.100 148.400 113.800 149.000 ;
        RECT 26.745 146.335 28.325 146.665 ;
        RECT 45.255 146.335 46.835 146.665 ;
        RECT 63.765 146.335 65.345 146.665 ;
        RECT 82.275 146.335 83.855 146.665 ;
        RECT 99.100 145.780 99.700 148.400 ;
        RECT 113.200 146.900 113.800 148.400 ;
        RECT 116.400 146.900 117.000 154.700 ;
        RECT 119.300 146.900 119.900 164.220 ;
        RECT 122.300 146.900 122.900 173.740 ;
        RECT 125.300 146.900 125.900 183.260 ;
        RECT 128.300 146.900 128.900 192.780 ;
        RECT 131.200 148.805 131.800 202.300 ;
        RECT 131.200 148.200 131.805 148.805 ;
        RECT 87.805 145.630 88.135 145.645 ;
        RECT 93.520 145.630 99.700 145.780 ;
        RECT 87.805 145.330 99.700 145.630 ;
        RECT 87.805 145.315 88.135 145.330 ;
        RECT 93.520 145.180 99.700 145.330 ;
        RECT 104.700 145.230 107.900 145.830 ;
        RECT 36.000 143.615 37.580 143.945 ;
        RECT 54.510 143.615 56.090 143.945 ;
        RECT 73.020 143.615 74.600 143.945 ;
        RECT 91.530 143.615 93.110 143.945 ;
        RECT 26.745 140.895 28.325 141.225 ;
        RECT 45.255 140.895 46.835 141.225 ;
        RECT 63.765 140.895 65.345 141.225 ;
        RECT 82.275 140.895 83.855 141.225 ;
        RECT 36.000 138.175 37.580 138.505 ;
        RECT 54.510 138.175 56.090 138.505 ;
        RECT 73.020 138.175 74.600 138.505 ;
        RECT 91.530 138.175 93.110 138.505 ;
        RECT 104.700 136.260 105.300 145.230 ;
        RECT 90.565 136.110 90.895 136.125 ;
        RECT 93.520 136.110 105.300 136.260 ;
        RECT 90.565 135.810 105.300 136.110 ;
        RECT 90.565 135.795 90.895 135.810 ;
        RECT 26.745 135.455 28.325 135.785 ;
        RECT 45.255 135.455 46.835 135.785 ;
        RECT 63.765 135.455 65.345 135.785 ;
        RECT 82.275 135.455 83.855 135.785 ;
        RECT 93.520 135.660 105.300 135.810 ;
        RECT 36.000 132.735 37.580 133.065 ;
        RECT 54.510 132.735 56.090 133.065 ;
        RECT 73.020 132.735 74.600 133.065 ;
        RECT 91.530 132.735 93.110 133.065 ;
        RECT 26.550 126.500 28.150 126.530 ;
        RECT 63.800 126.500 65.400 126.530 ;
        RECT 0.910 124.900 83.900 126.500 ;
        RECT 26.550 124.870 28.150 124.900 ;
        RECT 63.800 124.870 65.400 124.900 ;
        RECT 103.000 121.155 104.000 121.160 ;
        RECT 102.975 120.165 104.025 121.155 ;
        RECT 103.000 81.000 104.000 120.165 ;
        RECT 156.565 26.400 157.155 26.425 ;
        RECT 147.300 25.800 157.160 26.400 ;
        RECT 156.565 25.775 157.155 25.800 ;
      LAYER via3 ;
        RECT 114.380 222.380 114.700 222.700 ;
        RECT 118.060 221.395 118.380 221.715 ;
        RECT 121.725 220.435 122.045 220.755 ;
        RECT 125.420 219.355 125.740 219.675 ;
        RECT 129.100 218.190 129.420 218.510 ;
        RECT 132.760 216.950 133.080 217.270 ;
        RECT 136.460 215.710 136.780 216.030 ;
        RECT 140.120 214.750 140.440 215.070 ;
        RECT 143.820 213.630 144.140 213.950 ;
        RECT 147.460 212.660 147.780 212.980 ;
        RECT 151.180 211.685 151.500 212.005 ;
        RECT 154.865 210.710 155.185 211.030 ;
        RECT 26.775 206.180 27.095 206.500 ;
        RECT 27.175 206.180 27.495 206.500 ;
        RECT 27.575 206.180 27.895 206.500 ;
        RECT 27.975 206.180 28.295 206.500 ;
        RECT 45.285 206.180 45.605 206.500 ;
        RECT 45.685 206.180 46.005 206.500 ;
        RECT 46.085 206.180 46.405 206.500 ;
        RECT 46.485 206.180 46.805 206.500 ;
        RECT 63.795 206.180 64.115 206.500 ;
        RECT 64.195 206.180 64.515 206.500 ;
        RECT 64.595 206.180 64.915 206.500 ;
        RECT 64.995 206.180 65.315 206.500 ;
        RECT 82.305 206.180 82.625 206.500 ;
        RECT 82.705 206.180 83.025 206.500 ;
        RECT 83.105 206.180 83.425 206.500 ;
        RECT 83.505 206.180 83.825 206.500 ;
        RECT 36.030 203.460 36.350 203.780 ;
        RECT 36.430 203.460 36.750 203.780 ;
        RECT 36.830 203.460 37.150 203.780 ;
        RECT 37.230 203.460 37.550 203.780 ;
        RECT 54.540 203.460 54.860 203.780 ;
        RECT 54.940 203.460 55.260 203.780 ;
        RECT 55.340 203.460 55.660 203.780 ;
        RECT 55.740 203.460 56.060 203.780 ;
        RECT 73.050 203.460 73.370 203.780 ;
        RECT 73.450 203.460 73.770 203.780 ;
        RECT 73.850 203.460 74.170 203.780 ;
        RECT 74.250 203.460 74.570 203.780 ;
        RECT 91.560 203.460 91.880 203.780 ;
        RECT 91.960 203.460 92.280 203.780 ;
        RECT 92.360 203.460 92.680 203.780 ;
        RECT 92.760 203.460 93.080 203.780 ;
        RECT 26.775 200.740 27.095 201.060 ;
        RECT 27.175 200.740 27.495 201.060 ;
        RECT 27.575 200.740 27.895 201.060 ;
        RECT 27.975 200.740 28.295 201.060 ;
        RECT 45.285 200.740 45.605 201.060 ;
        RECT 45.685 200.740 46.005 201.060 ;
        RECT 46.085 200.740 46.405 201.060 ;
        RECT 46.485 200.740 46.805 201.060 ;
        RECT 63.795 200.740 64.115 201.060 ;
        RECT 64.195 200.740 64.515 201.060 ;
        RECT 64.595 200.740 64.915 201.060 ;
        RECT 64.995 200.740 65.315 201.060 ;
        RECT 82.305 200.740 82.625 201.060 ;
        RECT 82.705 200.740 83.025 201.060 ;
        RECT 83.105 200.740 83.425 201.060 ;
        RECT 83.505 200.740 83.825 201.060 ;
        RECT 36.030 198.020 36.350 198.340 ;
        RECT 36.430 198.020 36.750 198.340 ;
        RECT 36.830 198.020 37.150 198.340 ;
        RECT 37.230 198.020 37.550 198.340 ;
        RECT 54.540 198.020 54.860 198.340 ;
        RECT 54.940 198.020 55.260 198.340 ;
        RECT 55.340 198.020 55.660 198.340 ;
        RECT 55.740 198.020 56.060 198.340 ;
        RECT 73.050 198.020 73.370 198.340 ;
        RECT 73.450 198.020 73.770 198.340 ;
        RECT 73.850 198.020 74.170 198.340 ;
        RECT 74.250 198.020 74.570 198.340 ;
        RECT 91.560 198.020 91.880 198.340 ;
        RECT 91.960 198.020 92.280 198.340 ;
        RECT 92.360 198.020 92.680 198.340 ;
        RECT 92.760 198.020 93.080 198.340 ;
        RECT 26.775 195.300 27.095 195.620 ;
        RECT 27.175 195.300 27.495 195.620 ;
        RECT 27.575 195.300 27.895 195.620 ;
        RECT 27.975 195.300 28.295 195.620 ;
        RECT 45.285 195.300 45.605 195.620 ;
        RECT 45.685 195.300 46.005 195.620 ;
        RECT 46.085 195.300 46.405 195.620 ;
        RECT 46.485 195.300 46.805 195.620 ;
        RECT 63.795 195.300 64.115 195.620 ;
        RECT 64.195 195.300 64.515 195.620 ;
        RECT 64.595 195.300 64.915 195.620 ;
        RECT 64.995 195.300 65.315 195.620 ;
        RECT 82.305 195.300 82.625 195.620 ;
        RECT 82.705 195.300 83.025 195.620 ;
        RECT 83.105 195.300 83.425 195.620 ;
        RECT 83.505 195.300 83.825 195.620 ;
        RECT 36.030 192.580 36.350 192.900 ;
        RECT 36.430 192.580 36.750 192.900 ;
        RECT 36.830 192.580 37.150 192.900 ;
        RECT 37.230 192.580 37.550 192.900 ;
        RECT 54.540 192.580 54.860 192.900 ;
        RECT 54.940 192.580 55.260 192.900 ;
        RECT 55.340 192.580 55.660 192.900 ;
        RECT 55.740 192.580 56.060 192.900 ;
        RECT 73.050 192.580 73.370 192.900 ;
        RECT 73.450 192.580 73.770 192.900 ;
        RECT 73.850 192.580 74.170 192.900 ;
        RECT 74.250 192.580 74.570 192.900 ;
        RECT 91.560 192.580 91.880 192.900 ;
        RECT 91.960 192.580 92.280 192.900 ;
        RECT 92.360 192.580 92.680 192.900 ;
        RECT 92.760 192.580 93.080 192.900 ;
        RECT 26.775 189.860 27.095 190.180 ;
        RECT 27.175 189.860 27.495 190.180 ;
        RECT 27.575 189.860 27.895 190.180 ;
        RECT 27.975 189.860 28.295 190.180 ;
        RECT 45.285 189.860 45.605 190.180 ;
        RECT 45.685 189.860 46.005 190.180 ;
        RECT 46.085 189.860 46.405 190.180 ;
        RECT 46.485 189.860 46.805 190.180 ;
        RECT 63.795 189.860 64.115 190.180 ;
        RECT 64.195 189.860 64.515 190.180 ;
        RECT 64.595 189.860 64.915 190.180 ;
        RECT 64.995 189.860 65.315 190.180 ;
        RECT 82.305 189.860 82.625 190.180 ;
        RECT 82.705 189.860 83.025 190.180 ;
        RECT 83.105 189.860 83.425 190.180 ;
        RECT 83.505 189.860 83.825 190.180 ;
        RECT 36.030 187.140 36.350 187.460 ;
        RECT 36.430 187.140 36.750 187.460 ;
        RECT 36.830 187.140 37.150 187.460 ;
        RECT 37.230 187.140 37.550 187.460 ;
        RECT 54.540 187.140 54.860 187.460 ;
        RECT 54.940 187.140 55.260 187.460 ;
        RECT 55.340 187.140 55.660 187.460 ;
        RECT 55.740 187.140 56.060 187.460 ;
        RECT 73.050 187.140 73.370 187.460 ;
        RECT 73.450 187.140 73.770 187.460 ;
        RECT 73.850 187.140 74.170 187.460 ;
        RECT 74.250 187.140 74.570 187.460 ;
        RECT 91.560 187.140 91.880 187.460 ;
        RECT 91.960 187.140 92.280 187.460 ;
        RECT 92.360 187.140 92.680 187.460 ;
        RECT 92.760 187.140 93.080 187.460 ;
        RECT 26.775 184.420 27.095 184.740 ;
        RECT 27.175 184.420 27.495 184.740 ;
        RECT 27.575 184.420 27.895 184.740 ;
        RECT 27.975 184.420 28.295 184.740 ;
        RECT 45.285 184.420 45.605 184.740 ;
        RECT 45.685 184.420 46.005 184.740 ;
        RECT 46.085 184.420 46.405 184.740 ;
        RECT 46.485 184.420 46.805 184.740 ;
        RECT 63.795 184.420 64.115 184.740 ;
        RECT 64.195 184.420 64.515 184.740 ;
        RECT 64.595 184.420 64.915 184.740 ;
        RECT 64.995 184.420 65.315 184.740 ;
        RECT 82.305 184.420 82.625 184.740 ;
        RECT 82.705 184.420 83.025 184.740 ;
        RECT 83.105 184.420 83.425 184.740 ;
        RECT 83.505 184.420 83.825 184.740 ;
        RECT 36.030 181.700 36.350 182.020 ;
        RECT 36.430 181.700 36.750 182.020 ;
        RECT 36.830 181.700 37.150 182.020 ;
        RECT 37.230 181.700 37.550 182.020 ;
        RECT 54.540 181.700 54.860 182.020 ;
        RECT 54.940 181.700 55.260 182.020 ;
        RECT 55.340 181.700 55.660 182.020 ;
        RECT 55.740 181.700 56.060 182.020 ;
        RECT 73.050 181.700 73.370 182.020 ;
        RECT 73.450 181.700 73.770 182.020 ;
        RECT 73.850 181.700 74.170 182.020 ;
        RECT 74.250 181.700 74.570 182.020 ;
        RECT 91.560 181.700 91.880 182.020 ;
        RECT 91.960 181.700 92.280 182.020 ;
        RECT 92.360 181.700 92.680 182.020 ;
        RECT 92.760 181.700 93.080 182.020 ;
        RECT 26.775 178.980 27.095 179.300 ;
        RECT 27.175 178.980 27.495 179.300 ;
        RECT 27.575 178.980 27.895 179.300 ;
        RECT 27.975 178.980 28.295 179.300 ;
        RECT 45.285 178.980 45.605 179.300 ;
        RECT 45.685 178.980 46.005 179.300 ;
        RECT 46.085 178.980 46.405 179.300 ;
        RECT 46.485 178.980 46.805 179.300 ;
        RECT 63.795 178.980 64.115 179.300 ;
        RECT 64.195 178.980 64.515 179.300 ;
        RECT 64.595 178.980 64.915 179.300 ;
        RECT 64.995 178.980 65.315 179.300 ;
        RECT 82.305 178.980 82.625 179.300 ;
        RECT 82.705 178.980 83.025 179.300 ;
        RECT 83.105 178.980 83.425 179.300 ;
        RECT 83.505 178.980 83.825 179.300 ;
        RECT 36.030 176.260 36.350 176.580 ;
        RECT 36.430 176.260 36.750 176.580 ;
        RECT 36.830 176.260 37.150 176.580 ;
        RECT 37.230 176.260 37.550 176.580 ;
        RECT 54.540 176.260 54.860 176.580 ;
        RECT 54.940 176.260 55.260 176.580 ;
        RECT 55.340 176.260 55.660 176.580 ;
        RECT 55.740 176.260 56.060 176.580 ;
        RECT 73.050 176.260 73.370 176.580 ;
        RECT 73.450 176.260 73.770 176.580 ;
        RECT 73.850 176.260 74.170 176.580 ;
        RECT 74.250 176.260 74.570 176.580 ;
        RECT 91.560 176.260 91.880 176.580 ;
        RECT 91.960 176.260 92.280 176.580 ;
        RECT 92.360 176.260 92.680 176.580 ;
        RECT 92.760 176.260 93.080 176.580 ;
        RECT 26.775 173.540 27.095 173.860 ;
        RECT 27.175 173.540 27.495 173.860 ;
        RECT 27.575 173.540 27.895 173.860 ;
        RECT 27.975 173.540 28.295 173.860 ;
        RECT 45.285 173.540 45.605 173.860 ;
        RECT 45.685 173.540 46.005 173.860 ;
        RECT 46.085 173.540 46.405 173.860 ;
        RECT 46.485 173.540 46.805 173.860 ;
        RECT 63.795 173.540 64.115 173.860 ;
        RECT 64.195 173.540 64.515 173.860 ;
        RECT 64.595 173.540 64.915 173.860 ;
        RECT 64.995 173.540 65.315 173.860 ;
        RECT 82.305 173.540 82.625 173.860 ;
        RECT 82.705 173.540 83.025 173.860 ;
        RECT 83.105 173.540 83.425 173.860 ;
        RECT 83.505 173.540 83.825 173.860 ;
        RECT 36.030 170.820 36.350 171.140 ;
        RECT 36.430 170.820 36.750 171.140 ;
        RECT 36.830 170.820 37.150 171.140 ;
        RECT 37.230 170.820 37.550 171.140 ;
        RECT 54.540 170.820 54.860 171.140 ;
        RECT 54.940 170.820 55.260 171.140 ;
        RECT 55.340 170.820 55.660 171.140 ;
        RECT 55.740 170.820 56.060 171.140 ;
        RECT 73.050 170.820 73.370 171.140 ;
        RECT 73.450 170.820 73.770 171.140 ;
        RECT 73.850 170.820 74.170 171.140 ;
        RECT 74.250 170.820 74.570 171.140 ;
        RECT 91.560 170.820 91.880 171.140 ;
        RECT 91.960 170.820 92.280 171.140 ;
        RECT 92.360 170.820 92.680 171.140 ;
        RECT 92.760 170.820 93.080 171.140 ;
        RECT 26.775 168.100 27.095 168.420 ;
        RECT 27.175 168.100 27.495 168.420 ;
        RECT 27.575 168.100 27.895 168.420 ;
        RECT 27.975 168.100 28.295 168.420 ;
        RECT 45.285 168.100 45.605 168.420 ;
        RECT 45.685 168.100 46.005 168.420 ;
        RECT 46.085 168.100 46.405 168.420 ;
        RECT 46.485 168.100 46.805 168.420 ;
        RECT 63.795 168.100 64.115 168.420 ;
        RECT 64.195 168.100 64.515 168.420 ;
        RECT 64.595 168.100 64.915 168.420 ;
        RECT 64.995 168.100 65.315 168.420 ;
        RECT 82.305 168.100 82.625 168.420 ;
        RECT 82.705 168.100 83.025 168.420 ;
        RECT 83.105 168.100 83.425 168.420 ;
        RECT 83.505 168.100 83.825 168.420 ;
        RECT 36.030 165.380 36.350 165.700 ;
        RECT 36.430 165.380 36.750 165.700 ;
        RECT 36.830 165.380 37.150 165.700 ;
        RECT 37.230 165.380 37.550 165.700 ;
        RECT 54.540 165.380 54.860 165.700 ;
        RECT 54.940 165.380 55.260 165.700 ;
        RECT 55.340 165.380 55.660 165.700 ;
        RECT 55.740 165.380 56.060 165.700 ;
        RECT 73.050 165.380 73.370 165.700 ;
        RECT 73.450 165.380 73.770 165.700 ;
        RECT 73.850 165.380 74.170 165.700 ;
        RECT 74.250 165.380 74.570 165.700 ;
        RECT 91.560 165.380 91.880 165.700 ;
        RECT 91.960 165.380 92.280 165.700 ;
        RECT 92.360 165.380 92.680 165.700 ;
        RECT 92.760 165.380 93.080 165.700 ;
        RECT 26.775 162.660 27.095 162.980 ;
        RECT 27.175 162.660 27.495 162.980 ;
        RECT 27.575 162.660 27.895 162.980 ;
        RECT 27.975 162.660 28.295 162.980 ;
        RECT 45.285 162.660 45.605 162.980 ;
        RECT 45.685 162.660 46.005 162.980 ;
        RECT 46.085 162.660 46.405 162.980 ;
        RECT 46.485 162.660 46.805 162.980 ;
        RECT 63.795 162.660 64.115 162.980 ;
        RECT 64.195 162.660 64.515 162.980 ;
        RECT 64.595 162.660 64.915 162.980 ;
        RECT 64.995 162.660 65.315 162.980 ;
        RECT 82.305 162.660 82.625 162.980 ;
        RECT 82.705 162.660 83.025 162.980 ;
        RECT 83.105 162.660 83.425 162.980 ;
        RECT 83.505 162.660 83.825 162.980 ;
        RECT 36.030 159.940 36.350 160.260 ;
        RECT 36.430 159.940 36.750 160.260 ;
        RECT 36.830 159.940 37.150 160.260 ;
        RECT 37.230 159.940 37.550 160.260 ;
        RECT 54.540 159.940 54.860 160.260 ;
        RECT 54.940 159.940 55.260 160.260 ;
        RECT 55.340 159.940 55.660 160.260 ;
        RECT 55.740 159.940 56.060 160.260 ;
        RECT 73.050 159.940 73.370 160.260 ;
        RECT 73.450 159.940 73.770 160.260 ;
        RECT 73.850 159.940 74.170 160.260 ;
        RECT 74.250 159.940 74.570 160.260 ;
        RECT 91.560 159.940 91.880 160.260 ;
        RECT 91.960 159.940 92.280 160.260 ;
        RECT 92.360 159.940 92.680 160.260 ;
        RECT 92.760 159.940 93.080 160.260 ;
        RECT 26.775 157.220 27.095 157.540 ;
        RECT 27.175 157.220 27.495 157.540 ;
        RECT 27.575 157.220 27.895 157.540 ;
        RECT 27.975 157.220 28.295 157.540 ;
        RECT 45.285 157.220 45.605 157.540 ;
        RECT 45.685 157.220 46.005 157.540 ;
        RECT 46.085 157.220 46.405 157.540 ;
        RECT 46.485 157.220 46.805 157.540 ;
        RECT 63.795 157.220 64.115 157.540 ;
        RECT 64.195 157.220 64.515 157.540 ;
        RECT 64.595 157.220 64.915 157.540 ;
        RECT 64.995 157.220 65.315 157.540 ;
        RECT 82.305 157.220 82.625 157.540 ;
        RECT 82.705 157.220 83.025 157.540 ;
        RECT 83.105 157.220 83.425 157.540 ;
        RECT 83.505 157.220 83.825 157.540 ;
        RECT 36.030 154.500 36.350 154.820 ;
        RECT 36.430 154.500 36.750 154.820 ;
        RECT 36.830 154.500 37.150 154.820 ;
        RECT 37.230 154.500 37.550 154.820 ;
        RECT 54.540 154.500 54.860 154.820 ;
        RECT 54.940 154.500 55.260 154.820 ;
        RECT 55.340 154.500 55.660 154.820 ;
        RECT 55.740 154.500 56.060 154.820 ;
        RECT 73.050 154.500 73.370 154.820 ;
        RECT 73.450 154.500 73.770 154.820 ;
        RECT 73.850 154.500 74.170 154.820 ;
        RECT 74.250 154.500 74.570 154.820 ;
        RECT 91.560 154.500 91.880 154.820 ;
        RECT 91.960 154.500 92.280 154.820 ;
        RECT 92.360 154.500 92.680 154.820 ;
        RECT 92.760 154.500 93.080 154.820 ;
        RECT 26.775 151.780 27.095 152.100 ;
        RECT 27.175 151.780 27.495 152.100 ;
        RECT 27.575 151.780 27.895 152.100 ;
        RECT 27.975 151.780 28.295 152.100 ;
        RECT 45.285 151.780 45.605 152.100 ;
        RECT 45.685 151.780 46.005 152.100 ;
        RECT 46.085 151.780 46.405 152.100 ;
        RECT 46.485 151.780 46.805 152.100 ;
        RECT 63.795 151.780 64.115 152.100 ;
        RECT 64.195 151.780 64.515 152.100 ;
        RECT 64.595 151.780 64.915 152.100 ;
        RECT 64.995 151.780 65.315 152.100 ;
        RECT 82.305 151.780 82.625 152.100 ;
        RECT 82.705 151.780 83.025 152.100 ;
        RECT 83.105 151.780 83.425 152.100 ;
        RECT 83.505 151.780 83.825 152.100 ;
        RECT 36.030 149.060 36.350 149.380 ;
        RECT 36.430 149.060 36.750 149.380 ;
        RECT 36.830 149.060 37.150 149.380 ;
        RECT 37.230 149.060 37.550 149.380 ;
        RECT 54.540 149.060 54.860 149.380 ;
        RECT 54.940 149.060 55.260 149.380 ;
        RECT 55.340 149.060 55.660 149.380 ;
        RECT 55.740 149.060 56.060 149.380 ;
        RECT 73.050 149.060 73.370 149.380 ;
        RECT 73.450 149.060 73.770 149.380 ;
        RECT 73.850 149.060 74.170 149.380 ;
        RECT 74.250 149.060 74.570 149.380 ;
        RECT 91.560 149.060 91.880 149.380 ;
        RECT 91.960 149.060 92.280 149.380 ;
        RECT 92.360 149.060 92.680 149.380 ;
        RECT 92.760 149.060 93.080 149.380 ;
        RECT 26.775 146.340 27.095 146.660 ;
        RECT 27.175 146.340 27.495 146.660 ;
        RECT 27.575 146.340 27.895 146.660 ;
        RECT 27.975 146.340 28.295 146.660 ;
        RECT 45.285 146.340 45.605 146.660 ;
        RECT 45.685 146.340 46.005 146.660 ;
        RECT 46.085 146.340 46.405 146.660 ;
        RECT 46.485 146.340 46.805 146.660 ;
        RECT 63.795 146.340 64.115 146.660 ;
        RECT 64.195 146.340 64.515 146.660 ;
        RECT 64.595 146.340 64.915 146.660 ;
        RECT 64.995 146.340 65.315 146.660 ;
        RECT 82.305 146.340 82.625 146.660 ;
        RECT 82.705 146.340 83.025 146.660 ;
        RECT 83.105 146.340 83.425 146.660 ;
        RECT 83.505 146.340 83.825 146.660 ;
        RECT 36.030 143.620 36.350 143.940 ;
        RECT 36.430 143.620 36.750 143.940 ;
        RECT 36.830 143.620 37.150 143.940 ;
        RECT 37.230 143.620 37.550 143.940 ;
        RECT 54.540 143.620 54.860 143.940 ;
        RECT 54.940 143.620 55.260 143.940 ;
        RECT 55.340 143.620 55.660 143.940 ;
        RECT 55.740 143.620 56.060 143.940 ;
        RECT 73.050 143.620 73.370 143.940 ;
        RECT 73.450 143.620 73.770 143.940 ;
        RECT 73.850 143.620 74.170 143.940 ;
        RECT 74.250 143.620 74.570 143.940 ;
        RECT 91.560 143.620 91.880 143.940 ;
        RECT 91.960 143.620 92.280 143.940 ;
        RECT 92.360 143.620 92.680 143.940 ;
        RECT 92.760 143.620 93.080 143.940 ;
        RECT 26.775 140.900 27.095 141.220 ;
        RECT 27.175 140.900 27.495 141.220 ;
        RECT 27.575 140.900 27.895 141.220 ;
        RECT 27.975 140.900 28.295 141.220 ;
        RECT 45.285 140.900 45.605 141.220 ;
        RECT 45.685 140.900 46.005 141.220 ;
        RECT 46.085 140.900 46.405 141.220 ;
        RECT 46.485 140.900 46.805 141.220 ;
        RECT 63.795 140.900 64.115 141.220 ;
        RECT 64.195 140.900 64.515 141.220 ;
        RECT 64.595 140.900 64.915 141.220 ;
        RECT 64.995 140.900 65.315 141.220 ;
        RECT 82.305 140.900 82.625 141.220 ;
        RECT 82.705 140.900 83.025 141.220 ;
        RECT 83.105 140.900 83.425 141.220 ;
        RECT 83.505 140.900 83.825 141.220 ;
        RECT 36.030 138.180 36.350 138.500 ;
        RECT 36.430 138.180 36.750 138.500 ;
        RECT 36.830 138.180 37.150 138.500 ;
        RECT 37.230 138.180 37.550 138.500 ;
        RECT 54.540 138.180 54.860 138.500 ;
        RECT 54.940 138.180 55.260 138.500 ;
        RECT 55.340 138.180 55.660 138.500 ;
        RECT 55.740 138.180 56.060 138.500 ;
        RECT 73.050 138.180 73.370 138.500 ;
        RECT 73.450 138.180 73.770 138.500 ;
        RECT 73.850 138.180 74.170 138.500 ;
        RECT 74.250 138.180 74.570 138.500 ;
        RECT 91.560 138.180 91.880 138.500 ;
        RECT 91.960 138.180 92.280 138.500 ;
        RECT 92.360 138.180 92.680 138.500 ;
        RECT 92.760 138.180 93.080 138.500 ;
        RECT 26.775 135.460 27.095 135.780 ;
        RECT 27.175 135.460 27.495 135.780 ;
        RECT 27.575 135.460 27.895 135.780 ;
        RECT 27.975 135.460 28.295 135.780 ;
        RECT 45.285 135.460 45.605 135.780 ;
        RECT 45.685 135.460 46.005 135.780 ;
        RECT 46.085 135.460 46.405 135.780 ;
        RECT 46.485 135.460 46.805 135.780 ;
        RECT 63.795 135.460 64.115 135.780 ;
        RECT 64.195 135.460 64.515 135.780 ;
        RECT 64.595 135.460 64.915 135.780 ;
        RECT 64.995 135.460 65.315 135.780 ;
        RECT 82.305 135.460 82.625 135.780 ;
        RECT 82.705 135.460 83.025 135.780 ;
        RECT 83.105 135.460 83.425 135.780 ;
        RECT 83.505 135.460 83.825 135.780 ;
        RECT 36.030 132.740 36.350 133.060 ;
        RECT 36.430 132.740 36.750 133.060 ;
        RECT 36.830 132.740 37.150 133.060 ;
        RECT 37.230 132.740 37.550 133.060 ;
        RECT 54.540 132.740 54.860 133.060 ;
        RECT 54.940 132.740 55.260 133.060 ;
        RECT 55.340 132.740 55.660 133.060 ;
        RECT 55.740 132.740 56.060 133.060 ;
        RECT 73.050 132.740 73.370 133.060 ;
        RECT 73.450 132.740 73.770 133.060 ;
        RECT 73.850 132.740 74.170 133.060 ;
        RECT 74.250 132.740 74.570 133.060 ;
        RECT 91.560 132.740 91.880 133.060 ;
        RECT 91.960 132.740 92.280 133.060 ;
        RECT 92.360 132.740 92.680 133.060 ;
        RECT 92.760 132.740 93.080 133.060 ;
        RECT 0.940 124.900 2.540 126.500 ;
        RECT 26.550 124.900 28.150 126.500 ;
        RECT 45.280 124.900 46.880 126.500 ;
        RECT 63.800 124.900 65.400 126.500 ;
        RECT 82.250 124.900 83.850 126.500 ;
        RECT 103.005 120.165 103.995 121.155 ;
        RECT 156.565 25.805 157.155 26.395 ;
      LAYER met4 ;
        RECT 3.950 224.760 3.990 225.350 ;
        RECT 88.620 224.760 88.630 225.260 ;
        RECT 121.735 224.760 121.750 225.585 ;
        RECT 132.770 224.760 132.790 225.585 ;
        RECT 140.130 224.760 140.150 225.585 ;
        RECT 147.470 224.760 147.510 225.625 ;
        RECT 155.170 224.760 155.175 225.370 ;
        RECT 3.950 223.615 4.250 224.760 ;
        RECT 7.670 223.615 7.970 224.760 ;
        RECT 11.350 223.615 11.650 224.760 ;
        RECT 15.030 223.615 15.330 224.760 ;
        RECT 18.710 223.615 19.010 224.760 ;
        RECT 22.390 223.615 22.690 224.760 ;
        RECT 26.070 223.615 26.370 224.760 ;
        RECT 29.750 223.615 30.050 224.760 ;
        RECT 33.430 223.615 33.730 224.760 ;
        RECT 37.110 223.615 37.410 224.760 ;
        RECT 40.790 223.615 41.090 224.760 ;
        RECT 44.470 223.615 44.770 224.760 ;
        RECT 48.150 223.615 48.450 224.760 ;
        RECT 51.830 223.615 52.130 224.760 ;
        RECT 55.510 223.615 55.810 224.760 ;
        RECT 59.190 223.615 59.490 224.760 ;
        RECT 62.870 223.615 63.170 224.760 ;
        RECT 66.550 223.615 66.850 224.760 ;
        RECT 70.230 223.615 70.530 224.760 ;
        RECT 73.910 223.615 74.210 224.760 ;
        RECT 77.590 223.615 77.890 224.760 ;
        RECT 81.270 223.615 81.570 224.760 ;
        RECT 84.950 223.615 85.250 224.760 ;
        RECT 88.620 223.615 88.920 224.760 ;
        RECT 3.950 223.315 88.920 223.615 ;
        RECT 17.735 217.725 18.035 223.315 ;
        RECT 55.510 223.300 55.810 223.315 ;
        RECT 62.870 223.270 63.170 223.315 ;
        RECT 114.390 222.705 114.690 224.760 ;
        RECT 114.375 222.375 114.705 222.705 ;
        RECT 118.070 221.720 118.370 224.760 ;
        RECT 118.055 221.390 118.385 221.720 ;
        RECT 121.735 220.760 122.035 224.760 ;
        RECT 121.720 220.430 122.050 220.760 ;
        RECT 125.430 219.680 125.730 224.760 ;
        RECT 125.415 219.350 125.745 219.680 ;
        RECT 129.110 218.515 129.410 224.760 ;
        RECT 129.095 218.185 129.425 218.515 ;
        RECT 8.340 217.425 8.440 217.725 ;
        RECT 9.940 217.425 18.035 217.725 ;
        RECT 132.770 217.275 133.070 224.760 ;
        RECT 132.755 216.945 133.085 217.275 ;
        RECT 136.470 216.035 136.770 224.760 ;
        RECT 136.455 215.705 136.785 216.035 ;
        RECT 140.130 215.075 140.430 224.760 ;
        RECT 140.115 214.745 140.445 215.075 ;
        RECT 143.830 213.955 144.130 224.760 ;
        RECT 143.815 213.625 144.145 213.955 ;
        RECT 147.470 212.985 147.770 224.760 ;
        RECT 147.455 212.655 147.785 212.985 ;
        RECT 151.190 212.010 151.490 224.760 ;
        RECT 151.175 211.680 151.505 212.010 ;
        RECT 154.875 211.035 155.175 224.760 ;
        RECT 154.860 210.705 155.190 211.035 ;
        RECT 26.735 136.700 28.335 206.580 ;
        RECT 26.550 132.660 28.335 136.700 ;
        RECT 35.990 135.350 37.590 206.580 ;
        RECT 35.950 132.660 37.590 135.350 ;
        RECT 45.245 137.090 46.845 206.580 ;
        RECT 45.245 132.660 46.880 137.090 ;
        RECT 54.500 135.550 56.100 206.580 ;
        RECT 63.755 137.470 65.355 206.580 ;
        RECT 54.500 132.660 56.150 135.550 ;
        RECT 63.755 132.660 65.400 137.470 ;
        RECT 73.010 135.850 74.610 206.580 ;
        RECT 82.265 137.750 83.865 206.580 ;
        RECT 26.550 126.505 28.150 132.660 ;
        RECT 0.935 124.895 1.000 126.505 ;
        RECT 2.500 126.500 2.545 126.505 ;
        RECT 2.500 124.900 2.550 126.500 ;
        RECT 2.500 124.895 2.545 124.900 ;
        RECT 26.545 124.895 28.155 126.505 ;
        RECT 35.950 121.450 37.450 132.660 ;
        RECT 45.280 126.505 46.880 132.660 ;
        RECT 45.275 124.895 46.885 126.505 ;
        RECT 54.650 121.450 56.150 132.660 ;
        RECT 63.800 126.505 65.400 132.660 ;
        RECT 72.950 132.660 74.610 135.850 ;
        RECT 82.250 132.660 83.865 137.750 ;
        RECT 91.520 132.660 93.120 206.580 ;
        RECT 63.795 124.895 65.405 126.505 ;
        RECT 72.950 121.450 74.450 132.660 ;
        RECT 82.250 126.505 83.850 132.660 ;
        RECT 82.245 124.895 83.855 126.505 ;
        RECT 9.940 121.160 93.950 121.450 ;
        RECT 9.940 120.160 104.000 121.160 ;
        RECT 9.940 119.950 93.950 120.160 ;
        RECT 156.560 1.000 157.160 26.400 ;
  END
END tt_um_mattvenn_r2r_dac
END LIBRARY

