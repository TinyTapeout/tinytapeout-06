module tt_um_dlmiles_muldiv8_sky130faha (VGND,
    VPWR,
    clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input VGND;
 input VPWR;
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net64;
 wire net65;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _262_;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;
 wire \muldiv.a0_0.GATE ;
 wire \muldiv.a0_0.Q ;
 wire \muldiv.a0_1.Q ;
 wire \muldiv.a0_2.Q ;
 wire \muldiv.a0_3.Q ;
 wire \muldiv.a0_4.Q ;
 wire \muldiv.a0_5.Q ;
 wire \muldiv.a0_6.Q ;
 wire \muldiv.a0_7.Q ;
 wire \muldiv.a1_0.GATE ;
 wire \muldiv.a1_0.Q ;
 wire \muldiv.a1_1.Q ;
 wire \muldiv.a1_2.Q ;
 wire \muldiv.a1_3.Q ;
 wire \muldiv.a1_4.Q ;
 wire \muldiv.a1_5.Q ;
 wire \muldiv.a1_6.Q ;
 wire \muldiv.a1_7.Q ;
 wire \muldiv.div2reg ;
 wire \muldiv.div8.DU_Q0D0d0.fA.A ;
 wire \muldiv.div8.DU_Q0D0d0.fA.B ;
 wire \muldiv.div8.DU_Q0D0d0.fA.CIN ;
 wire \muldiv.div8.DU_Q0D0d0.fA.COUT ;
 wire \muldiv.div8.DU_Q0D0d0.fA.SUM ;
 wire \muldiv.div8.DU_Q0D0d0.io_sel ;
 wire \muldiv.div8.DU_Q0D0d1.fA.A ;
 wire \muldiv.div8.DU_Q0D0d1.fA.B ;
 wire \muldiv.div8.DU_Q0D0d1.fA.COUT ;
 wire \muldiv.div8.DU_Q0D0d1.fA.SUM ;
 wire \muldiv.div8.DU_Q0D0d10_EXT.fA.A ;
 wire \muldiv.div8.DU_Q0D0d10_EXT.fA.CIN ;
 wire \muldiv.div8.DU_Q0D0d10_EXT.fA.COUT ;
 wire \muldiv.div8.DU_Q0D0d10_EXT.fA.SUM ;
 wire \muldiv.div8.DU_Q0D0d11_EXT.fA.A ;
 wire \muldiv.div8.DU_Q0D0d11_EXT.fA.COUT ;
 wire \muldiv.div8.DU_Q0D0d11_EXT.fA.SUM ;
 wire \muldiv.div8.DU_Q0D0d12_EXT.fA.A ;
 wire \muldiv.div8.DU_Q0D0d12_EXT.fA.SUM ;
 wire \muldiv.div8.DU_Q0D0d2.fA.A ;
 wire \muldiv.div8.DU_Q0D0d2.fA.B ;
 wire \muldiv.div8.DU_Q0D0d2.fA.COUT ;
 wire \muldiv.div8.DU_Q0D0d2.fA.SUM ;
 wire \muldiv.div8.DU_Q0D0d3.fA.A ;
 wire \muldiv.div8.DU_Q0D0d3.fA.B ;
 wire \muldiv.div8.DU_Q0D0d3.fA.COUT ;
 wire \muldiv.div8.DU_Q0D0d3.fA.SUM ;
 wire \muldiv.div8.DU_Q0D0d4.fA.A ;
 wire \muldiv.div8.DU_Q0D0d4.fA.B ;
 wire \muldiv.div8.DU_Q0D0d4.fA.COUT ;
 wire \muldiv.div8.DU_Q0D0d4.fA.SUM ;
 wire \muldiv.div8.DU_Q0D0d5.fA.A ;
 wire \muldiv.div8.DU_Q0D0d5.fA.B ;
 wire \muldiv.div8.DU_Q0D0d5.fA.COUT ;
 wire \muldiv.div8.DU_Q0D0d5.fA.SUM ;
 wire \muldiv.div8.DU_Q0D0d6.fA.A ;
 wire \muldiv.div8.DU_Q0D0d6.fA.B ;
 wire \muldiv.div8.DU_Q0D0d6.fA.COUT ;
 wire \muldiv.div8.DU_Q0D0d6.fA.SUM ;
 wire \muldiv.div8.DU_Q0D0d7.fA.A ;
 wire \muldiv.div8.DU_Q0D0d7.fA.B ;
 wire \muldiv.div8.DU_Q0D0d7.fA.COUT ;
 wire \muldiv.div8.DU_Q0D0d7.fA.SUM ;
 wire \muldiv.div8.DU_Q0D0d8_EXT.fA.A ;
 wire \muldiv.div8.DU_Q0D0d8_EXT.fA.COUT ;
 wire \muldiv.div8.DU_Q0D0d8_EXT.fA.SUM ;
 wire \muldiv.div8.DU_Q0D0d9_EXT.fA.A ;
 wire \muldiv.div8.DU_Q0D0d9_EXT.fA.SUM ;
 wire \muldiv.div8.DU_Q1D1d0.fA.A ;
 wire \muldiv.div8.DU_Q1D1d0.fA.COUT ;
 wire \muldiv.div8.DU_Q1D1d0.fA.SUM ;
 wire \muldiv.div8.DU_Q1D1d0.io_sel ;
 wire \muldiv.div8.DU_Q1D1d1.fA.A ;
 wire \muldiv.div8.DU_Q1D1d1.fA.COUT ;
 wire \muldiv.div8.DU_Q1D1d1.fA.SUM ;
 wire \muldiv.div8.DU_Q1D1d10_EXT.fA.A ;
 wire \muldiv.div8.DU_Q1D1d10_EXT.fA.CIN ;
 wire \muldiv.div8.DU_Q1D1d10_EXT.fA.COUT ;
 wire \muldiv.div8.DU_Q1D1d10_EXT.fA.SUM ;
 wire \muldiv.div8.DU_Q1D1d11_EXT.fA.A ;
 wire \muldiv.div8.DU_Q1D1d11_EXT.fA.COUT ;
 wire \muldiv.div8.DU_Q1D1d11_EXT.fA.SUM ;
 wire \muldiv.div8.DU_Q1D1d12_EXT.fA.A ;
 wire \muldiv.div8.DU_Q1D1d12_EXT.fA.SUM ;
 wire \muldiv.div8.DU_Q1D1d2.fA.A ;
 wire \muldiv.div8.DU_Q1D1d2.fA.COUT ;
 wire \muldiv.div8.DU_Q1D1d2.fA.SUM ;
 wire \muldiv.div8.DU_Q1D1d3.fA.A ;
 wire \muldiv.div8.DU_Q1D1d3.fA.COUT ;
 wire \muldiv.div8.DU_Q1D1d3.fA.SUM ;
 wire \muldiv.div8.DU_Q1D1d4.fA.A ;
 wire \muldiv.div8.DU_Q1D1d4.fA.COUT ;
 wire \muldiv.div8.DU_Q1D1d4.fA.SUM ;
 wire \muldiv.div8.DU_Q1D1d5.fA.A ;
 wire \muldiv.div8.DU_Q1D1d5.fA.COUT ;
 wire \muldiv.div8.DU_Q1D1d5.fA.SUM ;
 wire \muldiv.div8.DU_Q1D1d6.fA.A ;
 wire \muldiv.div8.DU_Q1D1d6.fA.COUT ;
 wire \muldiv.div8.DU_Q1D1d6.fA.SUM ;
 wire \muldiv.div8.DU_Q1D1d7.fA.A ;
 wire \muldiv.div8.DU_Q1D1d7.fA.COUT ;
 wire \muldiv.div8.DU_Q1D1d7.fA.SUM ;
 wire \muldiv.div8.DU_Q1D1d8_EXT.fA.A ;
 wire \muldiv.div8.DU_Q1D1d8_EXT.fA.COUT ;
 wire \muldiv.div8.DU_Q1D1d8_EXT.fA.SUM ;
 wire \muldiv.div8.DU_Q1D1d9_EXT.fA.A ;
 wire \muldiv.div8.DU_Q1D1d9_EXT.fA.SUM ;
 wire \muldiv.div8.DU_Q2D2d0.fA.A ;
 wire \muldiv.div8.DU_Q2D2d0.fA.COUT ;
 wire \muldiv.div8.DU_Q2D2d0.fA.SUM ;
 wire \muldiv.div8.DU_Q2D2d0.io_sel ;
 wire \muldiv.div8.DU_Q2D2d1.fA.A ;
 wire \muldiv.div8.DU_Q2D2d1.fA.COUT ;
 wire \muldiv.div8.DU_Q2D2d1.fA.SUM ;
 wire \muldiv.div8.DU_Q2D2d10_EXT.fA.A ;
 wire \muldiv.div8.DU_Q2D2d10_EXT.fA.CIN ;
 wire \muldiv.div8.DU_Q2D2d10_EXT.fA.COUT ;
 wire \muldiv.div8.DU_Q2D2d10_EXT.fA.SUM ;
 wire \muldiv.div8.DU_Q2D2d11_EXT.fA.A ;
 wire \muldiv.div8.DU_Q2D2d11_EXT.fA.SUM ;
 wire \muldiv.div8.DU_Q2D2d2.fA.A ;
 wire \muldiv.div8.DU_Q2D2d2.fA.COUT ;
 wire \muldiv.div8.DU_Q2D2d2.fA.SUM ;
 wire \muldiv.div8.DU_Q2D2d3.fA.A ;
 wire \muldiv.div8.DU_Q2D2d3.fA.COUT ;
 wire \muldiv.div8.DU_Q2D2d3.fA.SUM ;
 wire \muldiv.div8.DU_Q2D2d4.fA.A ;
 wire \muldiv.div8.DU_Q2D2d4.fA.COUT ;
 wire \muldiv.div8.DU_Q2D2d4.fA.SUM ;
 wire \muldiv.div8.DU_Q2D2d5.fA.A ;
 wire \muldiv.div8.DU_Q2D2d5.fA.COUT ;
 wire \muldiv.div8.DU_Q2D2d5.fA.SUM ;
 wire \muldiv.div8.DU_Q2D2d6.fA.A ;
 wire \muldiv.div8.DU_Q2D2d6.fA.COUT ;
 wire \muldiv.div8.DU_Q2D2d6.fA.SUM ;
 wire \muldiv.div8.DU_Q2D2d7.fA.A ;
 wire \muldiv.div8.DU_Q2D2d7.fA.COUT ;
 wire \muldiv.div8.DU_Q2D2d7.fA.SUM ;
 wire \muldiv.div8.DU_Q2D2d8_EXT.fA.A ;
 wire \muldiv.div8.DU_Q2D2d8_EXT.fA.COUT ;
 wire \muldiv.div8.DU_Q2D2d8_EXT.fA.SUM ;
 wire \muldiv.div8.DU_Q2D2d9_EXT.fA.A ;
 wire \muldiv.div8.DU_Q2D2d9_EXT.fA.SUM ;
 wire \muldiv.div8.DU_Q3D3d0.fA.A ;
 wire \muldiv.div8.DU_Q3D3d0.fA.COUT ;
 wire \muldiv.div8.DU_Q3D3d0.fA.SUM ;
 wire \muldiv.div8.DU_Q3D3d0.io_sel ;
 wire \muldiv.div8.DU_Q3D3d1.fA.A ;
 wire \muldiv.div8.DU_Q3D3d1.fA.COUT ;
 wire \muldiv.div8.DU_Q3D3d1.fA.SUM ;
 wire \muldiv.div8.DU_Q3D3d10_EXT.fA.A ;
 wire \muldiv.div8.DU_Q3D3d10_EXT.fA.CIN ;
 wire \muldiv.div8.DU_Q3D3d10_EXT.fA.SUM ;
 wire \muldiv.div8.DU_Q3D3d2.fA.A ;
 wire \muldiv.div8.DU_Q3D3d2.fA.COUT ;
 wire \muldiv.div8.DU_Q3D3d2.fA.SUM ;
 wire \muldiv.div8.DU_Q3D3d3.fA.A ;
 wire \muldiv.div8.DU_Q3D3d3.fA.COUT ;
 wire \muldiv.div8.DU_Q3D3d3.fA.SUM ;
 wire \muldiv.div8.DU_Q3D3d4.fA.A ;
 wire \muldiv.div8.DU_Q3D3d4.fA.COUT ;
 wire \muldiv.div8.DU_Q3D3d4.fA.SUM ;
 wire \muldiv.div8.DU_Q3D3d5.fA.A ;
 wire \muldiv.div8.DU_Q3D3d5.fA.COUT ;
 wire \muldiv.div8.DU_Q3D3d5.fA.SUM ;
 wire \muldiv.div8.DU_Q3D3d6.fA.A ;
 wire \muldiv.div8.DU_Q3D3d6.fA.COUT ;
 wire \muldiv.div8.DU_Q3D3d6.fA.SUM ;
 wire \muldiv.div8.DU_Q3D3d7.fA.A ;
 wire \muldiv.div8.DU_Q3D3d7.fA.COUT ;
 wire \muldiv.div8.DU_Q3D3d7.fA.SUM ;
 wire \muldiv.div8.DU_Q3D3d8_EXT.fA.A ;
 wire \muldiv.div8.DU_Q3D3d8_EXT.fA.COUT ;
 wire \muldiv.div8.DU_Q3D3d8_EXT.fA.SUM ;
 wire \muldiv.div8.DU_Q3D3d9_EXT.fA.A ;
 wire \muldiv.div8.DU_Q3D3d9_EXT.fA.SUM ;
 wire \muldiv.div8.DU_Q4D4d0.fA.A ;
 wire \muldiv.div8.DU_Q4D4d0.fA.COUT ;
 wire \muldiv.div8.DU_Q4D4d0.fA.SUM ;
 wire \muldiv.div8.DU_Q4D4d0.io_sel ;
 wire \muldiv.div8.DU_Q4D4d1.fA.A ;
 wire \muldiv.div8.DU_Q4D4d1.fA.COUT ;
 wire \muldiv.div8.DU_Q4D4d1.fA.SUM ;
 wire \muldiv.div8.DU_Q4D4d2.fA.A ;
 wire \muldiv.div8.DU_Q4D4d2.fA.COUT ;
 wire \muldiv.div8.DU_Q4D4d2.fA.SUM ;
 wire \muldiv.div8.DU_Q4D4d3.fA.A ;
 wire \muldiv.div8.DU_Q4D4d3.fA.COUT ;
 wire \muldiv.div8.DU_Q4D4d3.fA.SUM ;
 wire \muldiv.div8.DU_Q4D4d4.fA.A ;
 wire \muldiv.div8.DU_Q4D4d4.fA.COUT ;
 wire \muldiv.div8.DU_Q4D4d4.fA.SUM ;
 wire \muldiv.div8.DU_Q4D4d5.fA.A ;
 wire \muldiv.div8.DU_Q4D4d5.fA.COUT ;
 wire \muldiv.div8.DU_Q4D4d5.fA.SUM ;
 wire \muldiv.div8.DU_Q4D4d6.fA.A ;
 wire \muldiv.div8.DU_Q4D4d6.fA.COUT ;
 wire \muldiv.div8.DU_Q4D4d6.fA.SUM ;
 wire \muldiv.div8.DU_Q4D4d7.fA.A ;
 wire \muldiv.div8.DU_Q4D4d7.fA.COUT ;
 wire \muldiv.div8.DU_Q4D4d7.fA.SUM ;
 wire \muldiv.div8.DU_Q4D4d8_EXT.fA.A ;
 wire \muldiv.div8.DU_Q4D4d8_EXT.fA.COUT ;
 wire \muldiv.div8.DU_Q4D4d8_EXT.fA.SUM ;
 wire \muldiv.div8.DU_Q4D4d9_EXT.fA.A ;
 wire \muldiv.div8.DU_Q4D4d9_EXT.fA.SUM ;
 wire \muldiv.div8.DU_Q5D5d0.fA.A ;
 wire \muldiv.div8.DU_Q5D5d0.fA.COUT ;
 wire \muldiv.div8.DU_Q5D5d0.fA.SUM ;
 wire \muldiv.div8.DU_Q5D5d0.io_sel ;
 wire \muldiv.div8.DU_Q5D5d1.fA.A ;
 wire \muldiv.div8.DU_Q5D5d1.fA.COUT ;
 wire \muldiv.div8.DU_Q5D5d1.fA.SUM ;
 wire \muldiv.div8.DU_Q5D5d2.fA.A ;
 wire \muldiv.div8.DU_Q5D5d2.fA.COUT ;
 wire \muldiv.div8.DU_Q5D5d2.fA.SUM ;
 wire \muldiv.div8.DU_Q5D5d3.fA.A ;
 wire \muldiv.div8.DU_Q5D5d3.fA.COUT ;
 wire \muldiv.div8.DU_Q5D5d3.fA.SUM ;
 wire \muldiv.div8.DU_Q5D5d4.fA.A ;
 wire \muldiv.div8.DU_Q5D5d4.fA.COUT ;
 wire \muldiv.div8.DU_Q5D5d4.fA.SUM ;
 wire \muldiv.div8.DU_Q5D5d5.fA.A ;
 wire \muldiv.div8.DU_Q5D5d5.fA.COUT ;
 wire \muldiv.div8.DU_Q5D5d5.fA.SUM ;
 wire \muldiv.div8.DU_Q5D5d6.fA.A ;
 wire \muldiv.div8.DU_Q5D5d6.fA.COUT ;
 wire \muldiv.div8.DU_Q5D5d6.fA.SUM ;
 wire \muldiv.div8.DU_Q5D5d7.fA.A ;
 wire \muldiv.div8.DU_Q5D5d7.fA.COUT ;
 wire \muldiv.div8.DU_Q5D5d7.fA.SUM ;
 wire \muldiv.div8.DU_Q5D5d8_EXT.fA.A ;
 wire \muldiv.div8.DU_Q5D5d8_EXT.fA.SUM ;
 wire \muldiv.div8.DU_Q6D6d0.fA.A ;
 wire \muldiv.div8.DU_Q6D6d0.fA.COUT ;
 wire \muldiv.div8.DU_Q6D6d0.fA.SUM ;
 wire \muldiv.div8.DU_Q6D6d0.io_sel ;
 wire \muldiv.div8.DU_Q6D6d1.fA.A ;
 wire \muldiv.div8.DU_Q6D6d1.fA.COUT ;
 wire \muldiv.div8.DU_Q6D6d1.fA.SUM ;
 wire \muldiv.div8.DU_Q6D6d2.fA.A ;
 wire \muldiv.div8.DU_Q6D6d2.fA.COUT ;
 wire \muldiv.div8.DU_Q6D6d2.fA.SUM ;
 wire \muldiv.div8.DU_Q6D6d3.fA.A ;
 wire \muldiv.div8.DU_Q6D6d3.fA.COUT ;
 wire \muldiv.div8.DU_Q6D6d3.fA.SUM ;
 wire \muldiv.div8.DU_Q6D6d4.fA.A ;
 wire \muldiv.div8.DU_Q6D6d4.fA.COUT ;
 wire \muldiv.div8.DU_Q6D6d4.fA.SUM ;
 wire \muldiv.div8.DU_Q6D6d5.fA.A ;
 wire \muldiv.div8.DU_Q6D6d5.fA.COUT ;
 wire \muldiv.div8.DU_Q6D6d5.fA.SUM ;
 wire \muldiv.div8.DU_Q6D6d6.fA.A ;
 wire \muldiv.div8.DU_Q6D6d6.fA.COUT ;
 wire \muldiv.div8.DU_Q6D6d6.fA.SUM ;
 wire \muldiv.div8.DU_Q6D6d7.fA.A ;
 wire \muldiv.div8.DU_Q6D6d7.fA.SUM ;
 wire \muldiv.div8.DU_Q7D7d0.fA.A ;
 wire \muldiv.div8.DU_Q7D7d0.fA.COUT ;
 wire \muldiv.div8.DU_Q7D7d0.fA.SUM ;
 wire \muldiv.div8.DU_Q7D7d0.io_sel ;
 wire \muldiv.div8.DU_Q7D7d1.fA.COUT ;
 wire \muldiv.div8.DU_Q7D7d1.fA.SUM ;
 wire \muldiv.div8.DU_Q7D7d2.fA.COUT ;
 wire \muldiv.div8.DU_Q7D7d2.fA.SUM ;
 wire \muldiv.div8.DU_Q7D7d3.fA.COUT ;
 wire \muldiv.div8.DU_Q7D7d3.fA.SUM ;
 wire \muldiv.div8.DU_Q7D7d4.fA.COUT ;
 wire \muldiv.div8.DU_Q7D7d4.fA.SUM ;
 wire \muldiv.div8.DU_Q7D7d5.fA.COUT ;
 wire \muldiv.div8.DU_Q7D7d5.fA.SUM ;
 wire \muldiv.div8.DU_Q7D7d6.fA.COUT ;
 wire \muldiv.div8.DU_Q7D7d6.fA.SUM ;
 wire \muldiv.div8.DU_Q7D7d7.fA.SUM ;
 wire \muldiv.div8.HAD_DVD_TWOS_0.A ;
 wire \muldiv.div8.HAD_DVD_TWOS_0.B ;
 wire \muldiv.div8.HAD_DVD_TWOS_0.COUT ;
 wire \muldiv.div8.HAD_DVD_TWOS_1.A ;
 wire \muldiv.div8.HAD_DVD_TWOS_1.COUT ;
 wire \muldiv.div8.HAD_DVD_TWOS_2.A ;
 wire \muldiv.div8.HAD_DVD_TWOS_2.COUT ;
 wire \muldiv.div8.HAD_DVD_TWOS_3.A ;
 wire \muldiv.div8.HAD_DVD_TWOS_3.COUT ;
 wire \muldiv.div8.HAD_DVD_TWOS_4.A ;
 wire \muldiv.div8.HAD_DVD_TWOS_4.COUT ;
 wire \muldiv.div8.HAD_DVD_TWOS_5.A ;
 wire \muldiv.div8.HAD_DVD_TWOS_5.COUT ;
 wire \muldiv.div8.HAD_DVD_TWOS_6.A ;
 wire \muldiv.div8.HAD_DVD_TWOS_6.COUT ;
 wire \muldiv.div8.HAD_DVD_TWOS_7.A ;
 wire \muldiv.div8.HAD_DVD_TWOS_7.COUT ;
 wire \muldiv.div8.HAQ0_SIGN.A ;
 wire \muldiv.div8.HAQ0_SIGN.B ;
 wire \muldiv.div8.HAQ0_SIGN.COUT ;
 wire \muldiv.div8.HAQ0_SIGN.SUM ;
 wire \muldiv.div8.HAQ1_SIGN.A ;
 wire \muldiv.div8.HAQ1_SIGN.COUT ;
 wire \muldiv.div8.HAQ1_SIGN.SUM ;
 wire \muldiv.div8.HAQ2_SIGN.A ;
 wire \muldiv.div8.HAQ2_SIGN.COUT ;
 wire \muldiv.div8.HAQ2_SIGN.SUM ;
 wire \muldiv.div8.HAQ3_SIGN.A ;
 wire \muldiv.div8.HAQ3_SIGN.COUT ;
 wire \muldiv.div8.HAQ3_SIGN.SUM ;
 wire \muldiv.div8.HAQ4_SIGN.A ;
 wire \muldiv.div8.HAQ4_SIGN.COUT ;
 wire \muldiv.div8.HAQ4_SIGN.SUM ;
 wire \muldiv.div8.HAQ5_SIGN.A ;
 wire \muldiv.div8.HAQ5_SIGN.COUT ;
 wire \muldiv.div8.HAQ5_SIGN.SUM ;
 wire \muldiv.div8.HAQ6_SIGN.A ;
 wire \muldiv.div8.HAQ6_SIGN.COUT ;
 wire \muldiv.div8.HAQ6_SIGN.SUM ;
 wire \muldiv.div8.HAQ7_SIGN.A ;
 wire \muldiv.div8.HAQ7_SIGN.COUT ;
 wire \muldiv.div8.HAQ7_SIGN.SUM ;
 wire \muldiv.div8.HAR0_SIGN.A ;
 wire \muldiv.div8.HAR0_SIGN.COUT ;
 wire \muldiv.div8.HAR0_SIGN.SUM ;
 wire \muldiv.div8.HAR1_SIGN.A ;
 wire \muldiv.div8.HAR1_SIGN.COUT ;
 wire \muldiv.div8.HAR1_SIGN.SUM ;
 wire \muldiv.div8.HAR2_SIGN.A ;
 wire \muldiv.div8.HAR2_SIGN.COUT ;
 wire \muldiv.div8.HAR2_SIGN.SUM ;
 wire \muldiv.div8.HAR3_SIGN.A ;
 wire \muldiv.div8.HAR3_SIGN.COUT ;
 wire \muldiv.div8.HAR3_SIGN.SUM ;
 wire \muldiv.div8.HAR4_SIGN.A ;
 wire \muldiv.div8.HAR4_SIGN.COUT ;
 wire \muldiv.div8.HAR4_SIGN.SUM ;
 wire \muldiv.div8.HAR5_SIGN.A ;
 wire \muldiv.div8.HAR5_SIGN.COUT ;
 wire \muldiv.div8.HAR5_SIGN.SUM ;
 wire \muldiv.div8.HAR6_SIGN.A ;
 wire \muldiv.div8.HAR6_SIGN.COUT ;
 wire \muldiv.div8.HAR6_SIGN.SUM ;
 wire \muldiv.div8.HAR7_SIGN.A ;
 wire \muldiv.div8.HAR7_SIGN.COUT ;
 wire \muldiv.div8.HAR7_SIGN.SUM ;
 wire \muldiv.div8.io_edivoverflow ;
 wire \muldiv.div8.io_edivzero ;
 wire \muldiv.mul8.A0xB1_8 ;
 wire \muldiv.mul8.A0xB2_16 ;
 wire \muldiv.mul8.A0xB3_24 ;
 wire \muldiv.mul8.A0xB4_32 ;
 wire \muldiv.mul8.A0xB5_40 ;
 wire \muldiv.mul8.A0xB6_48 ;
 wire \muldiv.mul8.A1xB0_1 ;
 wire \muldiv.mul8.A1xB1_9 ;
 wire \muldiv.mul8.A1xB2_17 ;
 wire \muldiv.mul8.A1xB3_25 ;
 wire \muldiv.mul8.A1xB4_33 ;
 wire \muldiv.mul8.A1xB5_41 ;
 wire \muldiv.mul8.A1xB6_49 ;
 wire \muldiv.mul8.A2xB0_2 ;
 wire \muldiv.mul8.A2xB1_10 ;
 wire \muldiv.mul8.A2xB2_18 ;
 wire \muldiv.mul8.A2xB3_26 ;
 wire \muldiv.mul8.A2xB4_34 ;
 wire \muldiv.mul8.A2xB5_42 ;
 wire \muldiv.mul8.A2xB6_50 ;
 wire \muldiv.mul8.A3xB0_3 ;
 wire \muldiv.mul8.A3xB1_11 ;
 wire \muldiv.mul8.A3xB2_19 ;
 wire \muldiv.mul8.A3xB3_27 ;
 wire \muldiv.mul8.A3xB4_35 ;
 wire \muldiv.mul8.A3xB5_43 ;
 wire \muldiv.mul8.A3xB6_51 ;
 wire \muldiv.mul8.A4xB0_4 ;
 wire \muldiv.mul8.A4xB1_12 ;
 wire \muldiv.mul8.A4xB2_20 ;
 wire \muldiv.mul8.A4xB3_28 ;
 wire \muldiv.mul8.A4xB4_36 ;
 wire \muldiv.mul8.A4xB5_44 ;
 wire \muldiv.mul8.A4xB6_52 ;
 wire \muldiv.mul8.A5xB0_5 ;
 wire \muldiv.mul8.A5xB1_13 ;
 wire \muldiv.mul8.A5xB2_21 ;
 wire \muldiv.mul8.A5xB3_29 ;
 wire \muldiv.mul8.A5xB4_37 ;
 wire \muldiv.mul8.A5xB5_45 ;
 wire \muldiv.mul8.A5xB6_53 ;
 wire \muldiv.mul8.A6xB0_6 ;
 wire \muldiv.mul8.A6xB1_14 ;
 wire \muldiv.mul8.A6xB2_22 ;
 wire \muldiv.mul8.A6xB3_30 ;
 wire \muldiv.mul8.A6xB4_38 ;
 wire \muldiv.mul8.A6xB5_46 ;
 wire \muldiv.mul8.A6xB6_54 ;
 wire \muldiv.mul8.A7xB0_7 ;
 wire \muldiv.mul8.A7xB1_15 ;
 wire \muldiv.mul8.A7xB2_23 ;
 wire \muldiv.mul8.A7xB3_31 ;
 wire \muldiv.mul8.A7xB4_39 ;
 wire \muldiv.mul8.A7xB5_47 ;
 wire \muldiv.mul8.A7xB6_55 ;
 wire \muldiv.mul8.FA_P10A3B7.A ;
 wire \muldiv.mul8.FA_P10A3B7.B ;
 wire \muldiv.mul8.FA_P10A3B7.CIN ;
 wire \muldiv.mul8.FA_P10A3B7.COUT ;
 wire \muldiv.mul8.FA_P10A3B7.SUM ;
 wire \muldiv.mul8.FA_P10A4B6.A ;
 wire \muldiv.mul8.FA_P10A4B6.CIN ;
 wire \muldiv.mul8.FA_P10A4B6.COUT ;
 wire \muldiv.mul8.FA_P10A5B5.A ;
 wire \muldiv.mul8.FA_P10A5B5.CIN ;
 wire \muldiv.mul8.FA_P10A5B5.COUT ;
 wire \muldiv.mul8.FA_P10A6B4.A ;
 wire \muldiv.mul8.FA_P10A6B4.CIN ;
 wire \muldiv.mul8.FA_P10A6B4.COUT ;
 wire \muldiv.mul8.FA_P10A7B1.A ;
 wire \muldiv.mul8.FA_P10A7B1.B ;
 wire \muldiv.mul8.FA_P10A7B1.CIN ;
 wire \muldiv.mul8.FA_P10A7B1.COUT ;
 wire \muldiv.mul8.FA_P10A7B1.SUM ;
 wire \muldiv.mul8.FA_P10A7B2.B ;
 wire \muldiv.mul8.FA_P10A7B2.CIN ;
 wire \muldiv.mul8.FA_P10A7B2.COUT ;
 wire \muldiv.mul8.FA_P10A7B2.SUM ;
 wire \muldiv.mul8.FA_P10A7B3.CIN ;
 wire \muldiv.mul8.FA_P10A7B3.COUT ;
 wire \muldiv.mul8.FA_P11A4B7.A ;
 wire \muldiv.mul8.FA_P11A4B7.B ;
 wire \muldiv.mul8.FA_P11A4B7.COUT ;
 wire \muldiv.mul8.FA_P11A4B7.SUM ;
 wire \muldiv.mul8.FA_P11A5B6.A ;
 wire \muldiv.mul8.FA_P11A5B6.COUT ;
 wire \muldiv.mul8.FA_P11A6B5.A ;
 wire \muldiv.mul8.FA_P11A6B5.COUT ;
 wire \muldiv.mul8.FA_P11A7B1.COUT ;
 wire \muldiv.mul8.FA_P11A7B1.SUM ;
 wire \muldiv.mul8.FA_P11A7B2.COUT ;
 wire \muldiv.mul8.FA_P11A7B2.SUM ;
 wire \muldiv.mul8.FA_P11A7B3.B ;
 wire \muldiv.mul8.FA_P11A7B3.COUT ;
 wire \muldiv.mul8.FA_P11A7B3.SUM ;
 wire \muldiv.mul8.FA_P11A7B4.COUT ;
 wire \muldiv.mul8.FA_P12A5B7.A ;
 wire \muldiv.mul8.FA_P12A5B7.B ;
 wire \muldiv.mul8.FA_P12A5B7.COUT ;
 wire \muldiv.mul8.FA_P12A5B7.SUM ;
 wire \muldiv.mul8.FA_P12A6B6.A ;
 wire \muldiv.mul8.FA_P12A6B6.COUT ;
 wire \muldiv.mul8.FA_P12A7B1.COUT ;
 wire \muldiv.mul8.FA_P12A7B1.SUM ;
 wire \muldiv.mul8.FA_P12A7B2.COUT ;
 wire \muldiv.mul8.FA_P12A7B2.SUM ;
 wire \muldiv.mul8.FA_P12A7B3.COUT ;
 wire \muldiv.mul8.FA_P12A7B3.SUM ;
 wire \muldiv.mul8.FA_P12A7B4.B ;
 wire \muldiv.mul8.FA_P12A7B4.COUT ;
 wire \muldiv.mul8.FA_P12A7B4.SUM ;
 wire \muldiv.mul8.FA_P12A7B5.COUT ;
 wire \muldiv.mul8.FA_P13A6B7.A ;
 wire \muldiv.mul8.FA_P13A6B7.B ;
 wire \muldiv.mul8.FA_P13A6B7.COUT ;
 wire \muldiv.mul8.FA_P13A6B7.SUM ;
 wire \muldiv.mul8.FA_P13A7B1.COUT ;
 wire \muldiv.mul8.FA_P13A7B1.SUM ;
 wire \muldiv.mul8.FA_P13A7B2.COUT ;
 wire \muldiv.mul8.FA_P13A7B2.SUM ;
 wire \muldiv.mul8.FA_P13A7B3.COUT ;
 wire \muldiv.mul8.FA_P13A7B3.SUM ;
 wire \muldiv.mul8.FA_P13A7B4.COUT ;
 wire \muldiv.mul8.FA_P13A7B4.SUM ;
 wire \muldiv.mul8.FA_P13A7B5.B ;
 wire \muldiv.mul8.FA_P13A7B5.COUT ;
 wire \muldiv.mul8.FA_P13A7B5.SUM ;
 wire \muldiv.mul8.FA_P13A7B6.COUT ;
 wire \muldiv.mul8.FA_P14A7B1.COUT ;
 wire \muldiv.mul8.FA_P14A7B1.SUM ;
 wire \muldiv.mul8.FA_P14A7B2.COUT ;
 wire \muldiv.mul8.FA_P14A7B2.SUM ;
 wire \muldiv.mul8.FA_P14A7B3.COUT ;
 wire \muldiv.mul8.FA_P14A7B3.SUM ;
 wire \muldiv.mul8.FA_P14A7B4.COUT ;
 wire \muldiv.mul8.FA_P14A7B4.SUM ;
 wire \muldiv.mul8.FA_P14A7B5.COUT ;
 wire \muldiv.mul8.FA_P14A7B5.SUM ;
 wire \muldiv.mul8.FA_P14A7B6.B ;
 wire \muldiv.mul8.FA_P14A7B6.COUT ;
 wire \muldiv.mul8.FA_P14A7B6.SUM ;
 wire \muldiv.mul8.FA_P14A7B7.B ;
 wire \muldiv.mul8.FA_P14A7B7.COUT ;
 wire \muldiv.mul8.FA_P14A7B7.SUM ;
 wire \muldiv.mul8.FA_P15A7B1.COUT ;
 wire \muldiv.mul8.FA_P15A7B1.SUM ;
 wire \muldiv.mul8.FA_P15A7B2.COUT ;
 wire \muldiv.mul8.FA_P15A7B2.SUM ;
 wire \muldiv.mul8.FA_P15A7B3.COUT ;
 wire \muldiv.mul8.FA_P15A7B3.SUM ;
 wire \muldiv.mul8.FA_P15A7B4.COUT ;
 wire \muldiv.mul8.FA_P15A7B4.SUM ;
 wire \muldiv.mul8.FA_P15A7B5.COUT ;
 wire \muldiv.mul8.FA_P15A7B5.SUM ;
 wire \muldiv.mul8.FA_P15A7B6.COUT ;
 wire \muldiv.mul8.FA_P15A7B6.SUM ;
 wire \muldiv.mul8.FA_P15A7B7.B ;
 wire \muldiv.mul8.FA_P15A7B7.COUT ;
 wire \muldiv.mul8.FA_P15A7B7.SUM ;
 wire \muldiv.mul8.FA_P2A1B1.CIN ;
 wire \muldiv.mul8.FA_P2A1B1.COUT ;
 wire \muldiv.mul8.FA_P2A1B1.SUM ;
 wire \muldiv.mul8.FA_P3A1B2.A ;
 wire \muldiv.mul8.FA_P3A1B2.CIN ;
 wire \muldiv.mul8.FA_P3A1B2.COUT ;
 wire \muldiv.mul8.FA_P3A1B2.SUM ;
 wire \muldiv.mul8.FA_P3A2B1.COUT ;
 wire \muldiv.mul8.FA_P4A1B3.A ;
 wire \muldiv.mul8.FA_P4A1B3.CIN ;
 wire \muldiv.mul8.FA_P4A1B3.COUT ;
 wire \muldiv.mul8.FA_P4A1B3.SUM ;
 wire \muldiv.mul8.FA_P4A2B2.A ;
 wire \muldiv.mul8.FA_P4A2B2.COUT ;
 wire \muldiv.mul8.FA_P4A3B1.COUT ;
 wire \muldiv.mul8.FA_P5A1B4.A ;
 wire \muldiv.mul8.FA_P5A1B4.CIN ;
 wire \muldiv.mul8.FA_P5A1B4.COUT ;
 wire \muldiv.mul8.FA_P5A1B4.SUM ;
 wire \muldiv.mul8.FA_P5A2B3.A ;
 wire \muldiv.mul8.FA_P5A2B3.COUT ;
 wire \muldiv.mul8.FA_P5A3B2.A ;
 wire \muldiv.mul8.FA_P5A3B2.COUT ;
 wire \muldiv.mul8.FA_P5A4B1.COUT ;
 wire \muldiv.mul8.FA_P6A1B5.A ;
 wire \muldiv.mul8.FA_P6A1B5.CIN ;
 wire \muldiv.mul8.FA_P6A1B5.COUT ;
 wire \muldiv.mul8.FA_P6A1B5.SUM ;
 wire \muldiv.mul8.FA_P6A2B4.A ;
 wire \muldiv.mul8.FA_P6A2B4.COUT ;
 wire \muldiv.mul8.FA_P6A3B3.A ;
 wire \muldiv.mul8.FA_P6A3B3.COUT ;
 wire \muldiv.mul8.FA_P6A4B2.A ;
 wire \muldiv.mul8.FA_P6A4B2.COUT ;
 wire \muldiv.mul8.FA_P6A5B1.COUT ;
 wire \muldiv.mul8.FA_P7A0B7.A ;
 wire \muldiv.mul8.FA_P7A0B7.B ;
 wire \muldiv.mul8.FA_P7A0B7.COUT ;
 wire \muldiv.mul8.FA_P7A0B7.SUM ;
 wire \muldiv.mul8.FA_P7A1B6.A ;
 wire \muldiv.mul8.FA_P7A1B6.CIN ;
 wire \muldiv.mul8.FA_P7A1B6.COUT ;
 wire \muldiv.mul8.FA_P7A2B5.A ;
 wire \muldiv.mul8.FA_P7A2B5.COUT ;
 wire \muldiv.mul8.FA_P7A3B4.A ;
 wire \muldiv.mul8.FA_P7A3B4.COUT ;
 wire \muldiv.mul8.FA_P7A4B3.A ;
 wire \muldiv.mul8.FA_P7A4B3.COUT ;
 wire \muldiv.mul8.FA_P7A5B2.A ;
 wire \muldiv.mul8.FA_P7A5B2.COUT ;
 wire \muldiv.mul8.FA_P7A6B1.COUT ;
 wire \muldiv.mul8.FA_P8A1B7.A ;
 wire \muldiv.mul8.FA_P8A1B7.B ;
 wire \muldiv.mul8.FA_P8A1B7.COUT ;
 wire \muldiv.mul8.FA_P8A1B7.SUM ;
 wire \muldiv.mul8.FA_P8A2B6.A ;
 wire \muldiv.mul8.FA_P8A2B6.COUT ;
 wire \muldiv.mul8.FA_P8A3B5.A ;
 wire \muldiv.mul8.FA_P8A3B5.COUT ;
 wire \muldiv.mul8.FA_P8A4B4.A ;
 wire \muldiv.mul8.FA_P8A4B4.COUT ;
 wire \muldiv.mul8.FA_P8A5B3.A ;
 wire \muldiv.mul8.FA_P8A5B3.COUT ;
 wire \muldiv.mul8.FA_P8A6B2.A ;
 wire \muldiv.mul8.FA_P8A6B2.COUT ;
 wire \muldiv.mul8.FA_P8A7B1.COUT ;
 wire \muldiv.mul8.FA_P9A2B7.A ;
 wire \muldiv.mul8.FA_P9A2B7.B ;
 wire \muldiv.mul8.FA_P9A2B7.SUM ;
 wire \muldiv.mul8.FA_P9A3B6.A ;
 wire \muldiv.mul8.FA_P9A4B5.A ;
 wire \muldiv.mul8.FA_P9A5B4.A ;
 wire \muldiv.mul8.FA_P9A6B3.A ;
 wire \muldiv.mul8.FA_P9A7B1.SUM ;
 wire \muldiv.mul8.HA_P1A0B1.SUM ;
 wire \muldiv.mul8.HA_P2A0B2.SUM ;
 wire \muldiv.mul8.HA_P3A0B3.SUM ;
 wire \muldiv.mul8.HA_P4A0B4.SUM ;
 wire \muldiv.mul8.HA_P5A0B5.SUM ;
 wire \muldiv.mul8.HA_P6A0B6.SUM ;
 wire \muldiv.negedgeReg_1.area_io_q ;
 wire \muldiv.regR[0] ;
 wire \muldiv.regR[10] ;
 wire \muldiv.regR[11] ;
 wire \muldiv.regR[12] ;
 wire \muldiv.regR[13] ;
 wire \muldiv.regR[14] ;
 wire \muldiv.regR[15] ;
 wire \muldiv.regR[1] ;
 wire \muldiv.regR[2] ;
 wire \muldiv.regR[3] ;
 wire \muldiv.regR[4] ;
 wire \muldiv.regR[5] ;
 wire \muldiv.regR[6] ;
 wire \muldiv.regR[7] ;
 wire \muldiv.regR[8] ;
 wire \muldiv.regR[9] ;
 wire net1;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net2;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net3;
 wire net30;
 wire net31;
 wire net4;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net5;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net6;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;

 sky130_fd_sc_hd__decap_3 FILLER_0_0_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_113 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_125 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_141 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_153 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_165 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_169 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_181 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_193 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_197 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_209 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_221 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_225 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_237 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_249 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_253 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_265 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_277 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_281 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_293 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_305 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_309 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_321 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_0_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_41 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_69 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_85 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_97 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_107 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_10_129 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_10_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_183 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_220 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_232 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_10_264 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_10_291 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_10_299 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_10_315 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_322 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_10_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_10_98 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_11_106 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_11_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_138 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_150 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_162 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_182 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_11_217 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_225 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_11_237 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_244 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_11_256 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_27 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_11_304 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_11_329 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_11_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_11_80 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_90 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_11_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_12_112 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_120 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_147 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_12_158 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_12_171 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_12_179 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_12_187 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_12_220 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_228 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_12_248 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_12_258 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_12_298 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_306 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_309 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_321 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_12_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_12_71 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_13_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_13_121 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_13_160 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_13_211 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_251 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_263 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_27 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_275 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_293 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_305 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_317 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_13_329 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_39 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_13_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_13_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_13_86 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_14_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_115 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_14_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_14_162 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_14_192 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_14_202 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_211 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_14_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_14_239 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_14_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_259 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_14_271 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_14_301 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_309 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_321 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_14_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_14_63 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_88 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_14_92 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_15_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_15_143 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_15_159 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_15_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_173 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_15_186 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_228 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_15_260 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_27 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_308 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_320 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_15_332 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_39 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_16_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_16_131 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_16_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_172 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_16_189 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_16_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_201 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_16_218 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_16_249 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_16_267 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_273 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_29 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_16_304 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_309 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_321 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_41 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_16_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_16_61 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_17_102 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_17_122 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_17_165 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_17_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_173 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_17_188 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_201 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_17_215 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_17_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_231 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_248 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_17_258 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_27 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_299 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_311 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_323 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_39 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_17_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_17_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_63 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_82 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_17_94 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_98 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_18_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_18_129 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_18_161 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_18_191 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_18_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_212 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_18_224 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_232 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_18_246 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_271 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_29 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_294 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_306 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_309 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_321 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_41 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_18_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_18_80 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_85 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_97 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_19_104 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_19_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_135 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_19_160 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_19_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_177 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_19_188 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_19_196 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_19_218 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_19_246 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_19_254 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_27 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_299 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_311 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_323 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_19_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_47 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_19_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_57 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_69 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_19_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_90 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_1_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_113 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_125 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_137 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_149 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_1_161 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_169 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_181 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_193 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_205 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_1_217 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_225 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_237 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_249 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_261 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_1_273 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_281 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_293 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_305 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_317 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_1_329 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_39 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_81 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_93 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_20_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_118 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_20_126 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_132 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_141 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_20_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_157 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_20_165 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_173 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_20_191 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_20_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_201 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_209 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_20_221 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_20_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_257 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_306 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_309 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_321 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_36 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_20_59 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_20_70 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_20_78 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_21_116 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_21_124 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_149 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_21_161 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_169 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_181 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_21_193 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_21_205 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_21_217 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_263 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_21_275 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_21_290 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_21_298 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_21_306 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_316 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_21_328 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_43 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_21_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_21_78 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_22_106 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_22_114 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_144 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_22_156 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_172 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_197 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_22_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_231 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_239 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_22_262 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_277 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_289 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_22_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_22_327 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_22_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_22_58 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_23_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_23_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_121 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_23_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_23_149 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_23_188 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_23_196 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_23_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_229 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_246 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_23_256 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_23_264 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_23_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_23_277 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_281 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_23_293 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_31 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_23_326 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_23_42 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_23_49 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_23_61 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_67 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_76 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_23_88 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_92 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_24_104 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_113 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_24_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_24_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_24_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_24_193 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_197 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_24_209 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_24_224 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_253 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_24_265 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_271 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_280 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_292 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_24_304 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_319 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_24_331 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_24_45 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_24_70 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_24_78 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_24_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_24_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_129 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_25_136 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_25_142 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_150 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_181 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_25_193 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_25_240 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_244 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_25_257 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_267 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_25_275 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_288 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_25_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_25_327 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_25_40 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_44 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_57 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_25_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_93 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_101 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_123 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_144 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_26_156 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_164 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_197 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_209 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_26_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_26_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_26_300 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_26_330 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_45 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_63 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_26_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_27_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_131 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_143 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_27_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_27_164 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_27_191 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_27_203 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_27_222 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_27_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_27_232 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_27_278 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_27_301 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_308 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_27_330 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_27_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_27_47 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_27_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_57 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_74 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_27_80 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_27_91 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_28_101 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_112 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_124 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_28_136 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_28_150 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_28_171 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_183 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_28_214 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_233 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_28_245 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_28_25 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_28_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_28_261 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_288 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_28_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_28_300 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_28_40 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_28_59 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_28_79 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_29_101 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_29_129 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_29_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_29_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_169 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_181 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_29_193 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_207 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_241 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_253 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_265 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_29_277 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_29_306 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_46 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_29_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_74 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_86 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_29_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_109 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_121 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_2_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_141 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_153 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_165 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_177 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_2_189 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_197 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_209 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_221 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_233 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_2_245 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_253 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_265 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_277 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_289 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_2_301 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_309 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_321 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_97 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_30_117 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_30_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_30_160 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_30_189 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_30_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_30_205 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_30_217 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_30_246 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_30_25 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_30_261 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_280 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_30_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_301 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_30_328 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_45 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_30_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_63 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_30_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_102 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_31_113 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_31_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_31_154 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_31_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_173 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_31_201 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_31_219 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_31_233 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_31_256 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_262 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_31_294 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_31_324 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_31_332 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_31_37 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_31_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_76 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_31_94 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_32_115 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_32_127 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_32_141 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_32_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_32_153 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_32_165 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_32_192 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_32_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_32_213 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_219 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_32_249 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_32_285 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_32_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_291 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_32_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_32_325 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_32_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_38 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_32_61 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_32_69 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_32_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_32_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_33_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_33_116 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_124 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_33_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_145 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_33_153 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_33_165 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_33_221 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_33_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_33_23 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_293 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_33_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_33_326 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_33_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_33_43 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_33_50 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_33_74 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_33_86 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_33_98 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_34_115 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_119 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_34_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_34_158 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_34_170 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_176 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_190 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_34_249 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_34_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_34_261 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_265 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_34_296 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_34_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_34_328 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_34_45 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_34_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_34_72 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_34_90 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_35_129 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_35_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_35_176 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_233 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_35_248 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_252 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_35_261 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_265 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_35_295 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_35_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_35_303 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_35_323 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_35_34 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_35_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_35_73 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_94 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_36_114 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_36_126 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_36_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_36_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_231 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_36_24 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_36_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_36_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_36_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_36_300 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_36_329 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_36_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_36_71 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_36_79 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_36_89 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_37_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_37_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_37_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_37_163 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_37_177 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_37_218 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_37_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_244 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_37_295 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_37_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_37_306 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_37_47 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_37_73 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_10 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_38_102 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_106 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_38_118 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_122 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_38_126 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_38_14 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_38_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_145 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_38_162 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_18 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_38_183 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_191 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_38_22 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_231 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_38_239 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_243 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_38_249 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_265 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_38_287 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_38_294 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_298 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_313 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_38_32 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_38_329 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_38_38 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_42 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_38_46 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_50 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_38_6 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_38_62 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_66 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_38_70 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_74 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_38_78 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_38_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_38_92 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_98 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_113 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_125 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_3_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_149 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_3_161 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_198 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_210 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_222 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_252 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_264 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_3_276 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_281 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_293 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_305 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_317 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_3_329 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_93 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_102 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_114 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_126 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_150 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_158 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_4_170 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_174 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_203 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_4_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_4_261 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_282 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_294 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_306 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_309 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_321 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_4_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_91 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_5_102 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_113 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_5_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_5_212 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_220 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_237 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_276 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_299 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_311 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_323 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_5_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_116 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_6_128 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_6_168 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_176 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_209 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_6_221 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_227 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_6_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_6_264 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_268 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_315 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_6_327 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_6_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_73 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_7_103 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_116 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_7_128 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_134 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_7_172 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_7_180 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_186 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_205 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_7_217 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_7_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_229 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_257 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_7_269 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_27 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_275 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_306 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_7_326 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_39 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_7_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_112 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_125 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_8_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_8_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_8_148 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_156 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_8_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_172 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_176 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_8_188 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_8_207 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_211 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_215 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_227 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_239 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_8_249 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_253 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_265 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_306 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_8_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_8_63 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_70 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_88 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_9_106 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_131 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_9_143 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_9_164 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_9_178 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_182 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_9_186 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_9_217 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_9_228 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_9_258 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_9_266 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_27 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_9_272 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_9_286 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_9_330 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_9_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_9_47 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_9_84 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_9_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_49 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_50 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_52 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_56 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_58 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_40 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_59 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_60 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_61 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_62 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_63 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_64 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_66 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_67 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_68 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_70 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_71 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_72 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_73 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_74 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_75 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_76 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_42 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_43 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_44 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_45 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_46 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_47 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_48 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_78 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_79 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_80 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_81 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_82 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_83 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_84 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_85 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_86 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_87 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_88 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_138 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_139 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_140 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_141 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_142 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_143 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_144 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_145 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_146 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_147 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_148 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_149 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_150 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_151 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_152 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_153 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_154 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_155 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_156 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_157 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_158 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_159 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_160 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_161 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_162 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_163 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_164 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_165 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_166 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_167 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_168 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_169 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_170 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_171 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_172 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_173 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_174 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_175 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_176 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_177 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_178 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_179 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_180 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_181 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_182 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_183 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_184 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_185 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_186 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_187 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_188 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_189 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_190 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_191 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_192 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_89 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_90 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_91 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_92 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_93 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_193 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_194 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_195 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_196 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_197 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_198 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_199 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_200 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_201 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_202 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_203 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_204 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_205 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_206 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_207 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_208 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_209 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_210 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_211 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_212 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_213 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_214 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_215 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_216 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_217 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_218 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_219 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_220 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_221 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_222 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_223 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_224 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_225 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_226 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_227 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_228 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_229 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_230 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_231 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_232 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_233 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_234 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_235 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_236 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_237 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_238 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_239 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_240 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_241 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_242 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_243 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_244 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_245 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_246 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_247 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_94 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_95 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_96 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_97 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_98 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_99 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_248 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_249 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_250 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_251 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_252 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_253 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_254 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_255 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_256 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_257 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_258 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_259 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_260 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_261 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_262 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_263 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_264 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_265 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_266 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_267 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_268 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_269 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_270 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_271 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_272 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_273 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_274 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_275 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_276 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_277 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_278 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_279 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_280 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_281 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_282 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_283 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_284 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_285 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_286 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_287 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_288 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_289 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_290 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_291 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_292 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_293 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_294 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_295 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_296 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_297 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_298 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_299 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_300 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_301 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_302 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_100 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_101 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_102 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_103 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_104 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_105 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_106 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_107 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_108 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_109 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_110 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_111 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_112 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_113 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_114 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_115 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_116 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_117 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_118 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_119 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_120 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_121 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_122 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_123 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_124 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_125 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_126 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_127 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_128 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_129 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_130 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_131 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_132 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_133 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_134 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_135 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_136 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_137 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__and2_1 _290_ (.A(_023_),
    .B(\muldiv.a1_2.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_025_));
 sky130_fd_sc_hd__clkbuf_1 _291_ (.A(_025_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.mul8.A0xB2_16 ));
 sky130_fd_sc_hd__and2_1 _292_ (.A(_023_),
    .B(\muldiv.a1_3.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_026_));
 sky130_fd_sc_hd__clkbuf_1 _293_ (.A(_026_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.mul8.A0xB3_24 ));
 sky130_fd_sc_hd__and2_1 _294_ (.A(_023_),
    .B(\muldiv.a1_4.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_027_));
 sky130_fd_sc_hd__clkbuf_1 _295_ (.A(_027_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.mul8.A0xB4_32 ));
 sky130_fd_sc_hd__and2_1 _296_ (.A(_023_),
    .B(\muldiv.a1_5.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_028_));
 sky130_fd_sc_hd__clkbuf_1 _297_ (.A(_028_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.mul8.A0xB5_40 ));
 sky130_fd_sc_hd__and2_1 _298_ (.A(_023_),
    .B(\muldiv.a1_6.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_029_));
 sky130_fd_sc_hd__clkbuf_1 _299_ (.A(_029_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.mul8.A0xB6_48 ));
 sky130_fd_sc_hd__clkbuf_4 _300_ (.A(\muldiv.a1_0.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_030_));
 sky130_fd_sc_hd__and2_1 _301_ (.A(_030_),
    .B(\muldiv.a0_1.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_031_));
 sky130_fd_sc_hd__clkbuf_1 _302_ (.A(_031_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.mul8.A1xB0_1 ));
 sky130_fd_sc_hd__and2_1 _303_ (.A(\muldiv.a1_1.Q ),
    .B(\muldiv.a0_1.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_032_));
 sky130_fd_sc_hd__buf_1 _304_ (.A(_032_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.mul8.A1xB1_9 ));
 sky130_fd_sc_hd__and2_1 _305_ (.A(\muldiv.a1_2.Q ),
    .B(\muldiv.a0_1.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_033_));
 sky130_fd_sc_hd__buf_1 _306_ (.A(_033_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.mul8.A1xB2_17 ));
 sky130_fd_sc_hd__and2_1 _307_ (.A(\muldiv.a1_3.Q ),
    .B(\muldiv.a0_1.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_034_));
 sky130_fd_sc_hd__buf_1 _308_ (.A(_034_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.mul8.A1xB3_25 ));
 sky130_fd_sc_hd__and2_1 _309_ (.A(\muldiv.a1_4.Q ),
    .B(\muldiv.a0_1.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_035_));
 sky130_fd_sc_hd__clkbuf_1 _310_ (.A(_035_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.mul8.A1xB4_33 ));
 sky130_fd_sc_hd__and2_1 _311_ (.A(\muldiv.a1_5.Q ),
    .B(\muldiv.a0_1.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_036_));
 sky130_fd_sc_hd__buf_1 _312_ (.A(_036_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.mul8.A1xB5_41 ));
 sky130_fd_sc_hd__and2_1 _313_ (.A(\muldiv.a1_6.Q ),
    .B(\muldiv.a0_1.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_037_));
 sky130_fd_sc_hd__buf_1 _314_ (.A(_037_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.mul8.A1xB6_49 ));
 sky130_fd_sc_hd__and2_1 _315_ (.A(_030_),
    .B(\muldiv.a0_2.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_038_));
 sky130_fd_sc_hd__buf_1 _316_ (.A(_038_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.mul8.A2xB0_2 ));
 sky130_fd_sc_hd__and2_1 _317_ (.A(\muldiv.a1_1.Q ),
    .B(\muldiv.a0_2.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_039_));
 sky130_fd_sc_hd__buf_1 _318_ (.A(_039_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.mul8.A2xB1_10 ));
 sky130_fd_sc_hd__and2_1 _319_ (.A(\muldiv.a1_2.Q ),
    .B(\muldiv.a0_2.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_040_));
 sky130_fd_sc_hd__buf_1 _320_ (.A(_040_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.mul8.A2xB2_18 ));
 sky130_fd_sc_hd__and2_1 _321_ (.A(\muldiv.a1_3.Q ),
    .B(\muldiv.a0_2.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_041_));
 sky130_fd_sc_hd__clkbuf_1 _322_ (.A(_041_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.mul8.A2xB3_26 ));
 sky130_fd_sc_hd__and2_1 _323_ (.A(\muldiv.a1_4.Q ),
    .B(\muldiv.a0_2.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_042_));
 sky130_fd_sc_hd__buf_1 _324_ (.A(_042_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.mul8.A2xB4_34 ));
 sky130_fd_sc_hd__and2_1 _325_ (.A(\muldiv.a1_5.Q ),
    .B(\muldiv.a0_2.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_043_));
 sky130_fd_sc_hd__buf_1 _326_ (.A(_043_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.mul8.A2xB5_42 ));
 sky130_fd_sc_hd__and2_1 _327_ (.A(\muldiv.a1_6.Q ),
    .B(\muldiv.a0_2.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_044_));
 sky130_fd_sc_hd__clkbuf_1 _328_ (.A(_044_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.mul8.A2xB6_50 ));
 sky130_fd_sc_hd__and2_1 _329_ (.A(_030_),
    .B(\muldiv.a0_3.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_045_));
 sky130_fd_sc_hd__buf_1 _330_ (.A(_045_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.mul8.A3xB0_3 ));
 sky130_fd_sc_hd__and2_1 _331_ (.A(\muldiv.a1_1.Q ),
    .B(\muldiv.a0_3.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_046_));
 sky130_fd_sc_hd__buf_1 _332_ (.A(_046_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.mul8.A3xB1_11 ));
 sky130_fd_sc_hd__and2_1 _333_ (.A(\muldiv.a1_2.Q ),
    .B(\muldiv.a0_3.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_047_));
 sky130_fd_sc_hd__buf_1 _334_ (.A(_047_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.mul8.A3xB2_19 ));
 sky130_fd_sc_hd__and2_1 _335_ (.A(\muldiv.a1_3.Q ),
    .B(\muldiv.a0_3.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_048_));
 sky130_fd_sc_hd__buf_1 _336_ (.A(_048_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.mul8.A3xB3_27 ));
 sky130_fd_sc_hd__and2_1 _337_ (.A(\muldiv.a1_4.Q ),
    .B(\muldiv.a0_3.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_049_));
 sky130_fd_sc_hd__buf_1 _338_ (.A(_049_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.mul8.A3xB4_35 ));
 sky130_fd_sc_hd__and2_1 _339_ (.A(\muldiv.a1_5.Q ),
    .B(\muldiv.a0_3.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_050_));
 sky130_fd_sc_hd__buf_1 _340_ (.A(_050_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.mul8.A3xB5_43 ));
 sky130_fd_sc_hd__and2_1 _341_ (.A(\muldiv.a1_6.Q ),
    .B(\muldiv.a0_3.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_051_));
 sky130_fd_sc_hd__buf_1 _342_ (.A(_051_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.mul8.A3xB6_51 ));
 sky130_fd_sc_hd__and2_1 _343_ (.A(_030_),
    .B(\muldiv.a0_4.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_052_));
 sky130_fd_sc_hd__buf_1 _344_ (.A(_052_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.mul8.A4xB0_4 ));
 sky130_fd_sc_hd__and2_1 _345_ (.A(\muldiv.a1_1.Q ),
    .B(\muldiv.a0_4.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_053_));
 sky130_fd_sc_hd__buf_1 _346_ (.A(_053_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.mul8.A4xB1_12 ));
 sky130_fd_sc_hd__and2_1 _347_ (.A(\muldiv.a1_2.Q ),
    .B(\muldiv.a0_4.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_054_));
 sky130_fd_sc_hd__buf_1 _348_ (.A(_054_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.mul8.A4xB2_20 ));
 sky130_fd_sc_hd__and2_1 _349_ (.A(\muldiv.a1_3.Q ),
    .B(\muldiv.a0_4.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_055_));
 sky130_fd_sc_hd__clkbuf_1 _350_ (.A(_055_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.mul8.A4xB3_28 ));
 sky130_fd_sc_hd__and2_1 _351_ (.A(\muldiv.a1_4.Q ),
    .B(\muldiv.a0_4.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_056_));
 sky130_fd_sc_hd__buf_1 _352_ (.A(_056_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.mul8.A4xB4_36 ));
 sky130_fd_sc_hd__and2_1 _353_ (.A(\muldiv.a1_5.Q ),
    .B(\muldiv.a0_4.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_057_));
 sky130_fd_sc_hd__buf_1 _354_ (.A(_057_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.mul8.A4xB5_44 ));
 sky130_fd_sc_hd__and2_1 _355_ (.A(\muldiv.a1_6.Q ),
    .B(\muldiv.a0_4.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_058_));
 sky130_fd_sc_hd__buf_1 _356_ (.A(_058_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.mul8.A4xB6_52 ));
 sky130_fd_sc_hd__and2_1 _357_ (.A(_030_),
    .B(\muldiv.a0_5.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_059_));
 sky130_fd_sc_hd__buf_1 _358_ (.A(_059_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.mul8.A5xB0_5 ));
 sky130_fd_sc_hd__and2_1 _359_ (.A(\muldiv.a1_1.Q ),
    .B(\muldiv.a0_5.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_060_));
 sky130_fd_sc_hd__buf_1 _360_ (.A(_060_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.mul8.A5xB1_13 ));
 sky130_fd_sc_hd__and2_1 _361_ (.A(\muldiv.a1_2.Q ),
    .B(\muldiv.a0_5.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_061_));
 sky130_fd_sc_hd__buf_1 _362_ (.A(_061_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.mul8.A5xB2_21 ));
 sky130_fd_sc_hd__and2_1 _363_ (.A(\muldiv.a1_3.Q ),
    .B(\muldiv.a0_5.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_062_));
 sky130_fd_sc_hd__buf_1 _364_ (.A(_062_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.mul8.A5xB3_29 ));
 sky130_fd_sc_hd__and2_1 _365_ (.A(\muldiv.a1_4.Q ),
    .B(\muldiv.a0_5.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_063_));
 sky130_fd_sc_hd__buf_1 _366_ (.A(_063_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.mul8.A5xB4_37 ));
 sky130_fd_sc_hd__and2_1 _367_ (.A(\muldiv.a1_5.Q ),
    .B(\muldiv.a0_5.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_064_));
 sky130_fd_sc_hd__buf_1 _368_ (.A(_064_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.mul8.A5xB5_45 ));
 sky130_fd_sc_hd__and2_1 _369_ (.A(\muldiv.a1_6.Q ),
    .B(\muldiv.a0_5.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_065_));
 sky130_fd_sc_hd__clkbuf_1 _370_ (.A(_065_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.mul8.A5xB6_53 ));
 sky130_fd_sc_hd__and2_1 _371_ (.A(_030_),
    .B(\muldiv.a0_6.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_066_));
 sky130_fd_sc_hd__buf_1 _372_ (.A(_066_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.mul8.A6xB0_6 ));
 sky130_fd_sc_hd__and2_1 _373_ (.A(\muldiv.a1_1.Q ),
    .B(\muldiv.a0_6.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_067_));
 sky130_fd_sc_hd__buf_1 _374_ (.A(_067_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.mul8.A6xB1_14 ));
 sky130_fd_sc_hd__and2_1 _375_ (.A(\muldiv.a1_2.Q ),
    .B(\muldiv.a0_6.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_068_));
 sky130_fd_sc_hd__buf_1 _376_ (.A(_068_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.mul8.A6xB2_22 ));
 sky130_fd_sc_hd__and2_1 _377_ (.A(\muldiv.a1_3.Q ),
    .B(\muldiv.a0_6.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_069_));
 sky130_fd_sc_hd__clkbuf_1 _378_ (.A(_069_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.mul8.A6xB3_30 ));
 sky130_fd_sc_hd__and2_1 _379_ (.A(\muldiv.a1_4.Q ),
    .B(\muldiv.a0_6.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_070_));
 sky130_fd_sc_hd__buf_1 _380_ (.A(_070_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.mul8.A6xB4_38 ));
 sky130_fd_sc_hd__and2_1 _381_ (.A(\muldiv.a1_5.Q ),
    .B(\muldiv.a0_6.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_071_));
 sky130_fd_sc_hd__clkbuf_1 _382_ (.A(_071_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.mul8.A6xB5_46 ));
 sky130_fd_sc_hd__and2_1 _383_ (.A(\muldiv.a1_6.Q ),
    .B(\muldiv.a0_6.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_072_));
 sky130_fd_sc_hd__clkbuf_1 _384_ (.A(_072_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.mul8.A6xB6_54 ));
 sky130_fd_sc_hd__clkbuf_2 _385_ (.A(_020_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_073_));
 sky130_fd_sc_hd__and2_1 _386_ (.A(_073_),
    .B(_030_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_074_));
 sky130_fd_sc_hd__buf_1 _387_ (.A(_074_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.mul8.A7xB0_7 ));
 sky130_fd_sc_hd__and2_1 _388_ (.A(_073_),
    .B(\muldiv.a1_1.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_075_));
 sky130_fd_sc_hd__clkbuf_1 _389_ (.A(_075_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.mul8.A7xB1_15 ));
 sky130_fd_sc_hd__and2_1 _390_ (.A(_073_),
    .B(\muldiv.a1_2.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_076_));
 sky130_fd_sc_hd__buf_1 _391_ (.A(_076_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.mul8.A7xB2_23 ));
 sky130_fd_sc_hd__and2_1 _392_ (.A(_073_),
    .B(\muldiv.a1_3.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_077_));
 sky130_fd_sc_hd__buf_1 _393_ (.A(_077_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.mul8.A7xB3_31 ));
 sky130_fd_sc_hd__and2_1 _394_ (.A(_073_),
    .B(\muldiv.a1_4.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_078_));
 sky130_fd_sc_hd__buf_1 _395_ (.A(_078_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.mul8.A7xB4_39 ));
 sky130_fd_sc_hd__and2_1 _396_ (.A(_073_),
    .B(\muldiv.a1_5.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_079_));
 sky130_fd_sc_hd__buf_1 _397_ (.A(_079_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.mul8.A7xB5_47 ));
 sky130_fd_sc_hd__and2_1 _398_ (.A(_073_),
    .B(\muldiv.a1_6.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_080_));
 sky130_fd_sc_hd__buf_1 _399_ (.A(_080_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.mul8.A7xB6_55 ));
 sky130_fd_sc_hd__buf_2 _400_ (.A(net12),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_081_));
 sky130_fd_sc_hd__and3_1 _401_ (.A(_081_),
    .B(_073_),
    .C(_030_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_082_));
 sky130_fd_sc_hd__buf_4 _402_ (.A(_082_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.mul8.FA_P10A7B1.A ));
 sky130_fd_sc_hd__and3_1 _403_ (.A(_081_),
    .B(_020_),
    .C(\muldiv.a1_1.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_083_));
 sky130_fd_sc_hd__clkbuf_4 _404_ (.A(_083_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.mul8.FA_P10A7B1.B ));
 sky130_fd_sc_hd__and3_1 _405_ (.A(_081_),
    .B(_020_),
    .C(\muldiv.a1_2.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_084_));
 sky130_fd_sc_hd__clkbuf_4 _406_ (.A(_084_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.mul8.FA_P10A7B2.B ));
 sky130_fd_sc_hd__and3_1 _407_ (.A(_081_),
    .B(_020_),
    .C(\muldiv.a1_3.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_085_));
 sky130_fd_sc_hd__clkbuf_4 _408_ (.A(_085_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.mul8.FA_P11A7B3.B ));
 sky130_fd_sc_hd__and3_1 _409_ (.A(_081_),
    .B(_020_),
    .C(\muldiv.a1_4.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_086_));
 sky130_fd_sc_hd__buf_2 _410_ (.A(_086_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.mul8.FA_P12A7B4.B ));
 sky130_fd_sc_hd__and3_1 _411_ (.A(_081_),
    .B(_020_),
    .C(\muldiv.a1_5.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_087_));
 sky130_fd_sc_hd__clkbuf_2 _412_ (.A(_087_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.mul8.FA_P13A7B5.B ));
 sky130_fd_sc_hd__and3_1 _413_ (.A(_081_),
    .B(_020_),
    .C(\muldiv.a1_6.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_088_));
 sky130_fd_sc_hd__buf_1 _414_ (.A(_088_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.mul8.FA_P14A7B6.B ));
 sky130_fd_sc_hd__or2_1 _415_ (.A(_081_),
    .B(_020_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_089_));
 sky130_fd_sc_hd__and3_1 _416_ (.A(\muldiv.a1_7.Q ),
    .B(_021_),
    .C(_089_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_090_));
 sky130_fd_sc_hd__buf_1 _417_ (.A(_090_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.mul8.FA_P14A7B7.B ));
 sky130_fd_sc_hd__buf_8 _418_ (.A(_022_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_091_));
 sky130_fd_sc_hd__nor2_1 _419_ (.A(_073_),
    .B(net75),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\muldiv.mul8.FA_P15A7B7.B ));
 sky130_fd_sc_hd__and2b_1 _420_ (.A_N(\muldiv.negedgeReg_1.area_io_q ),
    .B(\muldiv.div2reg ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_092_));
 sky130_fd_sc_hd__clkbuf_2 _421_ (.A(_092_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.a1_0.GATE ));
 sky130_fd_sc_hd__and2b_1 _422_ (.A_N(\muldiv.div2reg ),
    .B(\muldiv.negedgeReg_1.area_io_q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_093_));
 sky130_fd_sc_hd__clkbuf_2 _423_ (.A(_093_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.a0_0.GATE ));
 sky130_fd_sc_hd__mux2_4 _424_ (.A0(\muldiv.div8.DU_Q1D1d0.fA.A ),
    .A1(\muldiv.div8.DU_Q1D1d0.fA.SUM ),
    .S(\muldiv.div8.DU_Q1D1d0.io_sel ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_094_));
 sky130_fd_sc_hd__buf_6 _425_ (.A(_094_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.div8.DU_Q0D0d1.fA.A ));
 sky130_fd_sc_hd__mux2_4 _426_ (.A0(\muldiv.div8.DU_Q2D2d0.fA.A ),
    .A1(\muldiv.div8.DU_Q2D2d0.fA.SUM ),
    .S(\muldiv.div8.DU_Q2D2d0.io_sel ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_095_));
 sky130_fd_sc_hd__buf_6 _427_ (.A(_095_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.div8.DU_Q1D1d1.fA.A ));
 sky130_fd_sc_hd__inv_2 _428_ (.A(\muldiv.div8.DU_Q1D1d0.io_sel ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_096_));
 sky130_fd_sc_hd__buf_4 _429_ (.A(_096_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_097_));
 sky130_fd_sc_hd__mux2_1 _430_ (.A0(\muldiv.div8.DU_Q1D1d1.fA.SUM ),
    .A1(\muldiv.div8.DU_Q1D1d1.fA.A ),
    .S(_097_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_098_));
 sky130_fd_sc_hd__buf_1 _431_ (.A(_098_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.div8.DU_Q0D0d2.fA.A ));
 sky130_fd_sc_hd__mux2_4 _432_ (.A0(\muldiv.div8.DU_Q3D3d0.fA.A ),
    .A1(\muldiv.div8.DU_Q3D3d0.fA.SUM ),
    .S(\muldiv.div8.DU_Q3D3d0.io_sel ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_099_));
 sky130_fd_sc_hd__buf_6 _433_ (.A(_099_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.div8.DU_Q2D2d1.fA.A ));
 sky130_fd_sc_hd__inv_2 _434_ (.A(\muldiv.div8.DU_Q2D2d0.io_sel ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_100_));
 sky130_fd_sc_hd__clkbuf_4 _435_ (.A(_100_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_101_));
 sky130_fd_sc_hd__mux2_1 _436_ (.A0(\muldiv.div8.DU_Q2D2d1.fA.SUM ),
    .A1(\muldiv.div8.DU_Q2D2d1.fA.A ),
    .S(_101_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_102_));
 sky130_fd_sc_hd__buf_1 _437_ (.A(_102_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.div8.DU_Q1D1d2.fA.A ));
 sky130_fd_sc_hd__mux2_1 _438_ (.A0(\muldiv.div8.DU_Q1D1d2.fA.SUM ),
    .A1(\muldiv.div8.DU_Q1D1d2.fA.A ),
    .S(_097_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_103_));
 sky130_fd_sc_hd__buf_1 _439_ (.A(_103_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.div8.DU_Q0D0d3.fA.A ));
 sky130_fd_sc_hd__mux2_4 _440_ (.A0(\muldiv.div8.DU_Q4D4d0.fA.A ),
    .A1(\muldiv.div8.DU_Q4D4d0.fA.SUM ),
    .S(\muldiv.div8.DU_Q4D4d0.io_sel ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_104_));
 sky130_fd_sc_hd__buf_6 _441_ (.A(_104_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.div8.DU_Q3D3d1.fA.A ));
 sky130_fd_sc_hd__inv_2 _442_ (.A(\muldiv.div8.DU_Q3D3d0.io_sel ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_105_));
 sky130_fd_sc_hd__mux2_1 _443_ (.A0(\muldiv.div8.DU_Q3D3d1.fA.SUM ),
    .A1(\muldiv.div8.DU_Q3D3d1.fA.A ),
    .S(_105_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_106_));
 sky130_fd_sc_hd__buf_1 _444_ (.A(_106_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.div8.DU_Q2D2d2.fA.A ));
 sky130_fd_sc_hd__mux2_1 _445_ (.A0(\muldiv.div8.DU_Q2D2d2.fA.SUM ),
    .A1(\muldiv.div8.DU_Q2D2d2.fA.A ),
    .S(_100_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_107_));
 sky130_fd_sc_hd__buf_1 _446_ (.A(_107_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.div8.DU_Q1D1d3.fA.A ));
 sky130_fd_sc_hd__mux2_1 _447_ (.A0(\muldiv.div8.DU_Q1D1d3.fA.SUM ),
    .A1(\muldiv.div8.DU_Q1D1d3.fA.A ),
    .S(_097_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_108_));
 sky130_fd_sc_hd__buf_1 _448_ (.A(_108_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.div8.DU_Q0D0d4.fA.A ));
 sky130_fd_sc_hd__mux2_4 _449_ (.A0(\muldiv.div8.DU_Q5D5d0.fA.A ),
    .A1(\muldiv.div8.DU_Q5D5d0.fA.SUM ),
    .S(\muldiv.div8.DU_Q5D5d0.io_sel ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_109_));
 sky130_fd_sc_hd__buf_6 _450_ (.A(_109_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.div8.DU_Q4D4d1.fA.A ));
 sky130_fd_sc_hd__inv_2 _451_ (.A(\muldiv.div8.DU_Q4D4d0.io_sel ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_110_));
 sky130_fd_sc_hd__and2_1 _452_ (.A(\muldiv.div8.DU_Q4D4d0.io_sel ),
    .B(\muldiv.div8.DU_Q4D4d1.fA.SUM ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_111_));
 sky130_fd_sc_hd__a21o_1 _453_ (.A1(_110_),
    .A2(\muldiv.div8.DU_Q4D4d1.fA.A ),
    .B1(_111_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.div8.DU_Q3D3d2.fA.A ));
 sky130_fd_sc_hd__a211o_1 _454_ (.A1(_110_),
    .A2(\muldiv.div8.DU_Q4D4d1.fA.A ),
    .B1(_111_),
    .C1(\muldiv.div8.DU_Q3D3d0.io_sel ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_112_));
 sky130_fd_sc_hd__clkbuf_4 _455_ (.A(_105_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_113_));
 sky130_fd_sc_hd__or2_1 _456_ (.A(_113_),
    .B(\muldiv.div8.DU_Q3D3d2.fA.SUM ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_114_));
 sky130_fd_sc_hd__and2_1 _457_ (.A(_112_),
    .B(_114_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_115_));
 sky130_fd_sc_hd__buf_1 _458_ (.A(_115_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.div8.DU_Q2D2d3.fA.A ));
 sky130_fd_sc_hd__and2_1 _459_ (.A(\muldiv.div8.DU_Q2D2d0.io_sel ),
    .B(\muldiv.div8.DU_Q2D2d3.fA.SUM ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_116_));
 sky130_fd_sc_hd__a31o_1 _460_ (.A1(_101_),
    .A2(_112_),
    .A3(_114_),
    .B1(_116_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.div8.DU_Q1D1d4.fA.A ));
 sky130_fd_sc_hd__mux2_1 _461_ (.A0(\muldiv.div8.DU_Q1D1d4.fA.SUM ),
    .A1(\muldiv.div8.DU_Q1D1d4.fA.A ),
    .S(_096_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_117_));
 sky130_fd_sc_hd__buf_1 _462_ (.A(_117_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.div8.DU_Q0D0d5.fA.A ));
 sky130_fd_sc_hd__buf_6 _463_ (.A(\muldiv.div8.DU_Q6D6d0.io_sel ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_118_));
 sky130_fd_sc_hd__mux2_4 _464_ (.A0(\muldiv.div8.DU_Q6D6d0.fA.A ),
    .A1(\muldiv.div8.DU_Q6D6d0.fA.SUM ),
    .S(_118_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_119_));
 sky130_fd_sc_hd__buf_6 _465_ (.A(_119_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.div8.DU_Q5D5d1.fA.A ));
 sky130_fd_sc_hd__inv_2 _466_ (.A(net69),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_120_));
 sky130_fd_sc_hd__and2_1 _467_ (.A(\muldiv.div8.DU_Q5D5d0.io_sel ),
    .B(\muldiv.div8.DU_Q5D5d1.fA.SUM ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_121_));
 sky130_fd_sc_hd__a21o_1 _468_ (.A1(_120_),
    .A2(\muldiv.div8.DU_Q5D5d1.fA.A ),
    .B1(_121_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.div8.DU_Q4D4d2.fA.A ));
 sky130_fd_sc_hd__a211o_1 _469_ (.A1(_120_),
    .A2(\muldiv.div8.DU_Q5D5d1.fA.A ),
    .B1(_121_),
    .C1(\muldiv.div8.DU_Q4D4d0.io_sel ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_122_));
 sky130_fd_sc_hd__or2_1 _470_ (.A(_110_),
    .B(\muldiv.div8.DU_Q4D4d2.fA.SUM ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_123_));
 sky130_fd_sc_hd__and2_1 _471_ (.A(_122_),
    .B(_123_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_124_));
 sky130_fd_sc_hd__buf_1 _472_ (.A(_124_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.div8.DU_Q3D3d3.fA.A ));
 sky130_fd_sc_hd__and2_1 _473_ (.A(\muldiv.div8.DU_Q3D3d0.io_sel ),
    .B(\muldiv.div8.DU_Q3D3d3.fA.SUM ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_125_));
 sky130_fd_sc_hd__a31o_1 _474_ (.A1(_113_),
    .A2(_122_),
    .A3(_123_),
    .B1(_125_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.div8.DU_Q2D2d4.fA.A ));
 sky130_fd_sc_hd__a311o_1 _475_ (.A1(_113_),
    .A2(_122_),
    .A3(_123_),
    .B1(_125_),
    .C1(\muldiv.div8.DU_Q2D2d0.io_sel ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_126_));
 sky130_fd_sc_hd__or2_1 _476_ (.A(_101_),
    .B(\muldiv.div8.DU_Q2D2d4.fA.SUM ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_127_));
 sky130_fd_sc_hd__and2_1 _477_ (.A(_126_),
    .B(_127_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_128_));
 sky130_fd_sc_hd__buf_1 _478_ (.A(_128_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.div8.DU_Q1D1d5.fA.A ));
 sky130_fd_sc_hd__and2_1 _479_ (.A(\muldiv.div8.DU_Q1D1d0.io_sel ),
    .B(\muldiv.div8.DU_Q1D1d5.fA.SUM ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_129_));
 sky130_fd_sc_hd__a31o_1 _480_ (.A1(_097_),
    .A2(_126_),
    .A3(_127_),
    .B1(_129_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.div8.DU_Q0D0d6.fA.A ));
 sky130_fd_sc_hd__buf_6 _481_ (.A(\muldiv.div8.DU_Q7D7d0.io_sel ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_130_));
 sky130_fd_sc_hd__mux2_4 _482_ (.A0(\muldiv.div8.DU_Q7D7d0.fA.A ),
    .A1(\muldiv.div8.DU_Q7D7d0.fA.SUM ),
    .S(_130_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_131_));
 sky130_fd_sc_hd__buf_6 _483_ (.A(_131_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.div8.DU_Q6D6d1.fA.A ));
 sky130_fd_sc_hd__or2b_1 _484_ (.A(\muldiv.div8.DU_Q6D6d1.fA.SUM ),
    .B_N(net76),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_132_));
 sky130_fd_sc_hd__o21a_1 _485_ (.A1(_118_),
    .A2(\muldiv.div8.DU_Q6D6d1.fA.A ),
    .B1(_132_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.div8.DU_Q5D5d2.fA.A ));
 sky130_fd_sc_hd__and2_1 _486_ (.A(\muldiv.div8.DU_Q5D5d0.io_sel ),
    .B(\muldiv.div8.DU_Q5D5d2.fA.SUM ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_133_));
 sky130_fd_sc_hd__o211a_1 _487_ (.A1(net76),
    .A2(\muldiv.div8.DU_Q6D6d1.fA.A ),
    .B1(_132_),
    .C1(_120_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_134_));
 sky130_fd_sc_hd__or2_1 _488_ (.A(_133_),
    .B(_134_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_135_));
 sky130_fd_sc_hd__buf_1 _489_ (.A(_135_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.div8.DU_Q4D4d3.fA.A ));
 sky130_fd_sc_hd__or2_1 _490_ (.A(_110_),
    .B(\muldiv.div8.DU_Q4D4d3.fA.SUM ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_136_));
 sky130_fd_sc_hd__o21a_1 _491_ (.A1(\muldiv.div8.DU_Q4D4d0.io_sel ),
    .A2(\muldiv.div8.DU_Q4D4d3.fA.A ),
    .B1(_136_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.div8.DU_Q3D3d4.fA.A ));
 sky130_fd_sc_hd__and2_1 _492_ (.A(\muldiv.div8.DU_Q3D3d0.io_sel ),
    .B(\muldiv.div8.DU_Q3D3d4.fA.SUM ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_137_));
 sky130_fd_sc_hd__o311a_1 _493_ (.A1(\muldiv.div8.DU_Q4D4d0.io_sel ),
    .A2(_133_),
    .A3(_134_),
    .B1(_136_),
    .C1(_113_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_138_));
 sky130_fd_sc_hd__or2_1 _494_ (.A(_137_),
    .B(_138_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_139_));
 sky130_fd_sc_hd__buf_1 _495_ (.A(_139_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.div8.DU_Q2D2d5.fA.A ));
 sky130_fd_sc_hd__or2_1 _496_ (.A(_101_),
    .B(\muldiv.div8.DU_Q2D2d5.fA.SUM ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_140_));
 sky130_fd_sc_hd__o21a_1 _497_ (.A1(\muldiv.div8.DU_Q2D2d0.io_sel ),
    .A2(\muldiv.div8.DU_Q2D2d5.fA.A ),
    .B1(_140_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.div8.DU_Q1D1d6.fA.A ));
 sky130_fd_sc_hd__and2_1 _498_ (.A(\muldiv.div8.DU_Q1D1d0.io_sel ),
    .B(\muldiv.div8.DU_Q1D1d6.fA.SUM ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_141_));
 sky130_fd_sc_hd__o311a_1 _499_ (.A1(\muldiv.div8.DU_Q2D2d0.io_sel ),
    .A2(_137_),
    .A3(_138_),
    .B1(_140_),
    .C1(_097_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_142_));
 sky130_fd_sc_hd__or2_1 _500_ (.A(_141_),
    .B(_142_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_143_));
 sky130_fd_sc_hd__buf_1 _501_ (.A(_143_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.div8.DU_Q0D0d7.fA.A ));
 sky130_fd_sc_hd__and2_1 _502_ (.A(_130_),
    .B(\muldiv.div8.DU_Q7D7d2.fA.SUM ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_144_));
 sky130_fd_sc_hd__buf_1 _503_ (.A(_144_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.div8.DU_Q6D6d3.fA.A ));
 sky130_fd_sc_hd__a21o_1 _504_ (.A1(net77),
    .A2(\muldiv.div8.DU_Q7D7d2.fA.SUM ),
    .B1(_118_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_145_));
 sky130_fd_sc_hd__or2b_1 _505_ (.A(\muldiv.div8.DU_Q6D6d3.fA.SUM ),
    .B_N(net73),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_146_));
 sky130_fd_sc_hd__and2_1 _506_ (.A(_145_),
    .B(_146_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_147_));
 sky130_fd_sc_hd__buf_1 _507_ (.A(_147_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.div8.DU_Q5D5d4.fA.A ));
 sky130_fd_sc_hd__and2_1 _508_ (.A(\muldiv.div8.DU_Q5D5d0.io_sel ),
    .B(\muldiv.div8.DU_Q5D5d4.fA.SUM ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_148_));
 sky130_fd_sc_hd__a31o_1 _509_ (.A1(_120_),
    .A2(_145_),
    .A3(_146_),
    .B1(_148_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.div8.DU_Q4D4d5.fA.A ));
 sky130_fd_sc_hd__mux2_1 _510_ (.A0(\muldiv.div8.DU_Q4D4d5.fA.SUM ),
    .A1(\muldiv.div8.DU_Q4D4d5.fA.A ),
    .S(_110_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_149_));
 sky130_fd_sc_hd__buf_1 _511_ (.A(_149_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.div8.DU_Q3D3d6.fA.A ));
 sky130_fd_sc_hd__mux2_1 _512_ (.A0(\muldiv.div8.DU_Q3D3d6.fA.SUM ),
    .A1(\muldiv.div8.DU_Q3D3d6.fA.A ),
    .S(_113_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_150_));
 sky130_fd_sc_hd__buf_1 _513_ (.A(_150_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.div8.DU_Q2D2d7.fA.A ));
 sky130_fd_sc_hd__mux2_1 _514_ (.A0(\muldiv.div8.DU_Q2D2d7.fA.SUM ),
    .A1(\muldiv.div8.DU_Q2D2d7.fA.A ),
    .S(_101_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_151_));
 sky130_fd_sc_hd__buf_1 _515_ (.A(_151_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.div8.DU_Q1D1d8_EXT.fA.A ));
 sky130_fd_sc_hd__mux2_1 _516_ (.A0(\muldiv.div8.DU_Q1D1d8_EXT.fA.SUM ),
    .A1(\muldiv.div8.DU_Q1D1d8_EXT.fA.A ),
    .S(_097_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_152_));
 sky130_fd_sc_hd__buf_1 _517_ (.A(_152_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.div8.DU_Q0D0d9_EXT.fA.A ));
 sky130_fd_sc_hd__and2_1 _518_ (.A(_130_),
    .B(\muldiv.div8.DU_Q7D7d3.fA.SUM ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_153_));
 sky130_fd_sc_hd__buf_1 _519_ (.A(_153_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.div8.DU_Q6D6d4.fA.A ));
 sky130_fd_sc_hd__a21o_1 _520_ (.A1(net77),
    .A2(\muldiv.div8.DU_Q7D7d3.fA.SUM ),
    .B1(_118_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_154_));
 sky130_fd_sc_hd__or2b_1 _521_ (.A(\muldiv.div8.DU_Q6D6d4.fA.SUM ),
    .B_N(net73),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_155_));
 sky130_fd_sc_hd__and2_1 _522_ (.A(_154_),
    .B(_155_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_156_));
 sky130_fd_sc_hd__buf_1 _523_ (.A(_156_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.div8.DU_Q5D5d5.fA.A ));
 sky130_fd_sc_hd__and2_1 _524_ (.A(net70),
    .B(\muldiv.div8.DU_Q5D5d5.fA.SUM ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_157_));
 sky130_fd_sc_hd__a31o_1 _525_ (.A1(_120_),
    .A2(_154_),
    .A3(_155_),
    .B1(_157_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.div8.DU_Q4D4d6.fA.A ));
 sky130_fd_sc_hd__mux2_1 _526_ (.A0(\muldiv.div8.DU_Q4D4d6.fA.SUM ),
    .A1(\muldiv.div8.DU_Q4D4d6.fA.A ),
    .S(_110_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_158_));
 sky130_fd_sc_hd__buf_1 _527_ (.A(_158_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.div8.DU_Q3D3d7.fA.A ));
 sky130_fd_sc_hd__mux2_1 _528_ (.A0(\muldiv.div8.DU_Q3D3d7.fA.SUM ),
    .A1(\muldiv.div8.DU_Q3D3d7.fA.A ),
    .S(_113_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_159_));
 sky130_fd_sc_hd__buf_1 _529_ (.A(_159_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.div8.DU_Q2D2d8_EXT.fA.A ));
 sky130_fd_sc_hd__mux2_1 _530_ (.A0(\muldiv.div8.DU_Q2D2d8_EXT.fA.SUM ),
    .A1(\muldiv.div8.DU_Q2D2d8_EXT.fA.A ),
    .S(_101_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_160_));
 sky130_fd_sc_hd__buf_1 _531_ (.A(_160_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.div8.DU_Q1D1d9_EXT.fA.A ));
 sky130_fd_sc_hd__mux2_1 _532_ (.A0(\muldiv.div8.DU_Q1D1d9_EXT.fA.SUM ),
    .A1(\muldiv.div8.DU_Q1D1d9_EXT.fA.A ),
    .S(_097_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_161_));
 sky130_fd_sc_hd__buf_1 _533_ (.A(_161_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.div8.DU_Q0D0d10_EXT.fA.A ));
 sky130_fd_sc_hd__and2_1 _534_ (.A(_130_),
    .B(\muldiv.div8.DU_Q7D7d4.fA.SUM ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_162_));
 sky130_fd_sc_hd__buf_1 _535_ (.A(_162_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.div8.DU_Q6D6d5.fA.A ));
 sky130_fd_sc_hd__a21o_1 _536_ (.A1(net72),
    .A2(\muldiv.div8.DU_Q7D7d4.fA.SUM ),
    .B1(net76),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_163_));
 sky130_fd_sc_hd__or2b_1 _537_ (.A(\muldiv.div8.DU_Q6D6d5.fA.SUM ),
    .B_N(\muldiv.div8.DU_Q6D6d0.io_sel ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_164_));
 sky130_fd_sc_hd__and2_1 _538_ (.A(_163_),
    .B(_164_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_165_));
 sky130_fd_sc_hd__buf_1 _539_ (.A(_165_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.div8.DU_Q5D5d6.fA.A ));
 sky130_fd_sc_hd__and2_1 _540_ (.A(net70),
    .B(\muldiv.div8.DU_Q5D5d6.fA.SUM ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_166_));
 sky130_fd_sc_hd__a31o_1 _541_ (.A1(_120_),
    .A2(_163_),
    .A3(_164_),
    .B1(_166_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.div8.DU_Q4D4d7.fA.A ));
 sky130_fd_sc_hd__mux2_1 _542_ (.A0(\muldiv.div8.DU_Q4D4d7.fA.SUM ),
    .A1(\muldiv.div8.DU_Q4D4d7.fA.A ),
    .S(_110_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_167_));
 sky130_fd_sc_hd__buf_1 _543_ (.A(_167_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.div8.DU_Q3D3d8_EXT.fA.A ));
 sky130_fd_sc_hd__mux2_1 _544_ (.A0(\muldiv.div8.DU_Q3D3d8_EXT.fA.SUM ),
    .A1(\muldiv.div8.DU_Q3D3d8_EXT.fA.A ),
    .S(_113_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_168_));
 sky130_fd_sc_hd__buf_1 _545_ (.A(_168_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.div8.DU_Q2D2d9_EXT.fA.A ));
 sky130_fd_sc_hd__mux2_1 _546_ (.A0(\muldiv.div8.DU_Q2D2d9_EXT.fA.SUM ),
    .A1(\muldiv.div8.DU_Q2D2d9_EXT.fA.A ),
    .S(_101_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_169_));
 sky130_fd_sc_hd__buf_1 _547_ (.A(_169_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.div8.DU_Q1D1d10_EXT.fA.A ));
 sky130_fd_sc_hd__mux2_1 _548_ (.A0(\muldiv.div8.DU_Q1D1d10_EXT.fA.SUM ),
    .A1(\muldiv.div8.DU_Q1D1d10_EXT.fA.A ),
    .S(_097_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_170_));
 sky130_fd_sc_hd__buf_1 _549_ (.A(_170_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.div8.DU_Q0D0d11_EXT.fA.A ));
 sky130_fd_sc_hd__and2_1 _550_ (.A(net77),
    .B(\muldiv.div8.DU_Q7D7d5.fA.SUM ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_171_));
 sky130_fd_sc_hd__buf_1 _551_ (.A(_171_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.div8.DU_Q6D6d6.fA.A ));
 sky130_fd_sc_hd__a21o_1 _552_ (.A1(net72),
    .A2(\muldiv.div8.DU_Q7D7d5.fA.SUM ),
    .B1(net76),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_172_));
 sky130_fd_sc_hd__or2b_1 _553_ (.A(\muldiv.div8.DU_Q6D6d6.fA.SUM ),
    .B_N(\muldiv.div8.DU_Q6D6d0.io_sel ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_173_));
 sky130_fd_sc_hd__and2_1 _554_ (.A(_172_),
    .B(_173_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_174_));
 sky130_fd_sc_hd__buf_1 _555_ (.A(_174_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.div8.DU_Q5D5d7.fA.A ));
 sky130_fd_sc_hd__and2_1 _556_ (.A(net70),
    .B(\muldiv.div8.DU_Q5D5d7.fA.SUM ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_175_));
 sky130_fd_sc_hd__a31o_1 _557_ (.A1(_120_),
    .A2(_172_),
    .A3(_173_),
    .B1(_175_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.div8.DU_Q4D4d8_EXT.fA.A ));
 sky130_fd_sc_hd__mux2_1 _558_ (.A0(\muldiv.div8.DU_Q4D4d8_EXT.fA.SUM ),
    .A1(\muldiv.div8.DU_Q4D4d8_EXT.fA.A ),
    .S(_110_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_176_));
 sky130_fd_sc_hd__buf_1 _559_ (.A(_176_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.div8.DU_Q3D3d9_EXT.fA.A ));
 sky130_fd_sc_hd__mux2_1 _560_ (.A0(\muldiv.div8.DU_Q3D3d9_EXT.fA.SUM ),
    .A1(\muldiv.div8.DU_Q3D3d9_EXT.fA.A ),
    .S(_113_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_177_));
 sky130_fd_sc_hd__buf_1 _561_ (.A(_177_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.div8.DU_Q2D2d10_EXT.fA.A ));
 sky130_fd_sc_hd__mux2_1 _562_ (.A0(\muldiv.div8.DU_Q2D2d10_EXT.fA.SUM ),
    .A1(\muldiv.div8.DU_Q2D2d10_EXT.fA.A ),
    .S(_101_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_178_));
 sky130_fd_sc_hd__buf_1 _563_ (.A(_178_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.div8.DU_Q1D1d11_EXT.fA.A ));
 sky130_fd_sc_hd__mux2_1 _564_ (.A0(\muldiv.div8.DU_Q1D1d11_EXT.fA.SUM ),
    .A1(\muldiv.div8.DU_Q1D1d11_EXT.fA.A ),
    .S(_097_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_179_));
 sky130_fd_sc_hd__buf_1 _565_ (.A(_179_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.div8.DU_Q0D0d12_EXT.fA.A ));
 sky130_fd_sc_hd__and2_1 _566_ (.A(_130_),
    .B(\muldiv.div8.DU_Q7D7d1.fA.SUM ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_180_));
 sky130_fd_sc_hd__buf_1 _567_ (.A(_180_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.div8.DU_Q6D6d2.fA.A ));
 sky130_fd_sc_hd__a21o_1 _568_ (.A1(net79),
    .A2(\muldiv.div8.DU_Q7D7d1.fA.SUM ),
    .B1(_118_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_181_));
 sky130_fd_sc_hd__or2b_1 _569_ (.A(\muldiv.div8.DU_Q6D6d2.fA.SUM ),
    .B_N(net73),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_182_));
 sky130_fd_sc_hd__and2_1 _570_ (.A(_181_),
    .B(_182_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_183_));
 sky130_fd_sc_hd__buf_1 _571_ (.A(_183_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.div8.DU_Q5D5d3.fA.A ));
 sky130_fd_sc_hd__and2_1 _572_ (.A(\muldiv.div8.DU_Q5D5d0.io_sel ),
    .B(\muldiv.div8.DU_Q5D5d3.fA.SUM ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_184_));
 sky130_fd_sc_hd__a31o_1 _573_ (.A1(_120_),
    .A2(_181_),
    .A3(_182_),
    .B1(_184_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.div8.DU_Q4D4d4.fA.A ));
 sky130_fd_sc_hd__mux2_1 _574_ (.A0(\muldiv.div8.DU_Q4D4d4.fA.SUM ),
    .A1(\muldiv.div8.DU_Q4D4d4.fA.A ),
    .S(_110_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_185_));
 sky130_fd_sc_hd__buf_1 _575_ (.A(_185_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.div8.DU_Q3D3d5.fA.A ));
 sky130_fd_sc_hd__mux2_1 _576_ (.A0(\muldiv.div8.DU_Q3D3d5.fA.SUM ),
    .A1(\muldiv.div8.DU_Q3D3d5.fA.A ),
    .S(_113_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_186_));
 sky130_fd_sc_hd__buf_1 _577_ (.A(_186_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.div8.DU_Q2D2d6.fA.A ));
 sky130_fd_sc_hd__mux2_1 _578_ (.A0(\muldiv.div8.DU_Q2D2d6.fA.SUM ),
    .A1(\muldiv.div8.DU_Q2D2d6.fA.A ),
    .S(_101_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_187_));
 sky130_fd_sc_hd__buf_1 _579_ (.A(_187_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.div8.DU_Q1D1d7.fA.A ));
 sky130_fd_sc_hd__mux2_1 _580_ (.A0(\muldiv.div8.DU_Q1D1d7.fA.SUM ),
    .A1(\muldiv.div8.DU_Q1D1d7.fA.A ),
    .S(_097_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_188_));
 sky130_fd_sc_hd__buf_1 _581_ (.A(_188_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.div8.DU_Q0D0d8_EXT.fA.A ));
 sky130_fd_sc_hd__and2_1 _582_ (.A(\muldiv.div8.DU_Q7D7d0.io_sel ),
    .B(\muldiv.div8.DU_Q7D7d6.fA.SUM ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_189_));
 sky130_fd_sc_hd__buf_1 _583_ (.A(_189_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.div8.DU_Q6D6d7.fA.A ));
 sky130_fd_sc_hd__mux2_1 _584_ (.A0(\muldiv.div8.DU_Q6D6d7.fA.A ),
    .A1(\muldiv.div8.DU_Q6D6d7.fA.SUM ),
    .S(net74),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_190_));
 sky130_fd_sc_hd__buf_1 _585_ (.A(_190_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.div8.DU_Q5D5d8_EXT.fA.A ));
 sky130_fd_sc_hd__mux2_1 _586_ (.A0(\muldiv.div8.DU_Q5D5d8_EXT.fA.SUM ),
    .A1(\muldiv.div8.DU_Q5D5d8_EXT.fA.A ),
    .S(_120_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_191_));
 sky130_fd_sc_hd__buf_1 _587_ (.A(_191_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.div8.DU_Q4D4d9_EXT.fA.A ));
 sky130_fd_sc_hd__mux2_1 _588_ (.A0(\muldiv.div8.DU_Q4D4d9_EXT.fA.SUM ),
    .A1(\muldiv.div8.DU_Q4D4d9_EXT.fA.A ),
    .S(_110_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_192_));
 sky130_fd_sc_hd__buf_1 _589_ (.A(_192_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.div8.DU_Q3D3d10_EXT.fA.A ));
 sky130_fd_sc_hd__mux2_1 _590_ (.A0(\muldiv.div8.DU_Q3D3d10_EXT.fA.SUM ),
    .A1(\muldiv.div8.DU_Q3D3d10_EXT.fA.A ),
    .S(_113_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_193_));
 sky130_fd_sc_hd__buf_1 _591_ (.A(_193_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.div8.DU_Q2D2d11_EXT.fA.A ));
 sky130_fd_sc_hd__mux2_1 _592_ (.A0(\muldiv.div8.DU_Q2D2d11_EXT.fA.SUM ),
    .A1(\muldiv.div8.DU_Q2D2d11_EXT.fA.A ),
    .S(_101_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_194_));
 sky130_fd_sc_hd__buf_1 _593_ (.A(_194_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.div8.DU_Q1D1d12_EXT.fA.A ));
 sky130_fd_sc_hd__inv_2 _594_ (.A(net10),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_195_));
 sky130_fd_sc_hd__nor2_2 _595_ (.A(net13),
    .B(_195_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_196_));
 sky130_fd_sc_hd__clkbuf_4 _596_ (.A(net10),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_197_));
 sky130_fd_sc_hd__and2_2 _597_ (.A(net13),
    .B(_197_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_198_));
 sky130_fd_sc_hd__a22o_1 _598_ (.A1(\muldiv.mul8.FA_P8A1B7.SUM ),
    .A2(_196_),
    .B1(_198_),
    .B2(\muldiv.div8.HAQ0_SIGN.SUM ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_199_));
 sky130_fd_sc_hd__and2_2 _599_ (.A(net13),
    .B(_195_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_200_));
 sky130_fd_sc_hd__nor2_2 _600_ (.A(net13),
    .B(net10),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_201_));
 sky130_fd_sc_hd__a31o_1 _601_ (.A1(_023_),
    .A2(\muldiv.a1_0.Q ),
    .A3(_201_),
    .B1(net11),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_202_));
 sky130_fd_sc_hd__a21o_1 _602_ (.A1(\muldiv.div8.HAR0_SIGN.SUM ),
    .A2(_200_),
    .B1(_202_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_203_));
 sky130_fd_sc_hd__mux2_1 _603_ (.A0(\muldiv.regR[0] ),
    .A1(\muldiv.regR[8] ),
    .S(_197_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_204_));
 sky130_fd_sc_hd__inv_2 _604_ (.A(net11),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_205_));
 sky130_fd_sc_hd__o22a_4 _605_ (.A1(_199_),
    .A2(_203_),
    .B1(_204_),
    .B2(_205_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[0]));
 sky130_fd_sc_hd__and2_1 _606_ (.A(\muldiv.mul8.FA_P9A2B7.SUM ),
    .B(_196_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_206_));
 sky130_fd_sc_hd__a221o_1 _607_ (.A1(net13),
    .A2(\muldiv.div8.HAR1_SIGN.SUM ),
    .B1(_201_),
    .B2(\muldiv.mul8.HA_P1A0B1.SUM ),
    .C1(_206_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_207_));
 sky130_fd_sc_hd__mux2_1 _608_ (.A0(_207_),
    .A1(\muldiv.div8.HAQ1_SIGN.SUM ),
    .S(_198_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_208_));
 sky130_fd_sc_hd__mux2_1 _609_ (.A0(\muldiv.regR[1] ),
    .A1(\muldiv.regR[9] ),
    .S(_197_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_209_));
 sky130_fd_sc_hd__mux2_1 _610_ (.A0(_208_),
    .A1(_209_),
    .S(net11),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_210_));
 sky130_fd_sc_hd__clkbuf_4 _611_ (.A(_210_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[1]));
 sky130_fd_sc_hd__buf_2 _612_ (.A(_196_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_211_));
 sky130_fd_sc_hd__clkbuf_4 _613_ (.A(_198_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_212_));
 sky130_fd_sc_hd__a22o_1 _614_ (.A1(\muldiv.mul8.FA_P10A3B7.SUM ),
    .A2(_211_),
    .B1(_212_),
    .B2(\muldiv.div8.HAQ2_SIGN.SUM ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_213_));
 sky130_fd_sc_hd__a221o_1 _615_ (.A1(\muldiv.div8.HAR2_SIGN.SUM ),
    .A2(_200_),
    .B1(_201_),
    .B2(\muldiv.mul8.HA_P2A0B2.SUM ),
    .C1(net11),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_214_));
 sky130_fd_sc_hd__and2_1 _616_ (.A(_195_),
    .B(net90),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_215_));
 sky130_fd_sc_hd__a211o_1 _617_ (.A1(_197_),
    .A2(\muldiv.regR[10] ),
    .B1(_215_),
    .C1(_205_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_216_));
 sky130_fd_sc_hd__o21a_4 _618_ (.A1(_213_),
    .A2(_214_),
    .B1(_216_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[2]));
 sky130_fd_sc_hd__a22o_1 _619_ (.A1(\muldiv.mul8.FA_P11A4B7.SUM ),
    .A2(_211_),
    .B1(_212_),
    .B2(\muldiv.div8.HAQ3_SIGN.SUM ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_217_));
 sky130_fd_sc_hd__a221o_1 _620_ (.A1(\muldiv.div8.HAR3_SIGN.SUM ),
    .A2(_200_),
    .B1(_201_),
    .B2(\muldiv.mul8.HA_P3A0B3.SUM ),
    .C1(net11),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_218_));
 sky130_fd_sc_hd__and2_1 _621_ (.A(_195_),
    .B(net91),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_219_));
 sky130_fd_sc_hd__a211o_1 _622_ (.A1(_197_),
    .A2(\muldiv.regR[11] ),
    .B1(_219_),
    .C1(_205_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_220_));
 sky130_fd_sc_hd__o21a_4 _623_ (.A1(_217_),
    .A2(_218_),
    .B1(_220_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[3]));
 sky130_fd_sc_hd__a22o_1 _624_ (.A1(\muldiv.mul8.FA_P12A5B7.SUM ),
    .A2(_211_),
    .B1(_198_),
    .B2(\muldiv.div8.HAQ4_SIGN.SUM ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_221_));
 sky130_fd_sc_hd__a221o_1 _625_ (.A1(\muldiv.div8.HAR4_SIGN.SUM ),
    .A2(_200_),
    .B1(_201_),
    .B2(\muldiv.mul8.HA_P4A0B4.SUM ),
    .C1(net11),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_222_));
 sky130_fd_sc_hd__and2_1 _626_ (.A(_195_),
    .B(net95),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_223_));
 sky130_fd_sc_hd__a211o_1 _627_ (.A1(_197_),
    .A2(\muldiv.regR[12] ),
    .B1(_223_),
    .C1(_205_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_224_));
 sky130_fd_sc_hd__o21a_4 _628_ (.A1(_221_),
    .A2(_222_),
    .B1(_224_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[4]));
 sky130_fd_sc_hd__a22o_1 _629_ (.A1(\muldiv.mul8.FA_P13A6B7.SUM ),
    .A2(_196_),
    .B1(_198_),
    .B2(\muldiv.div8.HAQ5_SIGN.SUM ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_225_));
 sky130_fd_sc_hd__a221o_1 _630_ (.A1(\muldiv.div8.HAR5_SIGN.SUM ),
    .A2(_200_),
    .B1(_201_),
    .B2(\muldiv.mul8.HA_P5A0B5.SUM ),
    .C1(net11),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_226_));
 sky130_fd_sc_hd__and2_1 _631_ (.A(_195_),
    .B(net93),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_227_));
 sky130_fd_sc_hd__a211o_1 _632_ (.A1(_197_),
    .A2(\muldiv.regR[13] ),
    .B1(_227_),
    .C1(_205_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_228_));
 sky130_fd_sc_hd__o21a_2 _633_ (.A1(_225_),
    .A2(_226_),
    .B1(_228_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[5]));
 sky130_fd_sc_hd__a22o_1 _634_ (.A1(\muldiv.mul8.FA_P14A7B7.SUM ),
    .A2(_196_),
    .B1(_198_),
    .B2(\muldiv.div8.HAQ6_SIGN.SUM ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_229_));
 sky130_fd_sc_hd__a221o_1 _635_ (.A1(\muldiv.div8.HAR6_SIGN.SUM ),
    .A2(_200_),
    .B1(_201_),
    .B2(\muldiv.mul8.HA_P6A0B6.SUM ),
    .C1(net11),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_230_));
 sky130_fd_sc_hd__and2_1 _636_ (.A(_195_),
    .B(net94),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_231_));
 sky130_fd_sc_hd__a211o_1 _637_ (.A1(_197_),
    .A2(\muldiv.regR[14] ),
    .B1(_231_),
    .C1(_205_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_232_));
 sky130_fd_sc_hd__o21a_2 _638_ (.A1(_229_),
    .A2(_230_),
    .B1(_232_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[6]));
 sky130_fd_sc_hd__a22o_1 _639_ (.A1(\muldiv.mul8.FA_P15A7B7.SUM ),
    .A2(_196_),
    .B1(_198_),
    .B2(\muldiv.div8.HAQ7_SIGN.SUM ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_233_));
 sky130_fd_sc_hd__a221o_1 _640_ (.A1(\muldiv.div8.HAR7_SIGN.SUM ),
    .A2(_200_),
    .B1(_201_),
    .B2(\muldiv.mul8.FA_P7A0B7.SUM ),
    .C1(net11),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_234_));
 sky130_fd_sc_hd__and2_1 _641_ (.A(_195_),
    .B(net92),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_235_));
 sky130_fd_sc_hd__a211o_1 _642_ (.A1(_197_),
    .A2(\muldiv.regR[15] ),
    .B1(_235_),
    .C1(_205_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_236_));
 sky130_fd_sc_hd__o21a_4 _643_ (.A1(_233_),
    .A2(_234_),
    .B1(_236_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[7]));
 sky130_fd_sc_hd__o22a_1 _644_ (.A1(\muldiv.a1_7.Q ),
    .A2(_021_),
    .B1(_022_),
    .B2(_020_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_237_));
 sky130_fd_sc_hd__buf_4 _645_ (.A(_237_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_238_));
 sky130_fd_sc_hd__inv_2 _646_ (.A(_238_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\muldiv.div8.HAQ0_SIGN.B ));
 sky130_fd_sc_hd__xnor2_1 _647_ (.A(_030_),
    .B(_091_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\muldiv.div8.HAD_DVD_TWOS_0.A ));
 sky130_fd_sc_hd__xnor2_1 _648_ (.A(\muldiv.a1_1.Q ),
    .B(_091_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\muldiv.div8.HAD_DVD_TWOS_1.A ));
 sky130_fd_sc_hd__xnor2_1 _649_ (.A(\muldiv.a1_2.Q ),
    .B(_091_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\muldiv.div8.HAD_DVD_TWOS_2.A ));
 sky130_fd_sc_hd__xnor2_1 _650_ (.A(\muldiv.a1_3.Q ),
    .B(_091_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\muldiv.div8.HAD_DVD_TWOS_3.A ));
 sky130_fd_sc_hd__xnor2_1 _651_ (.A(\muldiv.a1_4.Q ),
    .B(_091_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\muldiv.div8.HAD_DVD_TWOS_4.A ));
 sky130_fd_sc_hd__xnor2_1 _652_ (.A(\muldiv.a1_5.Q ),
    .B(net75),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\muldiv.div8.HAD_DVD_TWOS_5.A ));
 sky130_fd_sc_hd__xnor2_1 _653_ (.A(\muldiv.a1_6.Q ),
    .B(net75),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\muldiv.div8.HAD_DVD_TWOS_6.A ));
 sky130_fd_sc_hd__and2b_1 _654_ (.A_N(_081_),
    .B(\muldiv.a1_7.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_239_));
 sky130_fd_sc_hd__clkbuf_2 _655_ (.A(_239_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.div8.HAD_DVD_TWOS_7.A ));
 sky130_fd_sc_hd__xor2_4 _656_ (.A(_023_),
    .B(net22),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.div8.DU_Q0D0d0.fA.B ));
 sky130_fd_sc_hd__xor2_4 _657_ (.A(\muldiv.a0_1.Q ),
    .B(net22),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.div8.DU_Q0D0d1.fA.B ));
 sky130_fd_sc_hd__xor2_4 _658_ (.A(\muldiv.a0_2.Q ),
    .B(net21),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.div8.DU_Q0D0d2.fA.B ));
 sky130_fd_sc_hd__xor2_2 _659_ (.A(\muldiv.a0_3.Q ),
    .B(net21),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.div8.DU_Q0D0d3.fA.B ));
 sky130_fd_sc_hd__xor2_2 _660_ (.A(\muldiv.a0_4.Q ),
    .B(net21),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.div8.DU_Q0D0d4.fA.B ));
 sky130_fd_sc_hd__xor2_2 _661_ (.A(\muldiv.a0_5.Q ),
    .B(net21),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.div8.DU_Q0D0d5.fA.B ));
 sky130_fd_sc_hd__xor2_2 _662_ (.A(\muldiv.a0_6.Q ),
    .B(net21),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.div8.DU_Q0D0d6.fA.B ));
 sky130_fd_sc_hd__or2b_1 _663_ (.A(_081_),
    .B_N(_073_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_240_));
 sky130_fd_sc_hd__clkbuf_8 _664_ (.A(_240_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.div8.DU_Q0D0d7.fA.B ));
 sky130_fd_sc_hd__mux2_4 _665_ (.A0(\muldiv.div8.DU_Q0D0d0.fA.A ),
    .A1(\muldiv.div8.DU_Q0D0d0.fA.SUM ),
    .S(\muldiv.div8.DU_Q0D0d0.io_sel ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_241_));
 sky130_fd_sc_hd__xnor2_2 _666_ (.A(net75),
    .B(_241_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\muldiv.div8.HAR0_SIGN.A ));
 sky130_fd_sc_hd__mux2_1 _667_ (.A0(\muldiv.div8.DU_Q0D0d1.fA.A ),
    .A1(\muldiv.div8.DU_Q0D0d1.fA.SUM ),
    .S(\muldiv.div8.DU_Q0D0d0.io_sel ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_242_));
 sky130_fd_sc_hd__xnor2_1 _668_ (.A(net75),
    .B(_242_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\muldiv.div8.HAR1_SIGN.A ));
 sky130_fd_sc_hd__mux2_1 _669_ (.A0(\muldiv.div8.DU_Q0D0d2.fA.A ),
    .A1(\muldiv.div8.DU_Q0D0d2.fA.SUM ),
    .S(\muldiv.div8.DU_Q0D0d0.io_sel ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_243_));
 sky130_fd_sc_hd__xnor2_1 _670_ (.A(_022_),
    .B(_243_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\muldiv.div8.HAR2_SIGN.A ));
 sky130_fd_sc_hd__mux2_1 _671_ (.A0(\muldiv.div8.DU_Q0D0d3.fA.A ),
    .A1(\muldiv.div8.DU_Q0D0d3.fA.SUM ),
    .S(\muldiv.div8.DU_Q0D0d0.io_sel ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_244_));
 sky130_fd_sc_hd__xnor2_1 _672_ (.A(_022_),
    .B(_244_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\muldiv.div8.HAR3_SIGN.A ));
 sky130_fd_sc_hd__mux2_1 _673_ (.A0(\muldiv.div8.DU_Q0D0d4.fA.A ),
    .A1(\muldiv.div8.DU_Q0D0d4.fA.SUM ),
    .S(net67),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_245_));
 sky130_fd_sc_hd__xnor2_1 _674_ (.A(net71),
    .B(_245_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\muldiv.div8.HAR4_SIGN.A ));
 sky130_fd_sc_hd__mux2_1 _675_ (.A0(\muldiv.div8.DU_Q0D0d5.fA.A ),
    .A1(\muldiv.div8.DU_Q0D0d5.fA.SUM ),
    .S(net67),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_246_));
 sky130_fd_sc_hd__xnor2_1 _676_ (.A(net71),
    .B(_246_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\muldiv.div8.HAR5_SIGN.A ));
 sky130_fd_sc_hd__mux2_1 _677_ (.A0(\muldiv.div8.DU_Q0D0d6.fA.A ),
    .A1(\muldiv.div8.DU_Q0D0d6.fA.SUM ),
    .S(net67),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_247_));
 sky130_fd_sc_hd__xnor2_1 _678_ (.A(net71),
    .B(_247_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\muldiv.div8.HAR6_SIGN.A ));
 sky130_fd_sc_hd__or2b_1 _679_ (.A(\muldiv.div8.DU_Q0D0d7.fA.SUM ),
    .B_N(net67),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_248_));
 sky130_fd_sc_hd__o31a_1 _680_ (.A1(net67),
    .A2(_141_),
    .A3(_142_),
    .B1(_248_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_249_));
 sky130_fd_sc_hd__xnor2_1 _681_ (.A(net71),
    .B(_249_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\muldiv.div8.HAR7_SIGN.A ));
 sky130_fd_sc_hd__xnor2_2 _682_ (.A(\muldiv.div8.DU_Q0D0d0.io_sel ),
    .B(_238_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\muldiv.div8.HAQ0_SIGN.A ));
 sky130_fd_sc_hd__xnor2_1 _683_ (.A(\muldiv.div8.DU_Q1D1d0.io_sel ),
    .B(_238_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\muldiv.div8.HAQ1_SIGN.A ));
 sky130_fd_sc_hd__xnor2_1 _684_ (.A(\muldiv.div8.DU_Q2D2d0.io_sel ),
    .B(_238_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\muldiv.div8.HAQ2_SIGN.A ));
 sky130_fd_sc_hd__xnor2_1 _685_ (.A(\muldiv.div8.DU_Q3D3d0.io_sel ),
    .B(_238_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\muldiv.div8.HAQ3_SIGN.A ));
 sky130_fd_sc_hd__xnor2_1 _686_ (.A(\muldiv.div8.DU_Q4D4d0.io_sel ),
    .B(_238_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\muldiv.div8.HAQ4_SIGN.A ));
 sky130_fd_sc_hd__xnor2_1 _687_ (.A(net68),
    .B(_238_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\muldiv.div8.HAQ5_SIGN.A ));
 sky130_fd_sc_hd__xnor2_1 _688_ (.A(net76),
    .B(_238_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\muldiv.div8.HAQ6_SIGN.A ));
 sky130_fd_sc_hd__xnor2_1 _689_ (.A(net77),
    .B(_238_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\muldiv.div8.HAQ7_SIGN.A ));
 sky130_fd_sc_hd__or4_1 _690_ (.A(\muldiv.a0_7.Q ),
    .B(\muldiv.a0_0.Q ),
    .C(\muldiv.a0_1.Q ),
    .D(\muldiv.a0_4.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_250_));
 sky130_fd_sc_hd__or4b_1 _691_ (.A(\muldiv.a0_5.Q ),
    .B(_250_),
    .C(\muldiv.a0_6.Q ),
    .D_N(net13),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_251_));
 sky130_fd_sc_hd__nor3_1 _692_ (.A(\muldiv.a0_2.Q ),
    .B(\muldiv.a0_3.Q ),
    .C(_251_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\muldiv.div8.io_edivzero ));
 sky130_fd_sc_hd__and3_1 _693_ (.A(net77),
    .B(net13),
    .C(\muldiv.div8.DU_Q7D7d7.fA.SUM ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_252_));
 sky130_fd_sc_hd__clkbuf_1 _694_ (.A(_252_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.div8.io_edivoverflow ));
 sky130_fd_sc_hd__mux2_1 _695_ (.A0(\muldiv.div8.HAD_DVD_TWOS_0.B ),
    .A1(\muldiv.div8.HAD_DVD_TWOS_7.A ),
    .S(_023_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_253_));
 sky130_fd_sc_hd__clkbuf_1 _696_ (.A(_253_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.mul8.FA_P7A0B7.B ));
 sky130_fd_sc_hd__mux2_1 _697_ (.A0(\muldiv.div8.HAD_DVD_TWOS_0.B ),
    .A1(\muldiv.div8.HAD_DVD_TWOS_7.A ),
    .S(\muldiv.a0_1.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_254_));
 sky130_fd_sc_hd__buf_1 _698_ (.A(_254_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.mul8.FA_P8A1B7.B ));
 sky130_fd_sc_hd__mux2_1 _699_ (.A0(\muldiv.div8.HAD_DVD_TWOS_0.B ),
    .A1(\muldiv.div8.HAD_DVD_TWOS_7.A ),
    .S(\muldiv.a0_2.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_255_));
 sky130_fd_sc_hd__clkbuf_1 _700_ (.A(_255_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.mul8.FA_P9A2B7.B ));
 sky130_fd_sc_hd__mux2_1 _701_ (.A0(\muldiv.div8.HAD_DVD_TWOS_0.B ),
    .A1(\muldiv.div8.HAD_DVD_TWOS_7.A ),
    .S(\muldiv.a0_3.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_256_));
 sky130_fd_sc_hd__buf_1 _702_ (.A(_256_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.mul8.FA_P10A3B7.B ));
 sky130_fd_sc_hd__mux2_1 _703_ (.A0(\muldiv.div8.HAD_DVD_TWOS_0.B ),
    .A1(\muldiv.div8.HAD_DVD_TWOS_7.A ),
    .S(\muldiv.a0_4.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_257_));
 sky130_fd_sc_hd__clkbuf_1 _704_ (.A(_257_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.mul8.FA_P11A4B7.B ));
 sky130_fd_sc_hd__mux2_1 _705_ (.A0(\muldiv.div8.HAD_DVD_TWOS_0.B ),
    .A1(\muldiv.div8.HAD_DVD_TWOS_7.A ),
    .S(\muldiv.a0_5.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_258_));
 sky130_fd_sc_hd__clkbuf_1 _706_ (.A(_258_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.mul8.FA_P12A5B7.B ));
 sky130_fd_sc_hd__mux2_1 _707_ (.A0(\muldiv.div8.HAD_DVD_TWOS_0.B ),
    .A1(\muldiv.div8.HAD_DVD_TWOS_7.A ),
    .S(\muldiv.a0_6.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_259_));
 sky130_fd_sc_hd__clkbuf_1 _708_ (.A(_259_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.mul8.FA_P13A6B7.B ));
 sky130_fd_sc_hd__inv_2 _709__1 (.A(clknet_1_1__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net66));
 sky130_fd_sc_hd__clkbuf_4 _710_ (.A(_195_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_260_));
 sky130_fd_sc_hd__and3_1 _711_ (.A(_023_),
    .B(_030_),
    .C(_196_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_261_));
 sky130_fd_sc_hd__a221o_1 _712_ (.A1(_260_),
    .A2(net88),
    .B1(_212_),
    .B2(\muldiv.div8.HAR0_SIGN.SUM ),
    .C1(_261_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_003_));
 sky130_fd_sc_hd__and3_1 _713_ (.A(net13),
    .B(\muldiv.div8.HAR1_SIGN.SUM ),
    .C(_197_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_262_));
 sky130_fd_sc_hd__a221o_1 _714_ (.A1(_260_),
    .A2(net87),
    .B1(_211_),
    .B2(\muldiv.mul8.HA_P1A0B1.SUM ),
    .C1(_262_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_004_));
 sky130_fd_sc_hd__a221o_1 _715_ (.A1(\muldiv.mul8.HA_P2A0B2.SUM ),
    .A2(_211_),
    .B1(_212_),
    .B2(\muldiv.div8.HAR2_SIGN.SUM ),
    .C1(_215_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_005_));
 sky130_fd_sc_hd__a221o_1 _716_ (.A1(\muldiv.mul8.HA_P3A0B3.SUM ),
    .A2(_211_),
    .B1(_212_),
    .B2(\muldiv.div8.HAR3_SIGN.SUM ),
    .C1(_219_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_006_));
 sky130_fd_sc_hd__a221o_1 _717_ (.A1(\muldiv.mul8.HA_P4A0B4.SUM ),
    .A2(_211_),
    .B1(_212_),
    .B2(\muldiv.div8.HAR4_SIGN.SUM ),
    .C1(_223_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_007_));
 sky130_fd_sc_hd__a221o_1 _718_ (.A1(\muldiv.mul8.HA_P5A0B5.SUM ),
    .A2(_211_),
    .B1(_212_),
    .B2(\muldiv.div8.HAR5_SIGN.SUM ),
    .C1(_227_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_008_));
 sky130_fd_sc_hd__a221o_1 _719_ (.A1(\muldiv.mul8.HA_P6A0B6.SUM ),
    .A2(_211_),
    .B1(_212_),
    .B2(\muldiv.div8.HAR6_SIGN.SUM ),
    .C1(_231_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_009_));
 sky130_fd_sc_hd__a221o_1 _720_ (.A1(\muldiv.mul8.FA_P7A0B7.SUM ),
    .A2(_211_),
    .B1(_212_),
    .B2(\muldiv.div8.HAR7_SIGN.SUM ),
    .C1(_235_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_010_));
 sky130_fd_sc_hd__a21o_1 _721_ (.A1(_260_),
    .A2(net83),
    .B1(_199_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_011_));
 sky130_fd_sc_hd__a221o_1 _722_ (.A1(_260_),
    .A2(net89),
    .B1(_212_),
    .B2(\muldiv.div8.HAQ1_SIGN.SUM ),
    .C1(_206_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_012_));
 sky130_fd_sc_hd__a21o_1 _723_ (.A1(_260_),
    .A2(net84),
    .B1(_213_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_013_));
 sky130_fd_sc_hd__a21o_1 _724_ (.A1(_260_),
    .A2(net82),
    .B1(_217_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_014_));
 sky130_fd_sc_hd__a21o_1 _725_ (.A1(_260_),
    .A2(net80),
    .B1(_221_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_015_));
 sky130_fd_sc_hd__a21o_1 _726_ (.A1(_260_),
    .A2(net81),
    .B1(_225_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_016_));
 sky130_fd_sc_hd__a21o_1 _727_ (.A1(_260_),
    .A2(net85),
    .B1(_229_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_017_));
 sky130_fd_sc_hd__a21o_1 _728_ (.A1(_260_),
    .A2(net86),
    .B1(_233_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_018_));
 sky130_fd_sc_hd__and2b_1 _729_ (.A_N(\muldiv.div2reg ),
    .B(net23),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_019_));
 sky130_fd_sc_hd__buf_1 _730_ (.A(_019_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_002_));
 sky130_fd_sc_hd__inv_2 _731_ (.A(_002_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_001_));
 sky130_fd_sc_hd__clkbuf_4 _732_ (.A(\muldiv.a0_7.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_020_));
 sky130_fd_sc_hd__nand2_1 _733_ (.A(net12),
    .B(_020_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_021_));
 sky130_fd_sc_hd__buf_1 _734_ (.A(_021_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.div8.DU_Q0D0d0.fA.CIN ));
 sky130_fd_sc_hd__nand2_8 _735_ (.A(net12),
    .B(\muldiv.a1_7.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_022_));
 sky130_fd_sc_hd__inv_2 _736_ (.A(_022_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\muldiv.div8.HAD_DVD_TWOS_0.B ));
 sky130_fd_sc_hd__buf_4 _737_ (.A(\muldiv.a0_0.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_023_));
 sky130_fd_sc_hd__and2_1 _738_ (.A(\muldiv.a1_1.Q ),
    .B(_023_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_024_));
 sky130_fd_sc_hd__clkbuf_1 _739_ (.A(_024_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\muldiv.mul8.A0xB1_8 ));
 sky130_fd_sc_hd__dfxtp_1 _740_ (.CLK(net66),
    .D(_001_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\muldiv.negedgeReg_1.area_io_q ));
 sky130_fd_sc_hd__dfxtp_1 _741_ (.CLK(clknet_1_1__leaf_clk),
    .D(_002_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\muldiv.div2reg ));
 sky130_fd_sc_hd__dfxtp_1 _742_ (.CLK(clknet_1_0__leaf_clk),
    .D(_003_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\muldiv.regR[0] ));
 sky130_fd_sc_hd__dfxtp_1 _743_ (.CLK(clknet_1_1__leaf_clk),
    .D(_004_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\muldiv.regR[1] ));
 sky130_fd_sc_hd__dfxtp_1 _744_ (.CLK(clknet_1_1__leaf_clk),
    .D(_005_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\muldiv.regR[2] ));
 sky130_fd_sc_hd__dfxtp_1 _745_ (.CLK(clknet_1_1__leaf_clk),
    .D(_006_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\muldiv.regR[3] ));
 sky130_fd_sc_hd__dfxtp_1 _746_ (.CLK(clknet_1_1__leaf_clk),
    .D(_007_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\muldiv.regR[4] ));
 sky130_fd_sc_hd__dfxtp_1 _747_ (.CLK(clknet_1_0__leaf_clk),
    .D(_008_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\muldiv.regR[5] ));
 sky130_fd_sc_hd__dfxtp_1 _748_ (.CLK(clknet_1_0__leaf_clk),
    .D(_009_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\muldiv.regR[6] ));
 sky130_fd_sc_hd__dfxtp_1 _749_ (.CLK(clknet_1_0__leaf_clk),
    .D(_010_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\muldiv.regR[7] ));
 sky130_fd_sc_hd__dfxtp_1 _750_ (.CLK(clknet_1_0__leaf_clk),
    .D(_011_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\muldiv.regR[8] ));
 sky130_fd_sc_hd__dfxtp_1 _751_ (.CLK(clknet_1_1__leaf_clk),
    .D(_012_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\muldiv.regR[9] ));
 sky130_fd_sc_hd__dfxtp_1 _752_ (.CLK(clknet_1_0__leaf_clk),
    .D(_013_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\muldiv.regR[10] ));
 sky130_fd_sc_hd__dfxtp_1 _753_ (.CLK(clknet_1_1__leaf_clk),
    .D(_014_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\muldiv.regR[11] ));
 sky130_fd_sc_hd__dfxtp_1 _754_ (.CLK(clknet_1_0__leaf_clk),
    .D(_015_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\muldiv.regR[12] ));
 sky130_fd_sc_hd__dfxtp_1 _755_ (.CLK(clknet_1_0__leaf_clk),
    .D(_016_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\muldiv.regR[13] ));
 sky130_fd_sc_hd__dfxtp_1 _756_ (.CLK(clknet_1_0__leaf_clk),
    .D(_017_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\muldiv.regR[14] ));
 sky130_fd_sc_hd__dfxtp_1 _757_ (.CLK(clknet_1_0__leaf_clk),
    .D(_018_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\muldiv.regR[15] ));
 sky130_fd_sc_hd__buf_2 _799_ (.A(\muldiv.div8.io_edivoverflow ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uio_out[4]));
 sky130_fd_sc_hd__clkbuf_4 _800_ (.A(\muldiv.div8.io_edivzero ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uio_out[5]));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_2 clone10 (.A(net96),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net76));
 sky130_fd_sc_hd__clkbuf_2 clone11 (.A(net78),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net77));
 sky130_fd_sc_hd__nand2_2 clone5 (.A(net12),
    .B(\muldiv.a1_7.Q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net71));
 sky130_fd_sc_hd__buf_4 clone9 (.A(_022_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net75));
 sky130_fd_sc_hd__buf_6 fanout21 (.A(\muldiv.div8.DU_Q0D0d0.fA.CIN ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net21));
 sky130_fd_sc_hd__buf_4 fanout22 (.A(\muldiv.div8.DU_Q0D0d0.fA.CIN ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net22));
 sky130_fd_sc_hd__buf_2 fanout23 (.A(net1),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_2 fanout24 (.A(net1),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net24));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(\muldiv.regR[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net80));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(\muldiv.regR[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net81));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(\muldiv.regR[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net82));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(\muldiv.regR[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net83));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(\muldiv.regR[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net84));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(\muldiv.regR[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net85));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(\muldiv.regR[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net86));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(\muldiv.regR[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net87));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(\muldiv.regR[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net88));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(\muldiv.regR[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net89));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(\muldiv.regR[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net90));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(\muldiv.regR[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net91));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(\muldiv.regR[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net92));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(\muldiv.regR[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net93));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(\muldiv.regR[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net94));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(\muldiv.regR[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net95));
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(rst_n),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net1));
 sky130_fd_sc_hd__buf_1 input10 (.A(uio_in[0]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net10));
 sky130_fd_sc_hd__buf_2 input11 (.A(uio_in[3]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net11));
 sky130_fd_sc_hd__buf_8 input12 (.A(uio_in[6]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net12));
 sky130_fd_sc_hd__buf_2 input13 (.A(uio_in[7]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(ui_in[0]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(ui_in[1]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(ui_in[2]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(ui_in[3]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(ui_in[4]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(ui_in[5]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(ui_in[6]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_1 input9 (.A(ui_in[7]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net9));
 sky130_fd_sc_hd__buf_4 max_cap14 (.A(\muldiv.div8.DU_Q0D0d6.fA.B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net14));
 sky130_fd_sc_hd__buf_4 max_cap15 (.A(\muldiv.div8.DU_Q0D0d5.fA.B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net15));
 sky130_fd_sc_hd__buf_4 max_cap16 (.A(\muldiv.div8.DU_Q0D0d4.fA.B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net16));
 sky130_fd_sc_hd__buf_4 max_cap17 (.A(\muldiv.div8.DU_Q0D0d3.fA.B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net17));
 sky130_fd_sc_hd__buf_4 max_cap18 (.A(\muldiv.div8.DU_Q0D0d2.fA.B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net18));
 sky130_fd_sc_hd__buf_4 max_cap19 (.A(\muldiv.div8.DU_Q0D0d1.fA.B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net19));
 sky130_fd_sc_hd__buf_4 max_cap20 (.A(\muldiv.div8.DU_Q0D0d0.fA.B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net20));
 sky130_fd_sc_hd__dlrtp_1 \muldiv.a0_0.genblk1.dlrtp_1  (.D(net2),
    .GATE(\muldiv.a0_0.GATE ),
    .RESET_B(net23),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\muldiv.a0_0.Q ));
 sky130_fd_sc_hd__dlrtp_4 \muldiv.a0_1.genblk1.dlrtp_1  (.D(net3),
    .GATE(\muldiv.a0_0.GATE ),
    .RESET_B(net24),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\muldiv.a0_1.Q ));
 sky130_fd_sc_hd__dlrtp_4 \muldiv.a0_2.genblk1.dlrtp_1  (.D(net4),
    .GATE(\muldiv.a0_0.GATE ),
    .RESET_B(net24),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\muldiv.a0_2.Q ));
 sky130_fd_sc_hd__dlrtp_4 \muldiv.a0_3.genblk1.dlrtp_1  (.D(net5),
    .GATE(\muldiv.a0_0.GATE ),
    .RESET_B(net24),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\muldiv.a0_3.Q ));
 sky130_fd_sc_hd__dlrtp_4 \muldiv.a0_4.genblk1.dlrtp_1  (.D(net6),
    .GATE(\muldiv.a0_0.GATE ),
    .RESET_B(net23),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\muldiv.a0_4.Q ));
 sky130_fd_sc_hd__dlrtp_4 \muldiv.a0_5.genblk1.dlrtp_1  (.D(net7),
    .GATE(\muldiv.a0_0.GATE ),
    .RESET_B(net23),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\muldiv.a0_5.Q ));
 sky130_fd_sc_hd__dlrtp_4 \muldiv.a0_6.genblk1.dlrtp_1  (.D(net8),
    .GATE(\muldiv.a0_0.GATE ),
    .RESET_B(net23),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\muldiv.a0_6.Q ));
 sky130_fd_sc_hd__dlrtp_1 \muldiv.a0_7.genblk1.dlrtp_1  (.D(net9),
    .GATE(\muldiv.a0_0.GATE ),
    .RESET_B(net23),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\muldiv.a0_7.Q ));
 sky130_fd_sc_hd__dlrtp_1 \muldiv.a1_0.genblk1.dlrtp_1  (.D(net2),
    .GATE(\muldiv.a1_0.GATE ),
    .RESET_B(net24),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\muldiv.a1_0.Q ));
 sky130_fd_sc_hd__dlrtp_4 \muldiv.a1_1.genblk1.dlrtp_1  (.D(net3),
    .GATE(\muldiv.a1_0.GATE ),
    .RESET_B(net24),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\muldiv.a1_1.Q ));
 sky130_fd_sc_hd__dlrtp_4 \muldiv.a1_2.genblk1.dlrtp_1  (.D(net4),
    .GATE(\muldiv.a1_0.GATE ),
    .RESET_B(net24),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\muldiv.a1_2.Q ));
 sky130_fd_sc_hd__dlrtp_4 \muldiv.a1_3.genblk1.dlrtp_1  (.D(net5),
    .GATE(\muldiv.a1_0.GATE ),
    .RESET_B(net24),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\muldiv.a1_3.Q ));
 sky130_fd_sc_hd__dlrtp_2 \muldiv.a1_4.genblk1.dlrtp_1  (.D(net6),
    .GATE(\muldiv.a1_0.GATE ),
    .RESET_B(net23),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\muldiv.a1_4.Q ));
 sky130_fd_sc_hd__dlrtp_2 \muldiv.a1_5.genblk1.dlrtp_1  (.D(net7),
    .GATE(\muldiv.a1_0.GATE ),
    .RESET_B(net23),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\muldiv.a1_5.Q ));
 sky130_fd_sc_hd__dlrtp_2 \muldiv.a1_6.genblk1.dlrtp_1  (.D(net8),
    .GATE(\muldiv.a1_0.GATE ),
    .RESET_B(net23),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\muldiv.a1_6.Q ));
 sky130_fd_sc_hd__dlrtp_2 \muldiv.a1_7.genblk1.dlrtp_1  (.D(net9),
    .GATE(\muldiv.a1_0.GATE ),
    .RESET_B(net23),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\muldiv.a1_7.Q ));
 sky130_fd_sc_hd__fa_1 \muldiv.div8.DU_Q0D0d0.fA.genblk1.fa_1  (.A(\muldiv.div8.DU_Q0D0d0.fA.A ),
    .B(\muldiv.div8.DU_Q0D0d0.fA.B ),
    .CIN(net22),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.div8.DU_Q0D0d0.fA.COUT ),
    .SUM(\muldiv.div8.DU_Q0D0d0.fA.SUM ));
 sky130_fd_sc_hd__fa_2 \muldiv.div8.DU_Q0D0d1.fA.genblk1.fa_1  (.A(\muldiv.div8.DU_Q0D0d1.fA.A ),
    .B(\muldiv.div8.DU_Q0D0d1.fA.B ),
    .CIN(\muldiv.div8.DU_Q0D0d0.fA.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.div8.DU_Q0D0d1.fA.COUT ),
    .SUM(\muldiv.div8.DU_Q0D0d1.fA.SUM ));
 sky130_fd_sc_hd__fa_2 \muldiv.div8.DU_Q0D0d10_EXT.fA.genblk1.fa_1  (.A(\muldiv.div8.DU_Q0D0d10_EXT.fA.A ),
    .B(net44),
    .CIN(\muldiv.div8.DU_Q0D0d10_EXT.fA.CIN ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.div8.DU_Q0D0d10_EXT.fA.COUT ),
    .SUM(\muldiv.div8.DU_Q0D0d10_EXT.fA.SUM ));
 sky130_fd_sc_hd__conb_1 \muldiv.div8.DU_Q0D0d10_EXT.fA.genblk1.fa_1_44  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(net44));
 sky130_fd_sc_hd__fa_2 \muldiv.div8.DU_Q0D0d11_EXT.fA.genblk1.fa_1  (.A(\muldiv.div8.DU_Q0D0d11_EXT.fA.A ),
    .B(net45),
    .CIN(\muldiv.div8.DU_Q0D0d10_EXT.fA.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.div8.DU_Q0D0d11_EXT.fA.COUT ),
    .SUM(\muldiv.div8.DU_Q0D0d11_EXT.fA.SUM ));
 sky130_fd_sc_hd__conb_1 \muldiv.div8.DU_Q0D0d11_EXT.fA.genblk1.fa_1_45  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(net45));
 sky130_fd_sc_hd__fa_2 \muldiv.div8.DU_Q0D0d12_EXT.fA.genblk1.fa_1  (.A(\muldiv.div8.DU_Q0D0d12_EXT.fA.A ),
    .B(net46),
    .CIN(\muldiv.div8.DU_Q0D0d11_EXT.fA.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.div8.DU_Q0D0d0.io_sel ),
    .SUM(\muldiv.div8.DU_Q0D0d12_EXT.fA.SUM ));
 sky130_fd_sc_hd__conb_1 \muldiv.div8.DU_Q0D0d12_EXT.fA.genblk1.fa_1_46  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(net46));
 sky130_fd_sc_hd__fa_2 \muldiv.div8.DU_Q0D0d2.fA.genblk1.fa_1  (.A(\muldiv.div8.DU_Q0D0d2.fA.A ),
    .B(net18),
    .CIN(\muldiv.div8.DU_Q0D0d1.fA.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.div8.DU_Q0D0d2.fA.COUT ),
    .SUM(\muldiv.div8.DU_Q0D0d2.fA.SUM ));
 sky130_fd_sc_hd__fa_2 \muldiv.div8.DU_Q0D0d3.fA.genblk1.fa_1  (.A(\muldiv.div8.DU_Q0D0d3.fA.A ),
    .B(net17),
    .CIN(\muldiv.div8.DU_Q0D0d2.fA.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.div8.DU_Q0D0d3.fA.COUT ),
    .SUM(\muldiv.div8.DU_Q0D0d3.fA.SUM ));
 sky130_fd_sc_hd__fa_2 \muldiv.div8.DU_Q0D0d4.fA.genblk1.fa_1  (.A(\muldiv.div8.DU_Q0D0d4.fA.A ),
    .B(net16),
    .CIN(\muldiv.div8.DU_Q0D0d3.fA.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.div8.DU_Q0D0d4.fA.COUT ),
    .SUM(\muldiv.div8.DU_Q0D0d4.fA.SUM ));
 sky130_fd_sc_hd__fa_2 \muldiv.div8.DU_Q0D0d5.fA.genblk1.fa_1  (.A(\muldiv.div8.DU_Q0D0d5.fA.A ),
    .B(net15),
    .CIN(\muldiv.div8.DU_Q0D0d4.fA.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.div8.DU_Q0D0d5.fA.COUT ),
    .SUM(\muldiv.div8.DU_Q0D0d5.fA.SUM ));
 sky130_fd_sc_hd__fa_2 \muldiv.div8.DU_Q0D0d6.fA.genblk1.fa_1  (.A(\muldiv.div8.DU_Q0D0d6.fA.A ),
    .B(net14),
    .CIN(\muldiv.div8.DU_Q0D0d5.fA.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.div8.DU_Q0D0d6.fA.COUT ),
    .SUM(\muldiv.div8.DU_Q0D0d6.fA.SUM ));
 sky130_fd_sc_hd__fa_2 \muldiv.div8.DU_Q0D0d7.fA.genblk1.fa_1  (.A(\muldiv.div8.DU_Q0D0d7.fA.A ),
    .B(\muldiv.div8.DU_Q0D0d7.fA.B ),
    .CIN(\muldiv.div8.DU_Q0D0d6.fA.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.div8.DU_Q0D0d7.fA.COUT ),
    .SUM(\muldiv.div8.DU_Q0D0d7.fA.SUM ));
 sky130_fd_sc_hd__fa_2 \muldiv.div8.DU_Q0D0d8_EXT.fA.genblk1.fa_1  (.A(\muldiv.div8.DU_Q0D0d8_EXT.fA.A ),
    .B(net47),
    .CIN(\muldiv.div8.DU_Q0D0d7.fA.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.div8.DU_Q0D0d8_EXT.fA.COUT ),
    .SUM(\muldiv.div8.DU_Q0D0d8_EXT.fA.SUM ));
 sky130_fd_sc_hd__conb_1 \muldiv.div8.DU_Q0D0d8_EXT.fA.genblk1.fa_1_47  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(net47));
 sky130_fd_sc_hd__fa_2 \muldiv.div8.DU_Q0D0d9_EXT.fA.genblk1.fa_1  (.A(\muldiv.div8.DU_Q0D0d9_EXT.fA.A ),
    .B(net48),
    .CIN(\muldiv.div8.DU_Q0D0d8_EXT.fA.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.div8.DU_Q0D0d10_EXT.fA.CIN ),
    .SUM(\muldiv.div8.DU_Q0D0d9_EXT.fA.SUM ));
 sky130_fd_sc_hd__conb_1 \muldiv.div8.DU_Q0D0d9_EXT.fA.genblk1.fa_1_48  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(net48));
 sky130_fd_sc_hd__fa_1 \muldiv.div8.DU_Q1D1d0.fA.genblk1.fa_1  (.A(\muldiv.div8.DU_Q1D1d0.fA.A ),
    .B(\muldiv.div8.DU_Q0D0d0.fA.B ),
    .CIN(net21),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.div8.DU_Q1D1d0.fA.COUT ),
    .SUM(\muldiv.div8.DU_Q1D1d0.fA.SUM ));
 sky130_fd_sc_hd__fa_2 \muldiv.div8.DU_Q1D1d1.fA.genblk1.fa_1  (.A(\muldiv.div8.DU_Q1D1d1.fA.A ),
    .B(\muldiv.div8.DU_Q0D0d1.fA.B ),
    .CIN(\muldiv.div8.DU_Q1D1d0.fA.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.div8.DU_Q1D1d1.fA.COUT ),
    .SUM(\muldiv.div8.DU_Q1D1d1.fA.SUM ));
 sky130_fd_sc_hd__fa_2 \muldiv.div8.DU_Q1D1d10_EXT.fA.genblk1.fa_1  (.A(\muldiv.div8.DU_Q1D1d10_EXT.fA.A ),
    .B(net49),
    .CIN(\muldiv.div8.DU_Q1D1d10_EXT.fA.CIN ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.div8.DU_Q1D1d10_EXT.fA.COUT ),
    .SUM(\muldiv.div8.DU_Q1D1d10_EXT.fA.SUM ));
 sky130_fd_sc_hd__conb_1 \muldiv.div8.DU_Q1D1d10_EXT.fA.genblk1.fa_1_49  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(net49));
 sky130_fd_sc_hd__fa_2 \muldiv.div8.DU_Q1D1d11_EXT.fA.genblk1.fa_1  (.A(\muldiv.div8.DU_Q1D1d11_EXT.fA.A ),
    .B(net50),
    .CIN(\muldiv.div8.DU_Q1D1d10_EXT.fA.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.div8.DU_Q1D1d11_EXT.fA.COUT ),
    .SUM(\muldiv.div8.DU_Q1D1d11_EXT.fA.SUM ));
 sky130_fd_sc_hd__conb_1 \muldiv.div8.DU_Q1D1d11_EXT.fA.genblk1.fa_1_50  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(net50));
 sky130_fd_sc_hd__fa_2 \muldiv.div8.DU_Q1D1d12_EXT.fA.genblk1.fa_1  (.A(\muldiv.div8.DU_Q1D1d12_EXT.fA.A ),
    .B(net51),
    .CIN(\muldiv.div8.DU_Q1D1d11_EXT.fA.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.div8.DU_Q1D1d0.io_sel ),
    .SUM(\muldiv.div8.DU_Q1D1d12_EXT.fA.SUM ));
 sky130_fd_sc_hd__conb_1 \muldiv.div8.DU_Q1D1d12_EXT.fA.genblk1.fa_1_51  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(net51));
 sky130_fd_sc_hd__fa_2 \muldiv.div8.DU_Q1D1d2.fA.genblk1.fa_1  (.A(\muldiv.div8.DU_Q1D1d2.fA.A ),
    .B(net18),
    .CIN(\muldiv.div8.DU_Q1D1d1.fA.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.div8.DU_Q1D1d2.fA.COUT ),
    .SUM(\muldiv.div8.DU_Q1D1d2.fA.SUM ));
 sky130_fd_sc_hd__fa_2 \muldiv.div8.DU_Q1D1d3.fA.genblk1.fa_1  (.A(\muldiv.div8.DU_Q1D1d3.fA.A ),
    .B(net17),
    .CIN(\muldiv.div8.DU_Q1D1d2.fA.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.div8.DU_Q1D1d3.fA.COUT ),
    .SUM(\muldiv.div8.DU_Q1D1d3.fA.SUM ));
 sky130_fd_sc_hd__fa_2 \muldiv.div8.DU_Q1D1d4.fA.genblk1.fa_1  (.A(\muldiv.div8.DU_Q1D1d4.fA.A ),
    .B(net16),
    .CIN(\muldiv.div8.DU_Q1D1d3.fA.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.div8.DU_Q1D1d4.fA.COUT ),
    .SUM(\muldiv.div8.DU_Q1D1d4.fA.SUM ));
 sky130_fd_sc_hd__fa_2 \muldiv.div8.DU_Q1D1d5.fA.genblk1.fa_1  (.A(\muldiv.div8.DU_Q1D1d5.fA.A ),
    .B(net15),
    .CIN(\muldiv.div8.DU_Q1D1d4.fA.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.div8.DU_Q1D1d5.fA.COUT ),
    .SUM(\muldiv.div8.DU_Q1D1d5.fA.SUM ));
 sky130_fd_sc_hd__fa_2 \muldiv.div8.DU_Q1D1d6.fA.genblk1.fa_1  (.A(\muldiv.div8.DU_Q1D1d6.fA.A ),
    .B(net14),
    .CIN(\muldiv.div8.DU_Q1D1d5.fA.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.div8.DU_Q1D1d6.fA.COUT ),
    .SUM(\muldiv.div8.DU_Q1D1d6.fA.SUM ));
 sky130_fd_sc_hd__fa_2 \muldiv.div8.DU_Q1D1d7.fA.genblk1.fa_1  (.A(\muldiv.div8.DU_Q1D1d7.fA.A ),
    .B(\muldiv.div8.DU_Q0D0d7.fA.B ),
    .CIN(\muldiv.div8.DU_Q1D1d6.fA.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.div8.DU_Q1D1d7.fA.COUT ),
    .SUM(\muldiv.div8.DU_Q1D1d7.fA.SUM ));
 sky130_fd_sc_hd__fa_2 \muldiv.div8.DU_Q1D1d8_EXT.fA.genblk1.fa_1  (.A(\muldiv.div8.DU_Q1D1d8_EXT.fA.A ),
    .B(net52),
    .CIN(\muldiv.div8.DU_Q1D1d7.fA.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.div8.DU_Q1D1d8_EXT.fA.COUT ),
    .SUM(\muldiv.div8.DU_Q1D1d8_EXT.fA.SUM ));
 sky130_fd_sc_hd__conb_1 \muldiv.div8.DU_Q1D1d8_EXT.fA.genblk1.fa_1_52  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(net52));
 sky130_fd_sc_hd__fa_2 \muldiv.div8.DU_Q1D1d9_EXT.fA.genblk1.fa_1  (.A(\muldiv.div8.DU_Q1D1d9_EXT.fA.A ),
    .B(net53),
    .CIN(\muldiv.div8.DU_Q1D1d8_EXT.fA.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.div8.DU_Q1D1d10_EXT.fA.CIN ),
    .SUM(\muldiv.div8.DU_Q1D1d9_EXT.fA.SUM ));
 sky130_fd_sc_hd__conb_1 \muldiv.div8.DU_Q1D1d9_EXT.fA.genblk1.fa_1_53  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(net53));
 sky130_fd_sc_hd__fa_1 \muldiv.div8.DU_Q2D2d0.fA.genblk1.fa_1  (.A(\muldiv.div8.DU_Q2D2d0.fA.A ),
    .B(\muldiv.div8.DU_Q0D0d0.fA.B ),
    .CIN(net22),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.div8.DU_Q2D2d0.fA.COUT ),
    .SUM(\muldiv.div8.DU_Q2D2d0.fA.SUM ));
 sky130_fd_sc_hd__fa_2 \muldiv.div8.DU_Q2D2d1.fA.genblk1.fa_1  (.A(\muldiv.div8.DU_Q2D2d1.fA.A ),
    .B(\muldiv.div8.DU_Q0D0d1.fA.B ),
    .CIN(\muldiv.div8.DU_Q2D2d0.fA.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.div8.DU_Q2D2d1.fA.COUT ),
    .SUM(\muldiv.div8.DU_Q2D2d1.fA.SUM ));
 sky130_fd_sc_hd__fa_2 \muldiv.div8.DU_Q2D2d10_EXT.fA.genblk1.fa_1  (.A(\muldiv.div8.DU_Q2D2d10_EXT.fA.A ),
    .B(net54),
    .CIN(\muldiv.div8.DU_Q2D2d10_EXT.fA.CIN ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.div8.DU_Q2D2d10_EXT.fA.COUT ),
    .SUM(\muldiv.div8.DU_Q2D2d10_EXT.fA.SUM ));
 sky130_fd_sc_hd__conb_1 \muldiv.div8.DU_Q2D2d10_EXT.fA.genblk1.fa_1_54  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(net54));
 sky130_fd_sc_hd__fa_2 \muldiv.div8.DU_Q2D2d11_EXT.fA.genblk1.fa_1  (.A(\muldiv.div8.DU_Q2D2d11_EXT.fA.A ),
    .B(net55),
    .CIN(\muldiv.div8.DU_Q2D2d10_EXT.fA.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.div8.DU_Q2D2d0.io_sel ),
    .SUM(\muldiv.div8.DU_Q2D2d11_EXT.fA.SUM ));
 sky130_fd_sc_hd__conb_1 \muldiv.div8.DU_Q2D2d11_EXT.fA.genblk1.fa_1_55  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(net55));
 sky130_fd_sc_hd__fa_2 \muldiv.div8.DU_Q2D2d2.fA.genblk1.fa_1  (.A(\muldiv.div8.DU_Q2D2d2.fA.A ),
    .B(net18),
    .CIN(\muldiv.div8.DU_Q2D2d1.fA.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.div8.DU_Q2D2d2.fA.COUT ),
    .SUM(\muldiv.div8.DU_Q2D2d2.fA.SUM ));
 sky130_fd_sc_hd__fa_2 \muldiv.div8.DU_Q2D2d3.fA.genblk1.fa_1  (.A(\muldiv.div8.DU_Q2D2d3.fA.A ),
    .B(net17),
    .CIN(\muldiv.div8.DU_Q2D2d2.fA.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.div8.DU_Q2D2d3.fA.COUT ),
    .SUM(\muldiv.div8.DU_Q2D2d3.fA.SUM ));
 sky130_fd_sc_hd__fa_2 \muldiv.div8.DU_Q2D2d4.fA.genblk1.fa_1  (.A(\muldiv.div8.DU_Q2D2d4.fA.A ),
    .B(net16),
    .CIN(\muldiv.div8.DU_Q2D2d3.fA.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.div8.DU_Q2D2d4.fA.COUT ),
    .SUM(\muldiv.div8.DU_Q2D2d4.fA.SUM ));
 sky130_fd_sc_hd__fa_2 \muldiv.div8.DU_Q2D2d5.fA.genblk1.fa_1  (.A(\muldiv.div8.DU_Q2D2d5.fA.A ),
    .B(net15),
    .CIN(\muldiv.div8.DU_Q2D2d4.fA.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.div8.DU_Q2D2d5.fA.COUT ),
    .SUM(\muldiv.div8.DU_Q2D2d5.fA.SUM ));
 sky130_fd_sc_hd__fa_2 \muldiv.div8.DU_Q2D2d6.fA.genblk1.fa_1  (.A(\muldiv.div8.DU_Q2D2d6.fA.A ),
    .B(net14),
    .CIN(\muldiv.div8.DU_Q2D2d5.fA.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.div8.DU_Q2D2d6.fA.COUT ),
    .SUM(\muldiv.div8.DU_Q2D2d6.fA.SUM ));
 sky130_fd_sc_hd__fa_2 \muldiv.div8.DU_Q2D2d7.fA.genblk1.fa_1  (.A(\muldiv.div8.DU_Q2D2d7.fA.A ),
    .B(\muldiv.div8.DU_Q0D0d7.fA.B ),
    .CIN(\muldiv.div8.DU_Q2D2d6.fA.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.div8.DU_Q2D2d7.fA.COUT ),
    .SUM(\muldiv.div8.DU_Q2D2d7.fA.SUM ));
 sky130_fd_sc_hd__fa_2 \muldiv.div8.DU_Q2D2d8_EXT.fA.genblk1.fa_1  (.A(\muldiv.div8.DU_Q2D2d8_EXT.fA.A ),
    .B(net56),
    .CIN(\muldiv.div8.DU_Q2D2d7.fA.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.div8.DU_Q2D2d8_EXT.fA.COUT ),
    .SUM(\muldiv.div8.DU_Q2D2d8_EXT.fA.SUM ));
 sky130_fd_sc_hd__conb_1 \muldiv.div8.DU_Q2D2d8_EXT.fA.genblk1.fa_1_56  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(net56));
 sky130_fd_sc_hd__fa_2 \muldiv.div8.DU_Q2D2d9_EXT.fA.genblk1.fa_1  (.A(\muldiv.div8.DU_Q2D2d9_EXT.fA.A ),
    .B(net57),
    .CIN(\muldiv.div8.DU_Q2D2d8_EXT.fA.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.div8.DU_Q2D2d10_EXT.fA.CIN ),
    .SUM(\muldiv.div8.DU_Q2D2d9_EXT.fA.SUM ));
 sky130_fd_sc_hd__conb_1 \muldiv.div8.DU_Q2D2d9_EXT.fA.genblk1.fa_1_57  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(net57));
 sky130_fd_sc_hd__fa_1 \muldiv.div8.DU_Q3D3d0.fA.genblk1.fa_1  (.A(\muldiv.div8.DU_Q3D3d0.fA.A ),
    .B(net20),
    .CIN(net22),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.div8.DU_Q3D3d0.fA.COUT ),
    .SUM(\muldiv.div8.DU_Q3D3d0.fA.SUM ));
 sky130_fd_sc_hd__fa_2 \muldiv.div8.DU_Q3D3d1.fA.genblk1.fa_1  (.A(\muldiv.div8.DU_Q3D3d1.fA.A ),
    .B(\muldiv.div8.DU_Q0D0d1.fA.B ),
    .CIN(\muldiv.div8.DU_Q3D3d0.fA.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.div8.DU_Q3D3d1.fA.COUT ),
    .SUM(\muldiv.div8.DU_Q3D3d1.fA.SUM ));
 sky130_fd_sc_hd__fa_2 \muldiv.div8.DU_Q3D3d10_EXT.fA.genblk1.fa_1  (.A(\muldiv.div8.DU_Q3D3d10_EXT.fA.A ),
    .B(net58),
    .CIN(\muldiv.div8.DU_Q3D3d10_EXT.fA.CIN ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.div8.DU_Q3D3d0.io_sel ),
    .SUM(\muldiv.div8.DU_Q3D3d10_EXT.fA.SUM ));
 sky130_fd_sc_hd__conb_1 \muldiv.div8.DU_Q3D3d10_EXT.fA.genblk1.fa_1_58  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(net58));
 sky130_fd_sc_hd__fa_2 \muldiv.div8.DU_Q3D3d2.fA.genblk1.fa_1  (.A(\muldiv.div8.DU_Q3D3d2.fA.A ),
    .B(net18),
    .CIN(\muldiv.div8.DU_Q3D3d1.fA.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.div8.DU_Q3D3d2.fA.COUT ),
    .SUM(\muldiv.div8.DU_Q3D3d2.fA.SUM ));
 sky130_fd_sc_hd__fa_2 \muldiv.div8.DU_Q3D3d3.fA.genblk1.fa_1  (.A(\muldiv.div8.DU_Q3D3d3.fA.A ),
    .B(net17),
    .CIN(\muldiv.div8.DU_Q3D3d2.fA.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.div8.DU_Q3D3d3.fA.COUT ),
    .SUM(\muldiv.div8.DU_Q3D3d3.fA.SUM ));
 sky130_fd_sc_hd__fa_2 \muldiv.div8.DU_Q3D3d4.fA.genblk1.fa_1  (.A(\muldiv.div8.DU_Q3D3d4.fA.A ),
    .B(net16),
    .CIN(\muldiv.div8.DU_Q3D3d3.fA.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.div8.DU_Q3D3d4.fA.COUT ),
    .SUM(\muldiv.div8.DU_Q3D3d4.fA.SUM ));
 sky130_fd_sc_hd__fa_2 \muldiv.div8.DU_Q3D3d5.fA.genblk1.fa_1  (.A(\muldiv.div8.DU_Q3D3d5.fA.A ),
    .B(net15),
    .CIN(\muldiv.div8.DU_Q3D3d4.fA.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.div8.DU_Q3D3d5.fA.COUT ),
    .SUM(\muldiv.div8.DU_Q3D3d5.fA.SUM ));
 sky130_fd_sc_hd__fa_2 \muldiv.div8.DU_Q3D3d6.fA.genblk1.fa_1  (.A(\muldiv.div8.DU_Q3D3d6.fA.A ),
    .B(net14),
    .CIN(\muldiv.div8.DU_Q3D3d5.fA.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.div8.DU_Q3D3d6.fA.COUT ),
    .SUM(\muldiv.div8.DU_Q3D3d6.fA.SUM ));
 sky130_fd_sc_hd__fa_2 \muldiv.div8.DU_Q3D3d7.fA.genblk1.fa_1  (.A(\muldiv.div8.DU_Q3D3d7.fA.A ),
    .B(\muldiv.div8.DU_Q0D0d7.fA.B ),
    .CIN(\muldiv.div8.DU_Q3D3d6.fA.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.div8.DU_Q3D3d7.fA.COUT ),
    .SUM(\muldiv.div8.DU_Q3D3d7.fA.SUM ));
 sky130_fd_sc_hd__fa_2 \muldiv.div8.DU_Q3D3d8_EXT.fA.genblk1.fa_1  (.A(\muldiv.div8.DU_Q3D3d8_EXT.fA.A ),
    .B(net59),
    .CIN(\muldiv.div8.DU_Q3D3d7.fA.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.div8.DU_Q3D3d8_EXT.fA.COUT ),
    .SUM(\muldiv.div8.DU_Q3D3d8_EXT.fA.SUM ));
 sky130_fd_sc_hd__conb_1 \muldiv.div8.DU_Q3D3d8_EXT.fA.genblk1.fa_1_59  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(net59));
 sky130_fd_sc_hd__fa_2 \muldiv.div8.DU_Q3D3d9_EXT.fA.genblk1.fa_1  (.A(\muldiv.div8.DU_Q3D3d9_EXT.fA.A ),
    .B(net60),
    .CIN(\muldiv.div8.DU_Q3D3d8_EXT.fA.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.div8.DU_Q3D3d10_EXT.fA.CIN ),
    .SUM(\muldiv.div8.DU_Q3D3d9_EXT.fA.SUM ));
 sky130_fd_sc_hd__conb_1 \muldiv.div8.DU_Q3D3d9_EXT.fA.genblk1.fa_1_60  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(net60));
 sky130_fd_sc_hd__fa_1 \muldiv.div8.DU_Q4D4d0.fA.genblk1.fa_1  (.A(\muldiv.div8.DU_Q4D4d0.fA.A ),
    .B(net20),
    .CIN(net21),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.div8.DU_Q4D4d0.fA.COUT ),
    .SUM(\muldiv.div8.DU_Q4D4d0.fA.SUM ));
 sky130_fd_sc_hd__fa_2 \muldiv.div8.DU_Q4D4d1.fA.genblk1.fa_1  (.A(\muldiv.div8.DU_Q4D4d1.fA.A ),
    .B(net19),
    .CIN(\muldiv.div8.DU_Q4D4d0.fA.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.div8.DU_Q4D4d1.fA.COUT ),
    .SUM(\muldiv.div8.DU_Q4D4d1.fA.SUM ));
 sky130_fd_sc_hd__fa_2 \muldiv.div8.DU_Q4D4d2.fA.genblk1.fa_1  (.A(\muldiv.div8.DU_Q4D4d2.fA.A ),
    .B(net18),
    .CIN(\muldiv.div8.DU_Q4D4d1.fA.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.div8.DU_Q4D4d2.fA.COUT ),
    .SUM(\muldiv.div8.DU_Q4D4d2.fA.SUM ));
 sky130_fd_sc_hd__fa_2 \muldiv.div8.DU_Q4D4d3.fA.genblk1.fa_1  (.A(\muldiv.div8.DU_Q4D4d3.fA.A ),
    .B(net17),
    .CIN(\muldiv.div8.DU_Q4D4d2.fA.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.div8.DU_Q4D4d3.fA.COUT ),
    .SUM(\muldiv.div8.DU_Q4D4d3.fA.SUM ));
 sky130_fd_sc_hd__fa_2 \muldiv.div8.DU_Q4D4d4.fA.genblk1.fa_1  (.A(\muldiv.div8.DU_Q4D4d4.fA.A ),
    .B(net16),
    .CIN(\muldiv.div8.DU_Q4D4d3.fA.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.div8.DU_Q4D4d4.fA.COUT ),
    .SUM(\muldiv.div8.DU_Q4D4d4.fA.SUM ));
 sky130_fd_sc_hd__fa_2 \muldiv.div8.DU_Q4D4d5.fA.genblk1.fa_1  (.A(\muldiv.div8.DU_Q4D4d5.fA.A ),
    .B(net15),
    .CIN(\muldiv.div8.DU_Q4D4d4.fA.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.div8.DU_Q4D4d5.fA.COUT ),
    .SUM(\muldiv.div8.DU_Q4D4d5.fA.SUM ));
 sky130_fd_sc_hd__fa_2 \muldiv.div8.DU_Q4D4d6.fA.genblk1.fa_1  (.A(\muldiv.div8.DU_Q4D4d6.fA.A ),
    .B(net14),
    .CIN(\muldiv.div8.DU_Q4D4d5.fA.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.div8.DU_Q4D4d6.fA.COUT ),
    .SUM(\muldiv.div8.DU_Q4D4d6.fA.SUM ));
 sky130_fd_sc_hd__fa_2 \muldiv.div8.DU_Q4D4d7.fA.genblk1.fa_1  (.A(\muldiv.div8.DU_Q4D4d7.fA.A ),
    .B(\muldiv.div8.DU_Q0D0d7.fA.B ),
    .CIN(\muldiv.div8.DU_Q4D4d6.fA.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.div8.DU_Q4D4d7.fA.COUT ),
    .SUM(\muldiv.div8.DU_Q4D4d7.fA.SUM ));
 sky130_fd_sc_hd__fa_2 \muldiv.div8.DU_Q4D4d8_EXT.fA.genblk1.fa_1  (.A(\muldiv.div8.DU_Q4D4d8_EXT.fA.A ),
    .B(net61),
    .CIN(\muldiv.div8.DU_Q4D4d7.fA.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.div8.DU_Q4D4d8_EXT.fA.COUT ),
    .SUM(\muldiv.div8.DU_Q4D4d8_EXT.fA.SUM ));
 sky130_fd_sc_hd__conb_1 \muldiv.div8.DU_Q4D4d8_EXT.fA.genblk1.fa_1_61  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(net61));
 sky130_fd_sc_hd__fa_2 \muldiv.div8.DU_Q4D4d9_EXT.fA.genblk1.fa_1  (.A(\muldiv.div8.DU_Q4D4d9_EXT.fA.A ),
    .B(net62),
    .CIN(\muldiv.div8.DU_Q4D4d8_EXT.fA.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.div8.DU_Q4D4d0.io_sel ),
    .SUM(\muldiv.div8.DU_Q4D4d9_EXT.fA.SUM ));
 sky130_fd_sc_hd__conb_1 \muldiv.div8.DU_Q4D4d9_EXT.fA.genblk1.fa_1_62  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(net62));
 sky130_fd_sc_hd__fa_1 \muldiv.div8.DU_Q5D5d0.fA.genblk1.fa_1  (.A(\muldiv.div8.DU_Q5D5d0.fA.A ),
    .B(net20),
    .CIN(net21),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.div8.DU_Q5D5d0.fA.COUT ),
    .SUM(\muldiv.div8.DU_Q5D5d0.fA.SUM ));
 sky130_fd_sc_hd__fa_2 \muldiv.div8.DU_Q5D5d1.fA.genblk1.fa_1  (.A(\muldiv.div8.DU_Q5D5d1.fA.A ),
    .B(net19),
    .CIN(\muldiv.div8.DU_Q5D5d0.fA.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.div8.DU_Q5D5d1.fA.COUT ),
    .SUM(\muldiv.div8.DU_Q5D5d1.fA.SUM ));
 sky130_fd_sc_hd__fa_2 \muldiv.div8.DU_Q5D5d2.fA.genblk1.fa_1  (.A(\muldiv.div8.DU_Q5D5d2.fA.A ),
    .B(\muldiv.div8.DU_Q0D0d2.fA.B ),
    .CIN(\muldiv.div8.DU_Q5D5d1.fA.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.div8.DU_Q5D5d2.fA.COUT ),
    .SUM(\muldiv.div8.DU_Q5D5d2.fA.SUM ));
 sky130_fd_sc_hd__fa_2 \muldiv.div8.DU_Q5D5d3.fA.genblk1.fa_1  (.A(\muldiv.div8.DU_Q5D5d3.fA.A ),
    .B(net17),
    .CIN(\muldiv.div8.DU_Q5D5d2.fA.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.div8.DU_Q5D5d3.fA.COUT ),
    .SUM(\muldiv.div8.DU_Q5D5d3.fA.SUM ));
 sky130_fd_sc_hd__fa_2 \muldiv.div8.DU_Q5D5d4.fA.genblk1.fa_1  (.A(\muldiv.div8.DU_Q5D5d4.fA.A ),
    .B(net16),
    .CIN(\muldiv.div8.DU_Q5D5d3.fA.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.div8.DU_Q5D5d4.fA.COUT ),
    .SUM(\muldiv.div8.DU_Q5D5d4.fA.SUM ));
 sky130_fd_sc_hd__fa_2 \muldiv.div8.DU_Q5D5d5.fA.genblk1.fa_1  (.A(\muldiv.div8.DU_Q5D5d5.fA.A ),
    .B(net15),
    .CIN(\muldiv.div8.DU_Q5D5d4.fA.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.div8.DU_Q5D5d5.fA.COUT ),
    .SUM(\muldiv.div8.DU_Q5D5d5.fA.SUM ));
 sky130_fd_sc_hd__fa_2 \muldiv.div8.DU_Q5D5d6.fA.genblk1.fa_1  (.A(\muldiv.div8.DU_Q5D5d6.fA.A ),
    .B(net14),
    .CIN(\muldiv.div8.DU_Q5D5d5.fA.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.div8.DU_Q5D5d6.fA.COUT ),
    .SUM(\muldiv.div8.DU_Q5D5d6.fA.SUM ));
 sky130_fd_sc_hd__fa_2 \muldiv.div8.DU_Q5D5d7.fA.genblk1.fa_1  (.A(\muldiv.div8.DU_Q5D5d7.fA.A ),
    .B(\muldiv.div8.DU_Q0D0d7.fA.B ),
    .CIN(\muldiv.div8.DU_Q5D5d6.fA.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.div8.DU_Q5D5d7.fA.COUT ),
    .SUM(\muldiv.div8.DU_Q5D5d7.fA.SUM ));
 sky130_fd_sc_hd__fa_2 \muldiv.div8.DU_Q5D5d8_EXT.fA.genblk1.fa_1  (.A(\muldiv.div8.DU_Q5D5d8_EXT.fA.A ),
    .B(net63),
    .CIN(\muldiv.div8.DU_Q5D5d7.fA.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.div8.DU_Q5D5d0.io_sel ),
    .SUM(\muldiv.div8.DU_Q5D5d8_EXT.fA.SUM ));
 sky130_fd_sc_hd__conb_1 \muldiv.div8.DU_Q5D5d8_EXT.fA.genblk1.fa_1_63  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(net63));
 sky130_fd_sc_hd__fa_1 \muldiv.div8.DU_Q6D6d0.fA.genblk1.fa_1  (.A(\muldiv.div8.DU_Q6D6d0.fA.A ),
    .B(net20),
    .CIN(net21),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.div8.DU_Q6D6d0.fA.COUT ),
    .SUM(\muldiv.div8.DU_Q6D6d0.fA.SUM ));
 sky130_fd_sc_hd__fa_2 \muldiv.div8.DU_Q6D6d1.fA.genblk1.fa_1  (.A(\muldiv.div8.DU_Q6D6d1.fA.A ),
    .B(net19),
    .CIN(\muldiv.div8.DU_Q6D6d0.fA.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.div8.DU_Q6D6d1.fA.COUT ),
    .SUM(\muldiv.div8.DU_Q6D6d1.fA.SUM ));
 sky130_fd_sc_hd__fa_2 \muldiv.div8.DU_Q6D6d2.fA.genblk1.fa_1  (.A(\muldiv.div8.DU_Q6D6d2.fA.A ),
    .B(\muldiv.div8.DU_Q0D0d2.fA.B ),
    .CIN(\muldiv.div8.DU_Q6D6d1.fA.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.div8.DU_Q6D6d2.fA.COUT ),
    .SUM(\muldiv.div8.DU_Q6D6d2.fA.SUM ));
 sky130_fd_sc_hd__fa_2 \muldiv.div8.DU_Q6D6d3.fA.genblk1.fa_1  (.A(\muldiv.div8.DU_Q6D6d3.fA.A ),
    .B(\muldiv.div8.DU_Q0D0d3.fA.B ),
    .CIN(\muldiv.div8.DU_Q6D6d2.fA.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.div8.DU_Q6D6d3.fA.COUT ),
    .SUM(\muldiv.div8.DU_Q6D6d3.fA.SUM ));
 sky130_fd_sc_hd__fa_2 \muldiv.div8.DU_Q6D6d4.fA.genblk1.fa_1  (.A(\muldiv.div8.DU_Q6D6d4.fA.A ),
    .B(\muldiv.div8.DU_Q0D0d4.fA.B ),
    .CIN(\muldiv.div8.DU_Q6D6d3.fA.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.div8.DU_Q6D6d4.fA.COUT ),
    .SUM(\muldiv.div8.DU_Q6D6d4.fA.SUM ));
 sky130_fd_sc_hd__fa_2 \muldiv.div8.DU_Q6D6d5.fA.genblk1.fa_1  (.A(\muldiv.div8.DU_Q6D6d5.fA.A ),
    .B(\muldiv.div8.DU_Q0D0d5.fA.B ),
    .CIN(\muldiv.div8.DU_Q6D6d4.fA.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.div8.DU_Q6D6d5.fA.COUT ),
    .SUM(\muldiv.div8.DU_Q6D6d5.fA.SUM ));
 sky130_fd_sc_hd__fa_2 \muldiv.div8.DU_Q6D6d6.fA.genblk1.fa_1  (.A(\muldiv.div8.DU_Q6D6d6.fA.A ),
    .B(\muldiv.div8.DU_Q0D0d6.fA.B ),
    .CIN(\muldiv.div8.DU_Q6D6d5.fA.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.div8.DU_Q6D6d6.fA.COUT ),
    .SUM(\muldiv.div8.DU_Q6D6d6.fA.SUM ));
 sky130_fd_sc_hd__fa_2 \muldiv.div8.DU_Q6D6d7.fA.genblk1.fa_1  (.A(\muldiv.div8.DU_Q6D6d7.fA.A ),
    .B(\muldiv.div8.DU_Q0D0d7.fA.B ),
    .CIN(\muldiv.div8.DU_Q6D6d6.fA.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.div8.DU_Q6D6d0.io_sel ),
    .SUM(\muldiv.div8.DU_Q6D6d7.fA.SUM ));
 sky130_fd_sc_hd__fa_2 \muldiv.div8.DU_Q7D7d0.fA.genblk1.fa_1  (.A(\muldiv.div8.DU_Q7D7d0.fA.A ),
    .B(net20),
    .CIN(net21),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.div8.DU_Q7D7d0.fA.COUT ),
    .SUM(\muldiv.div8.DU_Q7D7d0.fA.SUM ));
 sky130_fd_sc_hd__fa_2 \muldiv.div8.DU_Q7D7d1.fA.genblk1.fa_1  (.A(net25),
    .B(net19),
    .CIN(\muldiv.div8.DU_Q7D7d0.fA.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.div8.DU_Q7D7d1.fA.COUT ),
    .SUM(\muldiv.div8.DU_Q7D7d1.fA.SUM ));
 sky130_fd_sc_hd__conb_1 \muldiv.div8.DU_Q7D7d1.fA.genblk1.fa_1_25  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net25));
 sky130_fd_sc_hd__fa_2 \muldiv.div8.DU_Q7D7d2.fA.genblk1.fa_1  (.A(net26),
    .B(\muldiv.div8.DU_Q0D0d2.fA.B ),
    .CIN(\muldiv.div8.DU_Q7D7d1.fA.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.div8.DU_Q7D7d2.fA.COUT ),
    .SUM(\muldiv.div8.DU_Q7D7d2.fA.SUM ));
 sky130_fd_sc_hd__conb_1 \muldiv.div8.DU_Q7D7d2.fA.genblk1.fa_1_26  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net26));
 sky130_fd_sc_hd__fa_2 \muldiv.div8.DU_Q7D7d3.fA.genblk1.fa_1  (.A(net27),
    .B(\muldiv.div8.DU_Q0D0d3.fA.B ),
    .CIN(\muldiv.div8.DU_Q7D7d2.fA.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.div8.DU_Q7D7d3.fA.COUT ),
    .SUM(\muldiv.div8.DU_Q7D7d3.fA.SUM ));
 sky130_fd_sc_hd__conb_1 \muldiv.div8.DU_Q7D7d3.fA.genblk1.fa_1_27  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net27));
 sky130_fd_sc_hd__fa_2 \muldiv.div8.DU_Q7D7d4.fA.genblk1.fa_1  (.A(net28),
    .B(\muldiv.div8.DU_Q0D0d4.fA.B ),
    .CIN(\muldiv.div8.DU_Q7D7d3.fA.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.div8.DU_Q7D7d4.fA.COUT ),
    .SUM(\muldiv.div8.DU_Q7D7d4.fA.SUM ));
 sky130_fd_sc_hd__conb_1 \muldiv.div8.DU_Q7D7d4.fA.genblk1.fa_1_28  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net28));
 sky130_fd_sc_hd__fa_2 \muldiv.div8.DU_Q7D7d5.fA.genblk1.fa_1  (.A(net29),
    .B(\muldiv.div8.DU_Q0D0d5.fA.B ),
    .CIN(\muldiv.div8.DU_Q7D7d4.fA.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.div8.DU_Q7D7d5.fA.COUT ),
    .SUM(\muldiv.div8.DU_Q7D7d5.fA.SUM ));
 sky130_fd_sc_hd__conb_1 \muldiv.div8.DU_Q7D7d5.fA.genblk1.fa_1_29  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net29));
 sky130_fd_sc_hd__fa_2 \muldiv.div8.DU_Q7D7d6.fA.genblk1.fa_1  (.A(net30),
    .B(\muldiv.div8.DU_Q0D0d6.fA.B ),
    .CIN(\muldiv.div8.DU_Q7D7d5.fA.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.div8.DU_Q7D7d6.fA.COUT ),
    .SUM(\muldiv.div8.DU_Q7D7d6.fA.SUM ));
 sky130_fd_sc_hd__conb_1 \muldiv.div8.DU_Q7D7d6.fA.genblk1.fa_1_30  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net30));
 sky130_fd_sc_hd__fa_2 \muldiv.div8.DU_Q7D7d7.fA.genblk1.fa_1  (.A(net31),
    .B(\muldiv.div8.DU_Q0D0d7.fA.B ),
    .CIN(\muldiv.div8.DU_Q7D7d6.fA.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.div8.DU_Q7D7d0.io_sel ),
    .SUM(\muldiv.div8.DU_Q7D7d7.fA.SUM ));
 sky130_fd_sc_hd__conb_1 \muldiv.div8.DU_Q7D7d7.fA.genblk1.fa_1_31  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net31));
 sky130_fd_sc_hd__ha_2 \muldiv.div8.HAD_DVD_TWOS_0.genblk1.ha_1  (.A(\muldiv.div8.HAD_DVD_TWOS_0.A ),
    .B(\muldiv.div8.HAD_DVD_TWOS_0.B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.div8.HAD_DVD_TWOS_0.COUT ),
    .SUM(\muldiv.div8.DU_Q0D0d0.fA.A ));
 sky130_fd_sc_hd__ha_4 \muldiv.div8.HAD_DVD_TWOS_1.genblk1.ha_1  (.A(\muldiv.div8.HAD_DVD_TWOS_1.A ),
    .B(\muldiv.div8.HAD_DVD_TWOS_0.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.div8.HAD_DVD_TWOS_1.COUT ),
    .SUM(\muldiv.div8.DU_Q1D1d0.fA.A ));
 sky130_fd_sc_hd__ha_4 \muldiv.div8.HAD_DVD_TWOS_2.genblk1.ha_1  (.A(\muldiv.div8.HAD_DVD_TWOS_2.A ),
    .B(\muldiv.div8.HAD_DVD_TWOS_1.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.div8.HAD_DVD_TWOS_2.COUT ),
    .SUM(\muldiv.div8.DU_Q2D2d0.fA.A ));
 sky130_fd_sc_hd__ha_4 \muldiv.div8.HAD_DVD_TWOS_3.genblk1.ha_1  (.A(\muldiv.div8.HAD_DVD_TWOS_3.A ),
    .B(\muldiv.div8.HAD_DVD_TWOS_2.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.div8.HAD_DVD_TWOS_3.COUT ),
    .SUM(\muldiv.div8.DU_Q3D3d0.fA.A ));
 sky130_fd_sc_hd__ha_4 \muldiv.div8.HAD_DVD_TWOS_4.genblk1.ha_1  (.A(\muldiv.div8.HAD_DVD_TWOS_4.A ),
    .B(\muldiv.div8.HAD_DVD_TWOS_3.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.div8.HAD_DVD_TWOS_4.COUT ),
    .SUM(\muldiv.div8.DU_Q4D4d0.fA.A ));
 sky130_fd_sc_hd__ha_4 \muldiv.div8.HAD_DVD_TWOS_5.genblk1.ha_1  (.A(\muldiv.div8.HAD_DVD_TWOS_5.A ),
    .B(\muldiv.div8.HAD_DVD_TWOS_4.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.div8.HAD_DVD_TWOS_5.COUT ),
    .SUM(\muldiv.div8.DU_Q5D5d0.fA.A ));
 sky130_fd_sc_hd__ha_4 \muldiv.div8.HAD_DVD_TWOS_6.genblk1.ha_1  (.A(\muldiv.div8.HAD_DVD_TWOS_6.A ),
    .B(\muldiv.div8.HAD_DVD_TWOS_5.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.div8.HAD_DVD_TWOS_6.COUT ),
    .SUM(\muldiv.div8.DU_Q6D6d0.fA.A ));
 sky130_fd_sc_hd__ha_4 \muldiv.div8.HAD_DVD_TWOS_7.genblk1.ha_1  (.A(\muldiv.div8.HAD_DVD_TWOS_7.A ),
    .B(\muldiv.div8.HAD_DVD_TWOS_6.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.div8.HAD_DVD_TWOS_7.COUT ),
    .SUM(\muldiv.div8.DU_Q7D7d0.fA.A ));
 sky130_fd_sc_hd__ha_2 \muldiv.div8.HAQ0_SIGN.genblk1.ha_1  (.A(\muldiv.div8.HAQ0_SIGN.A ),
    .B(\muldiv.div8.HAQ0_SIGN.B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.div8.HAQ0_SIGN.COUT ),
    .SUM(\muldiv.div8.HAQ0_SIGN.SUM ));
 sky130_fd_sc_hd__ha_1 \muldiv.div8.HAQ1_SIGN.genblk1.ha_1  (.A(\muldiv.div8.HAQ1_SIGN.A ),
    .B(\muldiv.div8.HAQ0_SIGN.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.div8.HAQ1_SIGN.COUT ),
    .SUM(\muldiv.div8.HAQ1_SIGN.SUM ));
 sky130_fd_sc_hd__ha_1 \muldiv.div8.HAQ2_SIGN.genblk1.ha_1  (.A(\muldiv.div8.HAQ2_SIGN.A ),
    .B(\muldiv.div8.HAQ1_SIGN.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.div8.HAQ2_SIGN.COUT ),
    .SUM(\muldiv.div8.HAQ2_SIGN.SUM ));
 sky130_fd_sc_hd__ha_1 \muldiv.div8.HAQ3_SIGN.genblk1.ha_1  (.A(\muldiv.div8.HAQ3_SIGN.A ),
    .B(\muldiv.div8.HAQ2_SIGN.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.div8.HAQ3_SIGN.COUT ),
    .SUM(\muldiv.div8.HAQ3_SIGN.SUM ));
 sky130_fd_sc_hd__ha_1 \muldiv.div8.HAQ4_SIGN.genblk1.ha_1  (.A(\muldiv.div8.HAQ4_SIGN.A ),
    .B(\muldiv.div8.HAQ3_SIGN.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.div8.HAQ4_SIGN.COUT ),
    .SUM(\muldiv.div8.HAQ4_SIGN.SUM ));
 sky130_fd_sc_hd__ha_2 \muldiv.div8.HAQ5_SIGN.genblk1.ha_1  (.A(\muldiv.div8.HAQ5_SIGN.A ),
    .B(\muldiv.div8.HAQ4_SIGN.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.div8.HAQ5_SIGN.COUT ),
    .SUM(\muldiv.div8.HAQ5_SIGN.SUM ));
 sky130_fd_sc_hd__ha_2 \muldiv.div8.HAQ6_SIGN.genblk1.ha_1  (.A(\muldiv.div8.HAQ6_SIGN.A ),
    .B(\muldiv.div8.HAQ5_SIGN.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.div8.HAQ6_SIGN.COUT ),
    .SUM(\muldiv.div8.HAQ6_SIGN.SUM ));
 sky130_fd_sc_hd__ha_2 \muldiv.div8.HAQ7_SIGN.genblk1.ha_1  (.A(\muldiv.div8.HAQ7_SIGN.A ),
    .B(\muldiv.div8.HAQ6_SIGN.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.div8.HAQ7_SIGN.COUT ),
    .SUM(\muldiv.div8.HAQ7_SIGN.SUM ));
 sky130_fd_sc_hd__ha_2 \muldiv.div8.HAR0_SIGN.genblk1.ha_1  (.A(\muldiv.div8.HAR0_SIGN.A ),
    .B(\muldiv.div8.HAD_DVD_TWOS_0.B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.div8.HAR0_SIGN.COUT ),
    .SUM(\muldiv.div8.HAR0_SIGN.SUM ));
 sky130_fd_sc_hd__ha_4 \muldiv.div8.HAR1_SIGN.genblk1.ha_1  (.A(\muldiv.div8.HAR1_SIGN.A ),
    .B(\muldiv.div8.HAR0_SIGN.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.div8.HAR1_SIGN.COUT ),
    .SUM(\muldiv.div8.HAR1_SIGN.SUM ));
 sky130_fd_sc_hd__ha_4 \muldiv.div8.HAR2_SIGN.genblk1.ha_1  (.A(\muldiv.div8.HAR2_SIGN.A ),
    .B(\muldiv.div8.HAR1_SIGN.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.div8.HAR2_SIGN.COUT ),
    .SUM(\muldiv.div8.HAR2_SIGN.SUM ));
 sky130_fd_sc_hd__ha_4 \muldiv.div8.HAR3_SIGN.genblk1.ha_1  (.A(\muldiv.div8.HAR3_SIGN.A ),
    .B(\muldiv.div8.HAR2_SIGN.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.div8.HAR3_SIGN.COUT ),
    .SUM(\muldiv.div8.HAR3_SIGN.SUM ));
 sky130_fd_sc_hd__ha_4 \muldiv.div8.HAR4_SIGN.genblk1.ha_1  (.A(\muldiv.div8.HAR4_SIGN.A ),
    .B(\muldiv.div8.HAR3_SIGN.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.div8.HAR4_SIGN.COUT ),
    .SUM(\muldiv.div8.HAR4_SIGN.SUM ));
 sky130_fd_sc_hd__ha_4 \muldiv.div8.HAR5_SIGN.genblk1.ha_1  (.A(\muldiv.div8.HAR5_SIGN.A ),
    .B(\muldiv.div8.HAR4_SIGN.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.div8.HAR5_SIGN.COUT ),
    .SUM(\muldiv.div8.HAR5_SIGN.SUM ));
 sky130_fd_sc_hd__ha_4 \muldiv.div8.HAR6_SIGN.genblk1.ha_1  (.A(\muldiv.div8.HAR6_SIGN.A ),
    .B(\muldiv.div8.HAR5_SIGN.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.div8.HAR6_SIGN.COUT ),
    .SUM(\muldiv.div8.HAR6_SIGN.SUM ));
 sky130_fd_sc_hd__ha_4 \muldiv.div8.HAR7_SIGN.genblk1.ha_1  (.A(\muldiv.div8.HAR7_SIGN.A ),
    .B(\muldiv.div8.HAR6_SIGN.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.div8.HAR7_SIGN.COUT ),
    .SUM(\muldiv.div8.HAR7_SIGN.SUM ));
 sky130_fd_sc_hd__fa_1 \muldiv.mul8.FA_P10A3B7.genblk1.fa_1  (.A(\muldiv.mul8.FA_P10A3B7.A ),
    .B(\muldiv.mul8.FA_P10A3B7.B ),
    .CIN(\muldiv.mul8.FA_P10A3B7.CIN ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.mul8.FA_P10A3B7.COUT ),
    .SUM(\muldiv.mul8.FA_P10A3B7.SUM ));
 sky130_fd_sc_hd__fa_1 \muldiv.mul8.FA_P10A4B6.genblk1.fa_1  (.A(\muldiv.mul8.FA_P10A4B6.A ),
    .B(\muldiv.mul8.A4xB6_52 ),
    .CIN(\muldiv.mul8.FA_P10A4B6.CIN ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.mul8.FA_P10A4B6.COUT ),
    .SUM(\muldiv.mul8.FA_P10A3B7.A ));
 sky130_fd_sc_hd__fa_1 \muldiv.mul8.FA_P10A5B5.genblk1.fa_1  (.A(\muldiv.mul8.FA_P10A5B5.A ),
    .B(\muldiv.mul8.A5xB5_45 ),
    .CIN(\muldiv.mul8.FA_P10A5B5.CIN ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.mul8.FA_P10A5B5.COUT ),
    .SUM(\muldiv.mul8.FA_P10A4B6.A ));
 sky130_fd_sc_hd__fa_1 \muldiv.mul8.FA_P10A6B4.genblk1.fa_1  (.A(\muldiv.mul8.FA_P10A6B4.A ),
    .B(\muldiv.mul8.A6xB4_38 ),
    .CIN(\muldiv.mul8.FA_P10A6B4.CIN ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.mul8.FA_P10A6B4.COUT ),
    .SUM(\muldiv.mul8.FA_P10A5B5.A ));
 sky130_fd_sc_hd__fa_1 \muldiv.mul8.FA_P10A7B1.genblk1.fa_1  (.A(\muldiv.mul8.FA_P10A7B1.A ),
    .B(\muldiv.mul8.FA_P10A7B1.B ),
    .CIN(\muldiv.mul8.FA_P10A7B1.CIN ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.mul8.FA_P10A7B1.COUT ),
    .SUM(\muldiv.mul8.FA_P10A7B1.SUM ));
 sky130_fd_sc_hd__fa_1 \muldiv.mul8.FA_P10A7B2.genblk1.fa_1  (.A(\muldiv.mul8.FA_P10A7B1.SUM ),
    .B(\muldiv.mul8.FA_P10A7B2.B ),
    .CIN(\muldiv.mul8.FA_P10A7B2.CIN ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.mul8.FA_P10A7B2.COUT ),
    .SUM(\muldiv.mul8.FA_P10A7B2.SUM ));
 sky130_fd_sc_hd__fa_1 \muldiv.mul8.FA_P10A7B3.genblk1.fa_1  (.A(\muldiv.mul8.FA_P10A7B2.SUM ),
    .B(\muldiv.mul8.A7xB3_31 ),
    .CIN(\muldiv.mul8.FA_P10A7B3.CIN ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.mul8.FA_P10A7B3.COUT ),
    .SUM(\muldiv.mul8.FA_P10A6B4.A ));
 sky130_fd_sc_hd__fa_1 \muldiv.mul8.FA_P11A4B7.genblk1.fa_1  (.A(\muldiv.mul8.FA_P11A4B7.A ),
    .B(\muldiv.mul8.FA_P11A4B7.B ),
    .CIN(\muldiv.mul8.FA_P10A3B7.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.mul8.FA_P11A4B7.COUT ),
    .SUM(\muldiv.mul8.FA_P11A4B7.SUM ));
 sky130_fd_sc_hd__fa_1 \muldiv.mul8.FA_P11A5B6.genblk1.fa_1  (.A(\muldiv.mul8.FA_P11A5B6.A ),
    .B(\muldiv.mul8.A5xB6_53 ),
    .CIN(\muldiv.mul8.FA_P10A4B6.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.mul8.FA_P11A5B6.COUT ),
    .SUM(\muldiv.mul8.FA_P11A4B7.A ));
 sky130_fd_sc_hd__fa_1 \muldiv.mul8.FA_P11A6B5.genblk1.fa_1  (.A(\muldiv.mul8.FA_P11A6B5.A ),
    .B(\muldiv.mul8.A6xB5_46 ),
    .CIN(\muldiv.mul8.FA_P10A5B5.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.mul8.FA_P11A6B5.COUT ),
    .SUM(\muldiv.mul8.FA_P11A5B6.A ));
 sky130_fd_sc_hd__fa_1 \muldiv.mul8.FA_P11A7B1.genblk1.fa_1  (.A(\muldiv.mul8.FA_P10A7B1.A ),
    .B(\muldiv.mul8.FA_P10A7B1.B ),
    .CIN(\muldiv.mul8.FA_P10A7B1.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.mul8.FA_P11A7B1.COUT ),
    .SUM(\muldiv.mul8.FA_P11A7B1.SUM ));
 sky130_fd_sc_hd__fa_1 \muldiv.mul8.FA_P11A7B2.genblk1.fa_1  (.A(\muldiv.mul8.FA_P11A7B1.SUM ),
    .B(\muldiv.mul8.FA_P10A7B2.B ),
    .CIN(\muldiv.mul8.FA_P10A7B2.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.mul8.FA_P11A7B2.COUT ),
    .SUM(\muldiv.mul8.FA_P11A7B2.SUM ));
 sky130_fd_sc_hd__fa_1 \muldiv.mul8.FA_P11A7B3.genblk1.fa_1  (.A(\muldiv.mul8.FA_P11A7B2.SUM ),
    .B(\muldiv.mul8.FA_P11A7B3.B ),
    .CIN(\muldiv.mul8.FA_P10A7B3.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.mul8.FA_P11A7B3.COUT ),
    .SUM(\muldiv.mul8.FA_P11A7B3.SUM ));
 sky130_fd_sc_hd__fa_1 \muldiv.mul8.FA_P11A7B4.genblk1.fa_1  (.A(\muldiv.mul8.FA_P11A7B3.SUM ),
    .B(\muldiv.mul8.A7xB4_39 ),
    .CIN(\muldiv.mul8.FA_P10A6B4.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.mul8.FA_P11A7B4.COUT ),
    .SUM(\muldiv.mul8.FA_P11A6B5.A ));
 sky130_fd_sc_hd__fa_1 \muldiv.mul8.FA_P12A5B7.genblk1.fa_1  (.A(\muldiv.mul8.FA_P12A5B7.A ),
    .B(\muldiv.mul8.FA_P12A5B7.B ),
    .CIN(\muldiv.mul8.FA_P11A4B7.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.mul8.FA_P12A5B7.COUT ),
    .SUM(\muldiv.mul8.FA_P12A5B7.SUM ));
 sky130_fd_sc_hd__fa_1 \muldiv.mul8.FA_P12A6B6.genblk1.fa_1  (.A(\muldiv.mul8.FA_P12A6B6.A ),
    .B(\muldiv.mul8.A6xB6_54 ),
    .CIN(\muldiv.mul8.FA_P11A5B6.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.mul8.FA_P12A6B6.COUT ),
    .SUM(\muldiv.mul8.FA_P12A5B7.A ));
 sky130_fd_sc_hd__fa_1 \muldiv.mul8.FA_P12A7B1.genblk1.fa_1  (.A(\muldiv.mul8.FA_P10A7B1.A ),
    .B(\muldiv.mul8.FA_P10A7B1.B ),
    .CIN(\muldiv.mul8.FA_P11A7B1.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.mul8.FA_P12A7B1.COUT ),
    .SUM(\muldiv.mul8.FA_P12A7B1.SUM ));
 sky130_fd_sc_hd__fa_1 \muldiv.mul8.FA_P12A7B2.genblk1.fa_1  (.A(\muldiv.mul8.FA_P12A7B1.SUM ),
    .B(\muldiv.mul8.FA_P10A7B2.B ),
    .CIN(\muldiv.mul8.FA_P11A7B2.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.mul8.FA_P12A7B2.COUT ),
    .SUM(\muldiv.mul8.FA_P12A7B2.SUM ));
 sky130_fd_sc_hd__fa_1 \muldiv.mul8.FA_P12A7B3.genblk1.fa_1  (.A(\muldiv.mul8.FA_P12A7B2.SUM ),
    .B(\muldiv.mul8.FA_P11A7B3.B ),
    .CIN(\muldiv.mul8.FA_P11A7B3.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.mul8.FA_P12A7B3.COUT ),
    .SUM(\muldiv.mul8.FA_P12A7B3.SUM ));
 sky130_fd_sc_hd__fa_1 \muldiv.mul8.FA_P12A7B4.genblk1.fa_1  (.A(\muldiv.mul8.FA_P12A7B3.SUM ),
    .B(\muldiv.mul8.FA_P12A7B4.B ),
    .CIN(\muldiv.mul8.FA_P11A7B4.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.mul8.FA_P12A7B4.COUT ),
    .SUM(\muldiv.mul8.FA_P12A7B4.SUM ));
 sky130_fd_sc_hd__fa_1 \muldiv.mul8.FA_P12A7B5.genblk1.fa_1  (.A(\muldiv.mul8.FA_P12A7B4.SUM ),
    .B(\muldiv.mul8.A7xB5_47 ),
    .CIN(\muldiv.mul8.FA_P11A6B5.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.mul8.FA_P12A7B5.COUT ),
    .SUM(\muldiv.mul8.FA_P12A6B6.A ));
 sky130_fd_sc_hd__fa_1 \muldiv.mul8.FA_P13A6B7.genblk1.fa_1  (.A(\muldiv.mul8.FA_P13A6B7.A ),
    .B(\muldiv.mul8.FA_P13A6B7.B ),
    .CIN(\muldiv.mul8.FA_P12A5B7.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.mul8.FA_P13A6B7.COUT ),
    .SUM(\muldiv.mul8.FA_P13A6B7.SUM ));
 sky130_fd_sc_hd__fa_1 \muldiv.mul8.FA_P13A7B1.genblk1.fa_1  (.A(\muldiv.mul8.FA_P10A7B1.A ),
    .B(\muldiv.mul8.FA_P10A7B1.B ),
    .CIN(\muldiv.mul8.FA_P12A7B1.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.mul8.FA_P13A7B1.COUT ),
    .SUM(\muldiv.mul8.FA_P13A7B1.SUM ));
 sky130_fd_sc_hd__fa_1 \muldiv.mul8.FA_P13A7B2.genblk1.fa_1  (.A(\muldiv.mul8.FA_P13A7B1.SUM ),
    .B(\muldiv.mul8.FA_P10A7B2.B ),
    .CIN(\muldiv.mul8.FA_P12A7B2.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.mul8.FA_P13A7B2.COUT ),
    .SUM(\muldiv.mul8.FA_P13A7B2.SUM ));
 sky130_fd_sc_hd__fa_1 \muldiv.mul8.FA_P13A7B3.genblk1.fa_1  (.A(\muldiv.mul8.FA_P13A7B2.SUM ),
    .B(\muldiv.mul8.FA_P11A7B3.B ),
    .CIN(\muldiv.mul8.FA_P12A7B3.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.mul8.FA_P13A7B3.COUT ),
    .SUM(\muldiv.mul8.FA_P13A7B3.SUM ));
 sky130_fd_sc_hd__fa_1 \muldiv.mul8.FA_P13A7B4.genblk1.fa_1  (.A(\muldiv.mul8.FA_P13A7B3.SUM ),
    .B(\muldiv.mul8.FA_P12A7B4.B ),
    .CIN(\muldiv.mul8.FA_P12A7B4.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.mul8.FA_P13A7B4.COUT ),
    .SUM(\muldiv.mul8.FA_P13A7B4.SUM ));
 sky130_fd_sc_hd__fa_1 \muldiv.mul8.FA_P13A7B5.genblk1.fa_1  (.A(\muldiv.mul8.FA_P13A7B4.SUM ),
    .B(\muldiv.mul8.FA_P13A7B5.B ),
    .CIN(\muldiv.mul8.FA_P12A7B5.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.mul8.FA_P13A7B5.COUT ),
    .SUM(\muldiv.mul8.FA_P13A7B5.SUM ));
 sky130_fd_sc_hd__fa_1 \muldiv.mul8.FA_P13A7B6.genblk1.fa_1  (.A(\muldiv.mul8.FA_P13A7B5.SUM ),
    .B(\muldiv.mul8.A7xB6_55 ),
    .CIN(\muldiv.mul8.FA_P12A6B6.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.mul8.FA_P13A7B6.COUT ),
    .SUM(\muldiv.mul8.FA_P13A6B7.A ));
 sky130_fd_sc_hd__fa_1 \muldiv.mul8.FA_P14A7B1.genblk1.fa_1  (.A(\muldiv.mul8.FA_P10A7B1.A ),
    .B(\muldiv.mul8.FA_P10A7B1.B ),
    .CIN(\muldiv.mul8.FA_P13A7B1.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.mul8.FA_P14A7B1.COUT ),
    .SUM(\muldiv.mul8.FA_P14A7B1.SUM ));
 sky130_fd_sc_hd__fa_1 \muldiv.mul8.FA_P14A7B2.genblk1.fa_1  (.A(\muldiv.mul8.FA_P14A7B1.SUM ),
    .B(\muldiv.mul8.FA_P10A7B2.B ),
    .CIN(\muldiv.mul8.FA_P13A7B2.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.mul8.FA_P14A7B2.COUT ),
    .SUM(\muldiv.mul8.FA_P14A7B2.SUM ));
 sky130_fd_sc_hd__fa_1 \muldiv.mul8.FA_P14A7B3.genblk1.fa_1  (.A(\muldiv.mul8.FA_P14A7B2.SUM ),
    .B(\muldiv.mul8.FA_P11A7B3.B ),
    .CIN(\muldiv.mul8.FA_P13A7B3.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.mul8.FA_P14A7B3.COUT ),
    .SUM(\muldiv.mul8.FA_P14A7B3.SUM ));
 sky130_fd_sc_hd__fa_1 \muldiv.mul8.FA_P14A7B4.genblk1.fa_1  (.A(\muldiv.mul8.FA_P14A7B3.SUM ),
    .B(\muldiv.mul8.FA_P12A7B4.B ),
    .CIN(\muldiv.mul8.FA_P13A7B4.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.mul8.FA_P14A7B4.COUT ),
    .SUM(\muldiv.mul8.FA_P14A7B4.SUM ));
 sky130_fd_sc_hd__fa_1 \muldiv.mul8.FA_P14A7B5.genblk1.fa_1  (.A(\muldiv.mul8.FA_P14A7B4.SUM ),
    .B(\muldiv.mul8.FA_P13A7B5.B ),
    .CIN(\muldiv.mul8.FA_P13A7B5.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.mul8.FA_P14A7B5.COUT ),
    .SUM(\muldiv.mul8.FA_P14A7B5.SUM ));
 sky130_fd_sc_hd__fa_1 \muldiv.mul8.FA_P14A7B6.genblk1.fa_1  (.A(\muldiv.mul8.FA_P14A7B5.SUM ),
    .B(\muldiv.mul8.FA_P14A7B6.B ),
    .CIN(\muldiv.mul8.FA_P13A7B6.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.mul8.FA_P14A7B6.COUT ),
    .SUM(\muldiv.mul8.FA_P14A7B6.SUM ));
 sky130_fd_sc_hd__fa_1 \muldiv.mul8.FA_P14A7B7.genblk1.fa_1  (.A(\muldiv.mul8.FA_P14A7B6.SUM ),
    .B(\muldiv.mul8.FA_P14A7B7.B ),
    .CIN(\muldiv.mul8.FA_P13A6B7.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.mul8.FA_P14A7B7.COUT ),
    .SUM(\muldiv.mul8.FA_P14A7B7.SUM ));
 sky130_fd_sc_hd__fa_1 \muldiv.mul8.FA_P15A7B1.genblk1.fa_1  (.A(\muldiv.mul8.FA_P10A7B1.A ),
    .B(\muldiv.mul8.FA_P10A7B1.B ),
    .CIN(\muldiv.mul8.FA_P14A7B1.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.mul8.FA_P15A7B1.COUT ),
    .SUM(\muldiv.mul8.FA_P15A7B1.SUM ));
 sky130_fd_sc_hd__fa_1 \muldiv.mul8.FA_P15A7B2.genblk1.fa_1  (.A(\muldiv.mul8.FA_P15A7B1.SUM ),
    .B(\muldiv.mul8.FA_P10A7B2.B ),
    .CIN(\muldiv.mul8.FA_P14A7B2.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.mul8.FA_P15A7B2.COUT ),
    .SUM(\muldiv.mul8.FA_P15A7B2.SUM ));
 sky130_fd_sc_hd__fa_1 \muldiv.mul8.FA_P15A7B3.genblk1.fa_1  (.A(\muldiv.mul8.FA_P15A7B2.SUM ),
    .B(\muldiv.mul8.FA_P11A7B3.B ),
    .CIN(\muldiv.mul8.FA_P14A7B3.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.mul8.FA_P15A7B3.COUT ),
    .SUM(\muldiv.mul8.FA_P15A7B3.SUM ));
 sky130_fd_sc_hd__fa_1 \muldiv.mul8.FA_P15A7B4.genblk1.fa_1  (.A(\muldiv.mul8.FA_P15A7B3.SUM ),
    .B(\muldiv.mul8.FA_P12A7B4.B ),
    .CIN(\muldiv.mul8.FA_P14A7B4.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.mul8.FA_P15A7B4.COUT ),
    .SUM(\muldiv.mul8.FA_P15A7B4.SUM ));
 sky130_fd_sc_hd__fa_1 \muldiv.mul8.FA_P15A7B5.genblk1.fa_1  (.A(\muldiv.mul8.FA_P15A7B4.SUM ),
    .B(\muldiv.mul8.FA_P13A7B5.B ),
    .CIN(\muldiv.mul8.FA_P14A7B5.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.mul8.FA_P15A7B5.COUT ),
    .SUM(\muldiv.mul8.FA_P15A7B5.SUM ));
 sky130_fd_sc_hd__fa_1 \muldiv.mul8.FA_P15A7B6.genblk1.fa_1  (.A(\muldiv.mul8.FA_P15A7B5.SUM ),
    .B(\muldiv.mul8.FA_P14A7B6.B ),
    .CIN(\muldiv.mul8.FA_P14A7B6.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.mul8.FA_P15A7B6.COUT ),
    .SUM(\muldiv.mul8.FA_P15A7B6.SUM ));
 sky130_fd_sc_hd__fa_1 \muldiv.mul8.FA_P15A7B7.genblk1.fa_1  (.A(\muldiv.mul8.FA_P15A7B6.SUM ),
    .B(\muldiv.mul8.FA_P15A7B7.B ),
    .CIN(\muldiv.mul8.FA_P14A7B7.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.mul8.FA_P15A7B7.COUT ),
    .SUM(\muldiv.mul8.FA_P15A7B7.SUM ));
 sky130_fd_sc_hd__fa_1 \muldiv.mul8.FA_P2A1B1.genblk1.fa_1  (.A(\muldiv.mul8.A2xB0_2 ),
    .B(\muldiv.mul8.A1xB1_9 ),
    .CIN(\muldiv.mul8.FA_P2A1B1.CIN ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.mul8.FA_P2A1B1.COUT ),
    .SUM(\muldiv.mul8.FA_P2A1B1.SUM ));
 sky130_fd_sc_hd__fa_1 \muldiv.mul8.FA_P3A1B2.genblk1.fa_1  (.A(\muldiv.mul8.FA_P3A1B2.A ),
    .B(\muldiv.mul8.A1xB2_17 ),
    .CIN(\muldiv.mul8.FA_P3A1B2.CIN ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.mul8.FA_P3A1B2.COUT ),
    .SUM(\muldiv.mul8.FA_P3A1B2.SUM ));
 sky130_fd_sc_hd__fa_1 \muldiv.mul8.FA_P3A2B1.genblk1.fa_1  (.A(\muldiv.mul8.A3xB0_3 ),
    .B(\muldiv.mul8.A2xB1_10 ),
    .CIN(\muldiv.mul8.FA_P2A1B1.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.mul8.FA_P3A2B1.COUT ),
    .SUM(\muldiv.mul8.FA_P3A1B2.A ));
 sky130_fd_sc_hd__fa_2 \muldiv.mul8.FA_P4A1B3.genblk1.fa_1  (.A(\muldiv.mul8.FA_P4A1B3.A ),
    .B(\muldiv.mul8.A1xB3_25 ),
    .CIN(\muldiv.mul8.FA_P4A1B3.CIN ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.mul8.FA_P4A1B3.COUT ),
    .SUM(\muldiv.mul8.FA_P4A1B3.SUM ));
 sky130_fd_sc_hd__fa_2 \muldiv.mul8.FA_P4A2B2.genblk1.fa_1  (.A(\muldiv.mul8.FA_P4A2B2.A ),
    .B(\muldiv.mul8.A2xB2_18 ),
    .CIN(\muldiv.mul8.FA_P3A1B2.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.mul8.FA_P4A2B2.COUT ),
    .SUM(\muldiv.mul8.FA_P4A1B3.A ));
 sky130_fd_sc_hd__fa_2 \muldiv.mul8.FA_P4A3B1.genblk1.fa_1  (.A(\muldiv.mul8.A4xB0_4 ),
    .B(\muldiv.mul8.A3xB1_11 ),
    .CIN(\muldiv.mul8.FA_P3A2B1.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.mul8.FA_P4A3B1.COUT ),
    .SUM(\muldiv.mul8.FA_P4A2B2.A ));
 sky130_fd_sc_hd__fa_1 \muldiv.mul8.FA_P5A1B4.genblk1.fa_1  (.A(\muldiv.mul8.FA_P5A1B4.A ),
    .B(\muldiv.mul8.A1xB4_33 ),
    .CIN(\muldiv.mul8.FA_P5A1B4.CIN ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.mul8.FA_P5A1B4.COUT ),
    .SUM(\muldiv.mul8.FA_P5A1B4.SUM ));
 sky130_fd_sc_hd__fa_1 \muldiv.mul8.FA_P5A2B3.genblk1.fa_1  (.A(\muldiv.mul8.FA_P5A2B3.A ),
    .B(\muldiv.mul8.A2xB3_26 ),
    .CIN(\muldiv.mul8.FA_P4A1B3.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.mul8.FA_P5A2B3.COUT ),
    .SUM(\muldiv.mul8.FA_P5A1B4.A ));
 sky130_fd_sc_hd__fa_1 \muldiv.mul8.FA_P5A3B2.genblk1.fa_1  (.A(\muldiv.mul8.FA_P5A3B2.A ),
    .B(\muldiv.mul8.A3xB2_19 ),
    .CIN(\muldiv.mul8.FA_P4A2B2.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.mul8.FA_P5A3B2.COUT ),
    .SUM(\muldiv.mul8.FA_P5A2B3.A ));
 sky130_fd_sc_hd__fa_1 \muldiv.mul8.FA_P5A4B1.genblk1.fa_1  (.A(\muldiv.mul8.A5xB0_5 ),
    .B(\muldiv.mul8.A4xB1_12 ),
    .CIN(\muldiv.mul8.FA_P4A3B1.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.mul8.FA_P5A4B1.COUT ),
    .SUM(\muldiv.mul8.FA_P5A3B2.A ));
 sky130_fd_sc_hd__fa_1 \muldiv.mul8.FA_P6A1B5.genblk1.fa_1  (.A(\muldiv.mul8.FA_P6A1B5.A ),
    .B(\muldiv.mul8.A1xB5_41 ),
    .CIN(\muldiv.mul8.FA_P6A1B5.CIN ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.mul8.FA_P6A1B5.COUT ),
    .SUM(\muldiv.mul8.FA_P6A1B5.SUM ));
 sky130_fd_sc_hd__fa_1 \muldiv.mul8.FA_P6A2B4.genblk1.fa_1  (.A(\muldiv.mul8.FA_P6A2B4.A ),
    .B(\muldiv.mul8.A2xB4_34 ),
    .CIN(\muldiv.mul8.FA_P5A1B4.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.mul8.FA_P6A2B4.COUT ),
    .SUM(\muldiv.mul8.FA_P6A1B5.A ));
 sky130_fd_sc_hd__fa_1 \muldiv.mul8.FA_P6A3B3.genblk1.fa_1  (.A(\muldiv.mul8.FA_P6A3B3.A ),
    .B(\muldiv.mul8.A3xB3_27 ),
    .CIN(\muldiv.mul8.FA_P5A2B3.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.mul8.FA_P6A3B3.COUT ),
    .SUM(\muldiv.mul8.FA_P6A2B4.A ));
 sky130_fd_sc_hd__fa_1 \muldiv.mul8.FA_P6A4B2.genblk1.fa_1  (.A(\muldiv.mul8.FA_P6A4B2.A ),
    .B(\muldiv.mul8.A4xB2_20 ),
    .CIN(\muldiv.mul8.FA_P5A3B2.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.mul8.FA_P6A4B2.COUT ),
    .SUM(\muldiv.mul8.FA_P6A3B3.A ));
 sky130_fd_sc_hd__fa_1 \muldiv.mul8.FA_P6A5B1.genblk1.fa_1  (.A(\muldiv.mul8.A6xB0_6 ),
    .B(\muldiv.mul8.A5xB1_13 ),
    .CIN(\muldiv.mul8.FA_P5A4B1.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.mul8.FA_P6A5B1.COUT ),
    .SUM(\muldiv.mul8.FA_P6A4B2.A ));
 sky130_fd_sc_hd__fa_1 \muldiv.mul8.FA_P7A0B7.genblk1.fa_1  (.A(\muldiv.mul8.FA_P7A0B7.A ),
    .B(\muldiv.mul8.FA_P7A0B7.B ),
    .CIN(\muldiv.div8.HAD_DVD_TWOS_0.B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.mul8.FA_P7A0B7.COUT ),
    .SUM(\muldiv.mul8.FA_P7A0B7.SUM ));
 sky130_fd_sc_hd__fa_1 \muldiv.mul8.FA_P7A1B6.genblk1.fa_1  (.A(\muldiv.mul8.FA_P7A1B6.A ),
    .B(\muldiv.mul8.A1xB6_49 ),
    .CIN(\muldiv.mul8.FA_P7A1B6.CIN ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.mul8.FA_P7A1B6.COUT ),
    .SUM(\muldiv.mul8.FA_P7A0B7.A ));
 sky130_fd_sc_hd__fa_1 \muldiv.mul8.FA_P7A2B5.genblk1.fa_1  (.A(\muldiv.mul8.FA_P7A2B5.A ),
    .B(\muldiv.mul8.A2xB5_42 ),
    .CIN(\muldiv.mul8.FA_P6A1B5.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.mul8.FA_P7A2B5.COUT ),
    .SUM(\muldiv.mul8.FA_P7A1B6.A ));
 sky130_fd_sc_hd__fa_1 \muldiv.mul8.FA_P7A3B4.genblk1.fa_1  (.A(\muldiv.mul8.FA_P7A3B4.A ),
    .B(\muldiv.mul8.A3xB4_35 ),
    .CIN(\muldiv.mul8.FA_P6A2B4.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.mul8.FA_P7A3B4.COUT ),
    .SUM(\muldiv.mul8.FA_P7A2B5.A ));
 sky130_fd_sc_hd__fa_1 \muldiv.mul8.FA_P7A4B3.genblk1.fa_1  (.A(\muldiv.mul8.FA_P7A4B3.A ),
    .B(\muldiv.mul8.A4xB3_28 ),
    .CIN(\muldiv.mul8.FA_P6A3B3.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.mul8.FA_P7A4B3.COUT ),
    .SUM(\muldiv.mul8.FA_P7A3B4.A ));
 sky130_fd_sc_hd__fa_1 \muldiv.mul8.FA_P7A5B2.genblk1.fa_1  (.A(\muldiv.mul8.FA_P7A5B2.A ),
    .B(\muldiv.mul8.A5xB2_21 ),
    .CIN(\muldiv.mul8.FA_P6A4B2.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.mul8.FA_P7A5B2.COUT ),
    .SUM(\muldiv.mul8.FA_P7A4B3.A ));
 sky130_fd_sc_hd__fa_1 \muldiv.mul8.FA_P7A6B1.genblk1.fa_1  (.A(\muldiv.mul8.A7xB0_7 ),
    .B(\muldiv.mul8.A6xB1_14 ),
    .CIN(\muldiv.mul8.FA_P6A5B1.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.mul8.FA_P7A6B1.COUT ),
    .SUM(\muldiv.mul8.FA_P7A5B2.A ));
 sky130_fd_sc_hd__fa_1 \muldiv.mul8.FA_P8A1B7.genblk1.fa_1  (.A(\muldiv.mul8.FA_P8A1B7.A ),
    .B(\muldiv.mul8.FA_P8A1B7.B ),
    .CIN(\muldiv.mul8.FA_P7A0B7.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.mul8.FA_P8A1B7.COUT ),
    .SUM(\muldiv.mul8.FA_P8A1B7.SUM ));
 sky130_fd_sc_hd__fa_1 \muldiv.mul8.FA_P8A2B6.genblk1.fa_1  (.A(\muldiv.mul8.FA_P8A2B6.A ),
    .B(\muldiv.mul8.A2xB6_50 ),
    .CIN(\muldiv.mul8.FA_P7A1B6.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.mul8.FA_P8A2B6.COUT ),
    .SUM(\muldiv.mul8.FA_P8A1B7.A ));
 sky130_fd_sc_hd__fa_1 \muldiv.mul8.FA_P8A3B5.genblk1.fa_1  (.A(\muldiv.mul8.FA_P8A3B5.A ),
    .B(\muldiv.mul8.A3xB5_43 ),
    .CIN(\muldiv.mul8.FA_P7A2B5.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.mul8.FA_P8A3B5.COUT ),
    .SUM(\muldiv.mul8.FA_P8A2B6.A ));
 sky130_fd_sc_hd__fa_1 \muldiv.mul8.FA_P8A4B4.genblk1.fa_1  (.A(\muldiv.mul8.FA_P8A4B4.A ),
    .B(\muldiv.mul8.A4xB4_36 ),
    .CIN(\muldiv.mul8.FA_P7A3B4.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.mul8.FA_P8A4B4.COUT ),
    .SUM(\muldiv.mul8.FA_P8A3B5.A ));
 sky130_fd_sc_hd__fa_1 \muldiv.mul8.FA_P8A5B3.genblk1.fa_1  (.A(\muldiv.mul8.FA_P8A5B3.A ),
    .B(\muldiv.mul8.A5xB3_29 ),
    .CIN(\muldiv.mul8.FA_P7A4B3.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.mul8.FA_P8A5B3.COUT ),
    .SUM(\muldiv.mul8.FA_P8A4B4.A ));
 sky130_fd_sc_hd__fa_1 \muldiv.mul8.FA_P8A6B2.genblk1.fa_1  (.A(\muldiv.mul8.FA_P8A6B2.A ),
    .B(\muldiv.mul8.A6xB2_22 ),
    .CIN(\muldiv.mul8.FA_P7A5B2.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.mul8.FA_P8A6B2.COUT ),
    .SUM(\muldiv.mul8.FA_P8A5B3.A ));
 sky130_fd_sc_hd__fa_1 \muldiv.mul8.FA_P8A7B1.genblk1.fa_1  (.A(\muldiv.mul8.FA_P10A7B1.A ),
    .B(\muldiv.mul8.A7xB1_15 ),
    .CIN(\muldiv.mul8.FA_P7A6B1.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.mul8.FA_P8A7B1.COUT ),
    .SUM(\muldiv.mul8.FA_P8A6B2.A ));
 sky130_fd_sc_hd__fa_1 \muldiv.mul8.FA_P9A2B7.genblk1.fa_1  (.A(\muldiv.mul8.FA_P9A2B7.A ),
    .B(\muldiv.mul8.FA_P9A2B7.B ),
    .CIN(\muldiv.mul8.FA_P8A1B7.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.mul8.FA_P10A3B7.CIN ),
    .SUM(\muldiv.mul8.FA_P9A2B7.SUM ));
 sky130_fd_sc_hd__fa_1 \muldiv.mul8.FA_P9A3B6.genblk1.fa_1  (.A(\muldiv.mul8.FA_P9A3B6.A ),
    .B(\muldiv.mul8.A3xB6_51 ),
    .CIN(\muldiv.mul8.FA_P8A2B6.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.mul8.FA_P10A4B6.CIN ),
    .SUM(\muldiv.mul8.FA_P9A2B7.A ));
 sky130_fd_sc_hd__fa_1 \muldiv.mul8.FA_P9A4B5.genblk1.fa_1  (.A(\muldiv.mul8.FA_P9A4B5.A ),
    .B(\muldiv.mul8.A4xB5_44 ),
    .CIN(\muldiv.mul8.FA_P8A3B5.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.mul8.FA_P10A5B5.CIN ),
    .SUM(\muldiv.mul8.FA_P9A3B6.A ));
 sky130_fd_sc_hd__fa_1 \muldiv.mul8.FA_P9A5B4.genblk1.fa_1  (.A(\muldiv.mul8.FA_P9A5B4.A ),
    .B(\muldiv.mul8.A5xB4_37 ),
    .CIN(\muldiv.mul8.FA_P8A4B4.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.mul8.FA_P10A6B4.CIN ),
    .SUM(\muldiv.mul8.FA_P9A4B5.A ));
 sky130_fd_sc_hd__fa_1 \muldiv.mul8.FA_P9A6B3.genblk1.fa_1  (.A(\muldiv.mul8.FA_P9A6B3.A ),
    .B(\muldiv.mul8.A6xB3_30 ),
    .CIN(\muldiv.mul8.FA_P8A5B3.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.mul8.FA_P10A7B3.CIN ),
    .SUM(\muldiv.mul8.FA_P9A5B4.A ));
 sky130_fd_sc_hd__fa_1 \muldiv.mul8.FA_P9A7B1.genblk1.fa_1  (.A(\muldiv.mul8.FA_P10A7B1.A ),
    .B(\muldiv.mul8.FA_P10A7B1.B ),
    .CIN(\muldiv.mul8.FA_P8A7B1.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.mul8.FA_P10A7B1.CIN ),
    .SUM(\muldiv.mul8.FA_P9A7B1.SUM ));
 sky130_fd_sc_hd__fa_1 \muldiv.mul8.FA_P9A7B2.genblk1.fa_1  (.A(\muldiv.mul8.FA_P9A7B1.SUM ),
    .B(\muldiv.mul8.A7xB2_23 ),
    .CIN(\muldiv.mul8.FA_P8A6B2.COUT ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.mul8.FA_P10A7B2.CIN ),
    .SUM(\muldiv.mul8.FA_P9A6B3.A ));
 sky130_fd_sc_hd__ha_1 \muldiv.mul8.HA_P1A0B1.genblk1.ha_1  (.A(\muldiv.mul8.A1xB0_1 ),
    .B(\muldiv.mul8.A0xB1_8 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.mul8.FA_P2A1B1.CIN ),
    .SUM(\muldiv.mul8.HA_P1A0B1.SUM ));
 sky130_fd_sc_hd__ha_1 \muldiv.mul8.HA_P2A0B2.genblk1.ha_1  (.A(\muldiv.mul8.FA_P2A1B1.SUM ),
    .B(\muldiv.mul8.A0xB2_16 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.mul8.FA_P3A1B2.CIN ),
    .SUM(\muldiv.mul8.HA_P2A0B2.SUM ));
 sky130_fd_sc_hd__ha_1 \muldiv.mul8.HA_P3A0B3.genblk1.ha_1  (.A(\muldiv.mul8.FA_P3A1B2.SUM ),
    .B(\muldiv.mul8.A0xB3_24 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.mul8.FA_P4A1B3.CIN ),
    .SUM(\muldiv.mul8.HA_P3A0B3.SUM ));
 sky130_fd_sc_hd__ha_1 \muldiv.mul8.HA_P4A0B4.genblk1.ha_1  (.A(\muldiv.mul8.FA_P4A1B3.SUM ),
    .B(\muldiv.mul8.A0xB4_32 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.mul8.FA_P5A1B4.CIN ),
    .SUM(\muldiv.mul8.HA_P4A0B4.SUM ));
 sky130_fd_sc_hd__ha_1 \muldiv.mul8.HA_P5A0B5.genblk1.ha_1  (.A(\muldiv.mul8.FA_P5A1B4.SUM ),
    .B(\muldiv.mul8.A0xB5_40 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.mul8.FA_P6A1B5.CIN ),
    .SUM(\muldiv.mul8.HA_P5A0B5.SUM ));
 sky130_fd_sc_hd__ha_1 \muldiv.mul8.HA_P6A0B6.genblk1.ha_1  (.A(\muldiv.mul8.FA_P6A1B5.SUM ),
    .B(\muldiv.mul8.A0xB6_48 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .COUT(\muldiv.mul8.FA_P7A1B6.CIN ),
    .SUM(\muldiv.mul8.HA_P6A0B6.SUM ));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer1 (.A(\muldiv.div8.DU_Q6D6d0.io_sel ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net96));
 sky130_fd_sc_hd__buf_1 rebuffer12 (.A(\muldiv.div8.DU_Q7D7d0.io_sel ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net78));
 sky130_fd_sc_hd__clkbuf_1 rebuffer13 (.A(net78),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net79));
 sky130_fd_sc_hd__clkbuf_1 rebuffer2 (.A(net70),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net68));
 sky130_fd_sc_hd__clkbuf_1 rebuffer3 (.A(net70),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net69));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer4 (.A(\muldiv.div8.DU_Q6D6d0.io_sel ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net97));
 sky130_fd_sc_hd__buf_1 rebuffer6 (.A(net78),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net72));
 sky130_fd_sc_hd__clkbuf_1 rebuffer7 (.A(net97),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net73));
 sky130_fd_sc_hd__clkbuf_1 rebuffer8 (.A(\muldiv.div8.DU_Q6D6d0.io_sel ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net74));
 sky130_fd_sc_hd__clkbuf_2 split1 (.A(\muldiv.div8.DU_Q0D0d0.io_sel ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net67));
 sky130_fd_sc_hd__dlymetal6s2s_1 split4 (.A(\muldiv.div8.DU_Q5D5d0.io_sel ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net70));
 sky130_fd_sc_hd__conb_1 tt_um_dlmiles_muldiv8_sky130faha_32 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net32));
 sky130_fd_sc_hd__conb_1 tt_um_dlmiles_muldiv8_sky130faha_33 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net33));
 sky130_fd_sc_hd__conb_1 tt_um_dlmiles_muldiv8_sky130faha_34 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net34));
 sky130_fd_sc_hd__conb_1 tt_um_dlmiles_muldiv8_sky130faha_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net35));
 sky130_fd_sc_hd__conb_1 tt_um_dlmiles_muldiv8_sky130faha_36 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net36));
 sky130_fd_sc_hd__conb_1 tt_um_dlmiles_muldiv8_sky130faha_37 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net37));
 sky130_fd_sc_hd__conb_1 tt_um_dlmiles_muldiv8_sky130faha_38 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net38));
 sky130_fd_sc_hd__conb_1 tt_um_dlmiles_muldiv8_sky130faha_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net39));
 sky130_fd_sc_hd__conb_1 tt_um_dlmiles_muldiv8_sky130faha_40 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net40));
 sky130_fd_sc_hd__conb_1 tt_um_dlmiles_muldiv8_sky130faha_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net41));
 sky130_fd_sc_hd__conb_1 tt_um_dlmiles_muldiv8_sky130faha_42 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net42));
 sky130_fd_sc_hd__conb_1 tt_um_dlmiles_muldiv8_sky130faha_43 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net43));
 sky130_fd_sc_hd__conb_1 tt_um_dlmiles_muldiv8_sky130faha_64 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(net64));
 sky130_fd_sc_hd__conb_1 tt_um_dlmiles_muldiv8_sky130faha_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(net65));
 assign uio_oe[0] = net32;
 assign uio_oe[1] = net33;
 assign uio_oe[2] = net34;
 assign uio_oe[3] = net35;
 assign uio_oe[4] = net64;
 assign uio_oe[5] = net65;
 assign uio_oe[6] = net36;
 assign uio_oe[7] = net37;
 assign uio_out[0] = net38;
 assign uio_out[1] = net39;
 assign uio_out[2] = net40;
 assign uio_out[3] = net41;
 assign uio_out[6] = net42;
 assign uio_out[7] = net43;
endmodule
