VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_algofoogle_tt06_grab_bag
  CLASS BLOCK ;
  FOREIGN tt_um_algofoogle_tt06_grab_bag ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 154.870 224.760 155.170 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 158.550 224.760 158.850 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 151.190 224.760 151.490 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.480000 ;
    PORT
      LAYER met4 ;
        RECT 156.560 0.000 157.160 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 134.480 0.000 135.080 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 112.400 0.000 113.000 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 90.320 0.000 90.920 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 68.240 0.000 68.840 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 46.160 0.000 46.760 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 24.080 0.000 24.680 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 2.000 0.000 2.600 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.800000 ;
    PORT
      LAYER met4 ;
        RECT 147.510 224.760 147.810 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 140.150 224.760 140.450 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 136.470 224.760 136.770 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 129.110 224.760 129.410 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 125.430 224.760 125.730 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.070 224.760 118.370 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 114.390 224.760 114.690 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.030 224.760 107.330 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 103.350 224.760 103.650 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 95.990 224.760 96.290 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 92.310 224.760 92.610 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.591000 ;
    PORT
      LAYER met4 ;
        RECT 29.750 224.760 30.050 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.591000 ;
    PORT
      LAYER met4 ;
        RECT 26.070 224.760 26.370 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.591000 ;
    PORT
      LAYER met4 ;
        RECT 22.390 224.760 22.690 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.591000 ;
    PORT
      LAYER met4 ;
        RECT 18.710 224.760 19.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.591000 ;
    PORT
      LAYER met4 ;
        RECT 15.030 224.760 15.330 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.591000 ;
    PORT
      LAYER met4 ;
        RECT 11.350 224.760 11.650 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.591000 ;
    PORT
      LAYER met4 ;
        RECT 7.670 224.760 7.970 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.591000 ;
    PORT
      LAYER met4 ;
        RECT 3.990 224.760 4.290 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.591000 ;
    PORT
      LAYER met4 ;
        RECT 59.190 224.760 59.490 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.591000 ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.591000 ;
    PORT
      LAYER met4 ;
        RECT 51.830 224.760 52.130 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.591000 ;
    PORT
      LAYER met4 ;
        RECT 48.150 224.760 48.450 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.591000 ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.591000 ;
    PORT
      LAYER met4 ;
        RECT 40.790 224.760 41.090 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.591000 ;
    PORT
      LAYER met4 ;
        RECT 37.110 224.760 37.410 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.591000 ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.480000 ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.591000 ;
    PORT
      LAYER met4 ;
        RECT 84.950 224.760 85.250 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.591000 ;
    PORT
      LAYER met4 ;
        RECT 81.270 224.760 81.570 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.591000 ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.591000 ;
    PORT
      LAYER met4 ;
        RECT 73.910 224.760 74.210 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.591000 ;
    PORT
      LAYER met4 ;
        RECT 70.230 224.760 70.530 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.591000 ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.591000 ;
    PORT
      LAYER met4 ;
        RECT 62.870 224.760 63.170 225.760 ;
    END
  END uo_out[7]
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 2.500 220.760 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 49.000 5.000 50.500 220.760 ;
    END
  END VGND
  OBS
      LAYER nwell ;
        RECT 144.215 24.870 146.325 35.060 ;
      LAYER pwell ;
        RECT 147.030 26.935 149.140 33.035 ;
      LAYER li1 ;
        RECT 144.395 34.710 146.145 34.880 ;
        RECT 144.395 30.535 144.565 34.710 ;
        RECT 145.105 34.200 145.435 34.370 ;
        RECT 144.330 29.835 144.630 30.535 ;
        RECT 144.395 25.220 144.565 29.835 ;
        RECT 144.965 25.945 145.135 33.985 ;
        RECT 145.405 25.945 145.575 33.985 ;
        RECT 145.105 25.560 145.435 25.730 ;
        RECT 145.975 25.220 146.145 34.710 ;
        RECT 147.210 32.685 148.960 32.855 ;
        RECT 147.210 27.285 147.380 32.685 ;
        RECT 147.920 32.175 148.250 32.345 ;
        RECT 147.780 27.965 147.950 32.005 ;
        RECT 148.220 27.965 148.390 32.005 ;
        RECT 148.790 31.735 148.960 32.685 ;
        RECT 148.730 30.935 149.030 31.735 ;
        RECT 147.920 27.625 148.250 27.795 ;
        RECT 148.790 27.285 148.960 30.935 ;
        RECT 147.210 27.115 148.960 27.285 ;
        RECT 144.395 25.050 146.145 25.220 ;
      LAYER mcon ;
        RECT 145.185 34.200 145.355 34.370 ;
        RECT 144.330 29.835 144.630 30.535 ;
        RECT 144.965 26.025 145.135 33.905 ;
        RECT 145.405 26.025 145.575 33.905 ;
        RECT 145.185 25.560 145.355 25.730 ;
        RECT 148.000 32.175 148.170 32.345 ;
        RECT 147.780 28.045 147.950 31.925 ;
        RECT 148.220 28.045 148.390 31.925 ;
        RECT 148.730 30.935 149.030 31.735 ;
        RECT 148.000 27.625 148.170 27.795 ;
      LAYER met1 ;
        RECT 88.300 208.050 89.300 216.330 ;
        RECT 88.300 207.050 99.550 208.050 ;
        RECT 98.550 40.950 99.550 207.050 ;
        RECT 98.520 39.950 99.580 40.950 ;
        RECT 147.160 38.430 148.160 222.100 ;
        RECT 147.160 37.430 152.050 38.430 ;
        RECT 147.160 37.400 148.160 37.430 ;
        RECT 57.990 35.185 150.580 36.185 ;
        RECT 145.130 34.400 148.230 34.435 ;
        RECT 145.125 34.170 148.230 34.400 ;
        RECT 145.130 34.135 148.230 34.170 ;
        RECT 144.935 30.685 145.165 33.965 ;
        RECT 145.375 30.935 145.605 33.965 ;
        RECT 147.930 32.435 148.230 34.135 ;
        RECT 149.130 32.435 149.430 32.465 ;
        RECT 147.830 32.135 149.430 32.435 ;
        RECT 149.130 32.105 149.430 32.135 ;
        RECT 147.750 30.935 147.980 31.985 ;
        RECT 148.190 31.835 148.420 31.985 ;
        RECT 149.580 31.835 150.580 35.185 ;
        RECT 10.510 29.685 145.180 30.685 ;
        RECT 145.375 29.685 147.980 30.935 ;
        RECT 148.180 30.835 150.580 31.835 ;
        RECT 144.935 25.965 145.165 29.685 ;
        RECT 145.375 25.965 145.605 29.685 ;
        RECT 146.580 26.435 146.880 29.685 ;
        RECT 147.750 27.985 147.980 29.685 ;
        RECT 148.190 27.985 148.420 30.835 ;
        RECT 151.020 30.450 152.020 37.430 ;
        RECT 149.600 30.435 152.020 30.450 ;
        RECT 149.130 30.085 149.430 30.115 ;
        RECT 149.580 30.085 152.020 30.435 ;
        RECT 149.130 29.785 152.020 30.085 ;
        RECT 149.130 29.755 149.430 29.785 ;
        RECT 149.580 29.460 152.020 29.785 ;
        RECT 149.580 29.435 150.580 29.460 ;
        RECT 149.130 27.835 149.430 27.865 ;
        RECT 147.830 27.535 149.430 27.835 ;
        RECT 147.430 26.435 147.730 26.465 ;
        RECT 146.580 26.135 147.730 26.435 ;
        RECT 147.430 26.105 147.730 26.135 ;
        RECT 147.930 25.785 148.230 27.535 ;
        RECT 149.130 27.505 149.430 27.535 ;
        RECT 149.580 26.435 150.580 26.785 ;
        RECT 148.450 26.135 150.580 26.435 ;
        RECT 145.080 25.485 148.230 25.785 ;
        RECT 98.550 23.850 99.550 23.880 ;
        RECT 149.580 23.850 150.580 26.135 ;
        RECT 98.550 22.850 150.580 23.850 ;
        RECT 98.550 22.820 99.550 22.850 ;
        RECT 149.580 10.350 150.580 22.850 ;
        RECT 156.350 10.350 157.350 10.380 ;
        RECT 149.580 9.350 157.350 10.350 ;
        RECT 156.350 9.320 157.350 9.350 ;
      LAYER via ;
        RECT 147.510 221.750 147.810 222.050 ;
        RECT 88.300 215.300 89.300 216.300 ;
        RECT 98.550 39.950 99.550 40.950 ;
        RECT 58.020 35.185 59.020 36.185 ;
        RECT 149.130 32.135 149.430 32.435 ;
        RECT 10.540 29.685 11.540 30.685 ;
        RECT 149.130 27.535 149.430 27.835 ;
        RECT 147.430 26.135 147.730 26.435 ;
        RECT 148.480 26.135 148.780 26.435 ;
        RECT 156.350 9.350 157.350 10.350 ;
      LAYER met2 ;
        RECT 147.510 222.950 147.810 222.960 ;
        RECT 147.475 222.670 147.845 222.950 ;
        RECT 147.510 221.720 147.810 222.670 ;
        RECT 88.300 216.300 89.300 218.545 ;
        RECT 88.270 215.300 89.330 216.300 ;
        RECT 58.020 36.185 59.020 36.215 ;
        RECT 55.735 35.185 59.020 36.185 ;
        RECT 58.020 35.155 59.020 35.185 ;
        RECT 10.540 30.685 11.540 30.715 ;
        RECT 8.055 29.685 11.540 30.685 ;
        RECT 10.540 29.655 11.540 29.685 ;
        RECT 98.550 23.850 99.550 40.980 ;
        RECT 149.100 32.135 149.460 32.435 ;
        RECT 149.130 30.085 149.430 32.135 ;
        RECT 149.100 29.785 149.460 30.085 ;
        RECT 149.130 27.835 149.430 29.785 ;
        RECT 149.100 27.535 149.460 27.835 ;
        RECT 148.480 26.435 148.780 26.465 ;
        RECT 147.400 26.135 148.780 26.435 ;
        RECT 148.480 26.105 148.780 26.135 ;
        RECT 98.520 22.850 99.580 23.850 ;
        RECT 156.320 9.350 157.380 10.350 ;
        RECT 156.350 7.255 157.350 9.350 ;
      LAYER via2 ;
        RECT 147.520 222.670 147.800 222.950 ;
        RECT 88.300 217.500 89.300 218.500 ;
        RECT 55.780 35.185 56.780 36.185 ;
        RECT 8.100 29.685 9.100 30.685 ;
        RECT 156.350 7.300 157.350 8.300 ;
      LAYER met3 ;
        RECT 147.470 223.760 147.850 224.080 ;
        RECT 147.510 222.975 147.810 223.760 ;
        RECT 147.495 222.645 147.825 222.975 ;
        RECT 88.300 218.525 89.300 220.480 ;
        RECT 88.275 217.475 89.325 218.525 ;
        RECT 55.755 36.185 56.805 36.210 ;
        RECT 53.320 35.185 56.805 36.185 ;
        RECT 55.755 35.160 56.805 35.185 ;
        RECT 8.075 30.685 9.125 30.710 ;
        RECT 5.390 29.685 9.125 30.685 ;
        RECT 8.075 29.660 9.125 29.685 ;
        RECT 156.325 7.275 157.375 8.325 ;
        RECT 156.350 5.170 157.350 7.275 ;
      LAYER via3 ;
        RECT 147.500 223.760 147.820 224.080 ;
        RECT 88.300 219.450 89.300 220.450 ;
        RECT 53.350 35.185 54.350 36.185 ;
        RECT 5.420 29.685 6.420 30.685 ;
        RECT 156.350 5.200 157.350 6.200 ;
      LAYER met4 ;
        RECT 3.990 222.190 4.290 224.760 ;
        RECT 7.670 222.190 7.970 224.760 ;
        RECT 11.350 222.190 11.650 224.760 ;
        RECT 15.030 222.190 15.330 224.760 ;
        RECT 18.710 222.190 19.010 224.760 ;
        RECT 22.390 222.190 22.690 224.760 ;
        RECT 26.070 222.190 26.370 224.760 ;
        RECT 29.750 222.190 30.050 224.760 ;
        RECT 33.430 222.190 33.730 224.760 ;
        RECT 37.110 222.190 37.410 224.760 ;
        RECT 40.790 222.190 41.090 224.760 ;
        RECT 44.470 222.190 44.770 224.760 ;
        RECT 48.150 222.190 48.450 224.760 ;
        RECT 51.830 222.190 52.130 224.760 ;
        RECT 55.510 222.190 55.810 224.760 ;
        RECT 59.190 222.190 59.490 224.760 ;
        RECT 62.870 222.190 63.170 224.760 ;
        RECT 66.550 222.190 66.850 224.760 ;
        RECT 70.230 222.190 70.530 224.760 ;
        RECT 73.910 222.190 74.210 224.760 ;
        RECT 77.590 222.190 77.890 224.760 ;
        RECT 81.270 222.190 81.570 224.760 ;
        RECT 84.950 222.190 85.250 224.760 ;
        RECT 88.630 223.100 88.930 224.760 ;
        RECT 147.510 224.085 147.810 224.760 ;
        RECT 147.495 223.755 147.825 224.085 ;
        RECT 3.740 220.760 85.840 222.190 ;
        RECT 3.740 219.630 49.000 220.760 ;
        RECT 50.500 219.630 85.840 220.760 ;
        RECT 88.300 220.455 89.300 223.100 ;
        RECT 88.295 219.445 89.305 220.455 ;
        RECT 53.345 36.185 54.355 36.190 ;
        RECT 50.500 35.185 54.355 36.185 ;
        RECT 53.345 35.180 54.355 35.185 ;
        RECT 5.415 30.685 6.425 30.690 ;
        RECT 2.500 29.685 6.425 30.685 ;
        RECT 5.415 29.680 6.425 29.685 ;
        RECT 156.345 5.195 157.355 6.205 ;
        RECT 156.530 1.000 157.175 5.195 ;
        RECT 156.530 0.230 156.560 1.000 ;
        RECT 157.160 0.230 157.175 1.000 ;
  END
END tt_um_algofoogle_tt06_grab_bag
END LIBRARY

